VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO multi_project_harness
  CLASS BLOCK ;
  FOREIGN multi_project_harness ;
  ORIGIN 0.000 0.000 ;
  SIZE 1500.000 BY 400.000 ;
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 4.800 1500.000 5.400 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 109.520 1500.000 110.120 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 120.400 1500.000 121.000 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 130.600 1500.000 131.200 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 141.480 1500.000 142.080 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 151.680 1500.000 152.280 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 162.560 1500.000 163.160 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 172.760 1500.000 173.360 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 183.640 1500.000 184.240 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 193.840 1500.000 194.440 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 204.720 1500.000 205.320 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 15.000 1500.000 15.600 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 214.920 1500.000 215.520 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 225.120 1500.000 225.720 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 236.000 1500.000 236.600 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 246.200 1500.000 246.800 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 257.080 1500.000 257.680 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 267.280 1500.000 267.880 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 278.160 1500.000 278.760 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 288.360 1500.000 288.960 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 299.240 1500.000 299.840 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 309.440 1500.000 310.040 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 25.200 1500.000 25.800 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 320.320 1500.000 320.920 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 330.520 1500.000 331.120 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 341.400 1500.000 342.000 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 351.600 1500.000 352.200 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 362.480 1500.000 363.080 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 372.680 1500.000 373.280 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 383.560 1500.000 384.160 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 393.760 1500.000 394.360 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 36.080 1500.000 36.680 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 46.280 1500.000 46.880 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 57.160 1500.000 57.760 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 67.360 1500.000 67.960 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 78.240 1500.000 78.840 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 88.440 1500.000 89.040 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 1496.000 99.320 1500.000 99.920 ;
    END
  END io_in[9]
  PIN io_oeb[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 202.000 4.000 202.600 ;
    END
  END io_oeb[0]
  PIN io_oeb[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END io_oeb[10]
  PIN io_oeb[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 259.800 4.000 260.400 ;
    END
  END io_oeb[11]
  PIN io_oeb[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 264.560 4.000 265.160 ;
    END
  END io_oeb[12]
  PIN io_oeb[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.000 4.000 270.600 ;
    END
  END io_oeb[13]
  PIN io_oeb[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 275.440 4.000 276.040 ;
    END
  END io_oeb[14]
  PIN io_oeb[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 280.880 4.000 281.480 ;
    END
  END io_oeb[15]
  PIN io_oeb[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END io_oeb[16]
  PIN io_oeb[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 291.080 4.000 291.680 ;
    END
  END io_oeb[17]
  PIN io_oeb[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 296.520 4.000 297.120 ;
    END
  END io_oeb[18]
  PIN io_oeb[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END io_oeb[19]
  PIN io_oeb[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 206.760 4.000 207.360 ;
    END
  END io_oeb[1]
  PIN io_oeb[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 306.720 4.000 307.320 ;
    END
  END io_oeb[20]
  PIN io_oeb[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 312.160 4.000 312.760 ;
    END
  END io_oeb[21]
  PIN io_oeb[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 317.600 4.000 318.200 ;
    END
  END io_oeb[22]
  PIN io_oeb[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 322.360 4.000 322.960 ;
    END
  END io_oeb[23]
  PIN io_oeb[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 327.800 4.000 328.400 ;
    END
  END io_oeb[24]
  PIN io_oeb[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END io_oeb[25]
  PIN io_oeb[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 338.680 4.000 339.280 ;
    END
  END io_oeb[26]
  PIN io_oeb[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END io_oeb[27]
  PIN io_oeb[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 348.880 4.000 349.480 ;
    END
  END io_oeb[28]
  PIN io_oeb[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 354.320 4.000 354.920 ;
    END
  END io_oeb[29]
  PIN io_oeb[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 212.200 4.000 212.800 ;
    END
  END io_oeb[2]
  PIN io_oeb[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 359.760 4.000 360.360 ;
    END
  END io_oeb[30]
  PIN io_oeb[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END io_oeb[31]
  PIN io_oeb[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 369.960 4.000 370.560 ;
    END
  END io_oeb[32]
  PIN io_oeb[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 375.400 4.000 376.000 ;
    END
  END io_oeb[33]
  PIN io_oeb[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END io_oeb[34]
  PIN io_oeb[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 385.600 4.000 386.200 ;
    END
  END io_oeb[35]
  PIN io_oeb[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END io_oeb[36]
  PIN io_oeb[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 396.480 4.000 397.080 ;
    END
  END io_oeb[37]
  PIN io_oeb[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END io_oeb[3]
  PIN io_oeb[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 222.400 4.000 223.000 ;
    END
  END io_oeb[4]
  PIN io_oeb[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 227.840 4.000 228.440 ;
    END
  END io_oeb[5]
  PIN io_oeb[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 233.280 4.000 233.880 ;
    END
  END io_oeb[6]
  PIN io_oeb[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.720 4.000 239.320 ;
    END
  END io_oeb[7]
  PIN io_oeb[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 243.480 4.000 244.080 ;
    END
  END io_oeb[8]
  PIN io_oeb[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.920 4.000 249.520 ;
    END
  END io_oeb[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 2.080 4.000 2.680 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 54.440 4.000 55.040 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 59.880 4.000 60.480 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 70.080 4.000 70.680 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 75.520 4.000 76.120 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 80.960 4.000 81.560 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 85.720 4.000 86.320 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 91.160 4.000 91.760 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 96.600 4.000 97.200 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 102.040 4.000 102.640 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 6.840 4.000 7.440 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 106.800 4.000 107.400 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 117.680 4.000 118.280 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 127.880 4.000 128.480 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 133.320 4.000 133.920 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 138.760 4.000 139.360 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 143.520 4.000 144.120 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 148.960 4.000 149.560 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 154.400 4.000 155.000 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 12.280 4.000 12.880 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 164.600 4.000 165.200 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 175.480 4.000 176.080 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 180.920 4.000 181.520 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 185.680 4.000 186.280 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.120 4.000 191.720 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 196.560 4.000 197.160 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.720 4.000 18.320 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 22.480 4.000 23.080 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.920 4.000 28.520 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 33.360 4.000 33.960 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 38.800 4.000 39.400 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 43.560 4.000 44.160 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 49.000 4.000 49.600 ;
    END
  END io_out[9]
  PIN la_data_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 325.770 0.000 326.050 4.000 ;
    END
  END la_data_in[0]
  PIN la_data_in[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1243.930 0.000 1244.210 4.000 ;
    END
  END la_data_in[100]
  PIN la_data_in[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1253.130 0.000 1253.410 4.000 ;
    END
  END la_data_in[101]
  PIN la_data_in[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1262.330 0.000 1262.610 4.000 ;
    END
  END la_data_in[102]
  PIN la_data_in[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1271.530 0.000 1271.810 4.000 ;
    END
  END la_data_in[103]
  PIN la_data_in[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1280.730 0.000 1281.010 4.000 ;
    END
  END la_data_in[104]
  PIN la_data_in[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1289.930 0.000 1290.210 4.000 ;
    END
  END la_data_in[105]
  PIN la_data_in[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1299.130 0.000 1299.410 4.000 ;
    END
  END la_data_in[106]
  PIN la_data_in[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1308.330 0.000 1308.610 4.000 ;
    END
  END la_data_in[107]
  PIN la_data_in[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1317.530 0.000 1317.810 4.000 ;
    END
  END la_data_in[108]
  PIN la_data_in[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1326.730 0.000 1327.010 4.000 ;
    END
  END la_data_in[109]
  PIN la_data_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 417.770 0.000 418.050 4.000 ;
    END
  END la_data_in[10]
  PIN la_data_in[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1335.930 0.000 1336.210 4.000 ;
    END
  END la_data_in[110]
  PIN la_data_in[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1345.130 0.000 1345.410 4.000 ;
    END
  END la_data_in[111]
  PIN la_data_in[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1354.330 0.000 1354.610 4.000 ;
    END
  END la_data_in[112]
  PIN la_data_in[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1363.530 0.000 1363.810 4.000 ;
    END
  END la_data_in[113]
  PIN la_data_in[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1372.730 0.000 1373.010 4.000 ;
    END
  END la_data_in[114]
  PIN la_data_in[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1381.930 0.000 1382.210 4.000 ;
    END
  END la_data_in[115]
  PIN la_data_in[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1391.130 0.000 1391.410 4.000 ;
    END
  END la_data_in[116]
  PIN la_data_in[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1400.330 0.000 1400.610 4.000 ;
    END
  END la_data_in[117]
  PIN la_data_in[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1409.530 0.000 1409.810 4.000 ;
    END
  END la_data_in[118]
  PIN la_data_in[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1418.730 0.000 1419.010 4.000 ;
    END
  END la_data_in[119]
  PIN la_data_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 426.970 0.000 427.250 4.000 ;
    END
  END la_data_in[11]
  PIN la_data_in[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1427.930 0.000 1428.210 4.000 ;
    END
  END la_data_in[120]
  PIN la_data_in[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1437.130 0.000 1437.410 4.000 ;
    END
  END la_data_in[121]
  PIN la_data_in[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1446.330 0.000 1446.610 4.000 ;
    END
  END la_data_in[122]
  PIN la_data_in[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1455.530 0.000 1455.810 4.000 ;
    END
  END la_data_in[123]
  PIN la_data_in[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1464.730 0.000 1465.010 4.000 ;
    END
  END la_data_in[124]
  PIN la_data_in[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1473.930 0.000 1474.210 4.000 ;
    END
  END la_data_in[125]
  PIN la_data_in[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1483.130 0.000 1483.410 4.000 ;
    END
  END la_data_in[126]
  PIN la_data_in[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1492.330 0.000 1492.610 4.000 ;
    END
  END la_data_in[127]
  PIN la_data_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 436.170 0.000 436.450 4.000 ;
    END
  END la_data_in[12]
  PIN la_data_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 444.910 0.000 445.190 4.000 ;
    END
  END la_data_in[13]
  PIN la_data_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 454.110 0.000 454.390 4.000 ;
    END
  END la_data_in[14]
  PIN la_data_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 463.310 0.000 463.590 4.000 ;
    END
  END la_data_in[15]
  PIN la_data_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 472.510 0.000 472.790 4.000 ;
    END
  END la_data_in[16]
  PIN la_data_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 481.710 0.000 481.990 4.000 ;
    END
  END la_data_in[17]
  PIN la_data_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 490.910 0.000 491.190 4.000 ;
    END
  END la_data_in[18]
  PIN la_data_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 500.110 0.000 500.390 4.000 ;
    END
  END la_data_in[19]
  PIN la_data_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 334.970 0.000 335.250 4.000 ;
    END
  END la_data_in[1]
  PIN la_data_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 509.310 0.000 509.590 4.000 ;
    END
  END la_data_in[20]
  PIN la_data_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END la_data_in[21]
  PIN la_data_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 527.710 0.000 527.990 4.000 ;
    END
  END la_data_in[22]
  PIN la_data_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 536.910 0.000 537.190 4.000 ;
    END
  END la_data_in[23]
  PIN la_data_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 546.110 0.000 546.390 4.000 ;
    END
  END la_data_in[24]
  PIN la_data_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 555.310 0.000 555.590 4.000 ;
    END
  END la_data_in[25]
  PIN la_data_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 564.510 0.000 564.790 4.000 ;
    END
  END la_data_in[26]
  PIN la_data_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 573.710 0.000 573.990 4.000 ;
    END
  END la_data_in[27]
  PIN la_data_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 582.910 0.000 583.190 4.000 ;
    END
  END la_data_in[28]
  PIN la_data_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 592.110 0.000 592.390 4.000 ;
    END
  END la_data_in[29]
  PIN la_data_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 344.170 0.000 344.450 4.000 ;
    END
  END la_data_in[2]
  PIN la_data_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 601.310 0.000 601.590 4.000 ;
    END
  END la_data_in[30]
  PIN la_data_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 610.510 0.000 610.790 4.000 ;
    END
  END la_data_in[31]
  PIN la_data_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 619.710 0.000 619.990 4.000 ;
    END
  END la_data_in[32]
  PIN la_data_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 628.910 0.000 629.190 4.000 ;
    END
  END la_data_in[33]
  PIN la_data_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 638.110 0.000 638.390 4.000 ;
    END
  END la_data_in[34]
  PIN la_data_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 647.310 0.000 647.590 4.000 ;
    END
  END la_data_in[35]
  PIN la_data_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 656.510 0.000 656.790 4.000 ;
    END
  END la_data_in[36]
  PIN la_data_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 665.710 0.000 665.990 4.000 ;
    END
  END la_data_in[37]
  PIN la_data_in[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 674.910 0.000 675.190 4.000 ;
    END
  END la_data_in[38]
  PIN la_data_in[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 684.110 0.000 684.390 4.000 ;
    END
  END la_data_in[39]
  PIN la_data_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 4.000 ;
    END
  END la_data_in[3]
  PIN la_data_in[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 693.310 0.000 693.590 4.000 ;
    END
  END la_data_in[40]
  PIN la_data_in[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 702.510 0.000 702.790 4.000 ;
    END
  END la_data_in[41]
  PIN la_data_in[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 711.250 0.000 711.530 4.000 ;
    END
  END la_data_in[42]
  PIN la_data_in[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 720.450 0.000 720.730 4.000 ;
    END
  END la_data_in[43]
  PIN la_data_in[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 729.650 0.000 729.930 4.000 ;
    END
  END la_data_in[44]
  PIN la_data_in[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 738.850 0.000 739.130 4.000 ;
    END
  END la_data_in[45]
  PIN la_data_in[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 748.050 0.000 748.330 4.000 ;
    END
  END la_data_in[46]
  PIN la_data_in[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.250 0.000 757.530 4.000 ;
    END
  END la_data_in[47]
  PIN la_data_in[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 766.450 0.000 766.730 4.000 ;
    END
  END la_data_in[48]
  PIN la_data_in[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 775.650 0.000 775.930 4.000 ;
    END
  END la_data_in[49]
  PIN la_data_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 362.570 0.000 362.850 4.000 ;
    END
  END la_data_in[4]
  PIN la_data_in[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 784.850 0.000 785.130 4.000 ;
    END
  END la_data_in[50]
  PIN la_data_in[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 794.050 0.000 794.330 4.000 ;
    END
  END la_data_in[51]
  PIN la_data_in[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 803.250 0.000 803.530 4.000 ;
    END
  END la_data_in[52]
  PIN la_data_in[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 812.450 0.000 812.730 4.000 ;
    END
  END la_data_in[53]
  PIN la_data_in[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 821.650 0.000 821.930 4.000 ;
    END
  END la_data_in[54]
  PIN la_data_in[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 830.850 0.000 831.130 4.000 ;
    END
  END la_data_in[55]
  PIN la_data_in[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 840.050 0.000 840.330 4.000 ;
    END
  END la_data_in[56]
  PIN la_data_in[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 849.250 0.000 849.530 4.000 ;
    END
  END la_data_in[57]
  PIN la_data_in[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 858.450 0.000 858.730 4.000 ;
    END
  END la_data_in[58]
  PIN la_data_in[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 867.650 0.000 867.930 4.000 ;
    END
  END la_data_in[59]
  PIN la_data_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 371.770 0.000 372.050 4.000 ;
    END
  END la_data_in[5]
  PIN la_data_in[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.850 0.000 877.130 4.000 ;
    END
  END la_data_in[60]
  PIN la_data_in[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 886.050 0.000 886.330 4.000 ;
    END
  END la_data_in[61]
  PIN la_data_in[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 895.250 0.000 895.530 4.000 ;
    END
  END la_data_in[62]
  PIN la_data_in[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 904.450 0.000 904.730 4.000 ;
    END
  END la_data_in[63]
  PIN la_data_in[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 913.650 0.000 913.930 4.000 ;
    END
  END la_data_in[64]
  PIN la_data_in[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 922.850 0.000 923.130 4.000 ;
    END
  END la_data_in[65]
  PIN la_data_in[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 932.050 0.000 932.330 4.000 ;
    END
  END la_data_in[66]
  PIN la_data_in[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 941.250 0.000 941.530 4.000 ;
    END
  END la_data_in[67]
  PIN la_data_in[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 950.450 0.000 950.730 4.000 ;
    END
  END la_data_in[68]
  PIN la_data_in[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 959.650 0.000 959.930 4.000 ;
    END
  END la_data_in[69]
  PIN la_data_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 380.970 0.000 381.250 4.000 ;
    END
  END la_data_in[6]
  PIN la_data_in[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 968.850 0.000 969.130 4.000 ;
    END
  END la_data_in[70]
  PIN la_data_in[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 977.590 0.000 977.870 4.000 ;
    END
  END la_data_in[71]
  PIN la_data_in[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 986.790 0.000 987.070 4.000 ;
    END
  END la_data_in[72]
  PIN la_data_in[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 995.990 0.000 996.270 4.000 ;
    END
  END la_data_in[73]
  PIN la_data_in[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1005.190 0.000 1005.470 4.000 ;
    END
  END la_data_in[74]
  PIN la_data_in[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1014.390 0.000 1014.670 4.000 ;
    END
  END la_data_in[75]
  PIN la_data_in[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1023.590 0.000 1023.870 4.000 ;
    END
  END la_data_in[76]
  PIN la_data_in[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1032.790 0.000 1033.070 4.000 ;
    END
  END la_data_in[77]
  PIN la_data_in[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1041.990 0.000 1042.270 4.000 ;
    END
  END la_data_in[78]
  PIN la_data_in[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1051.190 0.000 1051.470 4.000 ;
    END
  END la_data_in[79]
  PIN la_data_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 390.170 0.000 390.450 4.000 ;
    END
  END la_data_in[7]
  PIN la_data_in[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1060.390 0.000 1060.670 4.000 ;
    END
  END la_data_in[80]
  PIN la_data_in[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1069.590 0.000 1069.870 4.000 ;
    END
  END la_data_in[81]
  PIN la_data_in[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1078.790 0.000 1079.070 4.000 ;
    END
  END la_data_in[82]
  PIN la_data_in[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1087.990 0.000 1088.270 4.000 ;
    END
  END la_data_in[83]
  PIN la_data_in[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1097.190 0.000 1097.470 4.000 ;
    END
  END la_data_in[84]
  PIN la_data_in[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1106.390 0.000 1106.670 4.000 ;
    END
  END la_data_in[85]
  PIN la_data_in[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1115.590 0.000 1115.870 4.000 ;
    END
  END la_data_in[86]
  PIN la_data_in[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1124.790 0.000 1125.070 4.000 ;
    END
  END la_data_in[87]
  PIN la_data_in[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1133.990 0.000 1134.270 4.000 ;
    END
  END la_data_in[88]
  PIN la_data_in[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1143.190 0.000 1143.470 4.000 ;
    END
  END la_data_in[89]
  PIN la_data_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END la_data_in[8]
  PIN la_data_in[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1152.390 0.000 1152.670 4.000 ;
    END
  END la_data_in[90]
  PIN la_data_in[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1161.590 0.000 1161.870 4.000 ;
    END
  END la_data_in[91]
  PIN la_data_in[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1170.790 0.000 1171.070 4.000 ;
    END
  END la_data_in[92]
  PIN la_data_in[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1179.990 0.000 1180.270 4.000 ;
    END
  END la_data_in[93]
  PIN la_data_in[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1189.190 0.000 1189.470 4.000 ;
    END
  END la_data_in[94]
  PIN la_data_in[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1198.390 0.000 1198.670 4.000 ;
    END
  END la_data_in[95]
  PIN la_data_in[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1207.590 0.000 1207.870 4.000 ;
    END
  END la_data_in[96]
  PIN la_data_in[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1216.790 0.000 1217.070 4.000 ;
    END
  END la_data_in[97]
  PIN la_data_in[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1225.990 0.000 1226.270 4.000 ;
    END
  END la_data_in[98]
  PIN la_data_in[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1235.190 0.000 1235.470 4.000 ;
    END
  END la_data_in[99]
  PIN la_data_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 408.570 0.000 408.850 4.000 ;
    END
  END la_data_in[9]
  PIN la_data_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 328.990 0.000 329.270 4.000 ;
    END
  END la_data_out[0]
  PIN la_data_out[100]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1247.150 0.000 1247.430 4.000 ;
    END
  END la_data_out[100]
  PIN la_data_out[101]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1256.350 0.000 1256.630 4.000 ;
    END
  END la_data_out[101]
  PIN la_data_out[102]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1265.550 0.000 1265.830 4.000 ;
    END
  END la_data_out[102]
  PIN la_data_out[103]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1274.750 0.000 1275.030 4.000 ;
    END
  END la_data_out[103]
  PIN la_data_out[104]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1283.950 0.000 1284.230 4.000 ;
    END
  END la_data_out[104]
  PIN la_data_out[105]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1293.150 0.000 1293.430 4.000 ;
    END
  END la_data_out[105]
  PIN la_data_out[106]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1302.350 0.000 1302.630 4.000 ;
    END
  END la_data_out[106]
  PIN la_data_out[107]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1311.550 0.000 1311.830 4.000 ;
    END
  END la_data_out[107]
  PIN la_data_out[108]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1320.750 0.000 1321.030 4.000 ;
    END
  END la_data_out[108]
  PIN la_data_out[109]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1329.950 0.000 1330.230 4.000 ;
    END
  END la_data_out[109]
  PIN la_data_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 420.530 0.000 420.810 4.000 ;
    END
  END la_data_out[10]
  PIN la_data_out[110]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1339.150 0.000 1339.430 4.000 ;
    END
  END la_data_out[110]
  PIN la_data_out[111]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1348.350 0.000 1348.630 4.000 ;
    END
  END la_data_out[111]
  PIN la_data_out[112]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1357.550 0.000 1357.830 4.000 ;
    END
  END la_data_out[112]
  PIN la_data_out[113]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1366.750 0.000 1367.030 4.000 ;
    END
  END la_data_out[113]
  PIN la_data_out[114]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1375.950 0.000 1376.230 4.000 ;
    END
  END la_data_out[114]
  PIN la_data_out[115]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1385.150 0.000 1385.430 4.000 ;
    END
  END la_data_out[115]
  PIN la_data_out[116]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1394.350 0.000 1394.630 4.000 ;
    END
  END la_data_out[116]
  PIN la_data_out[117]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1403.550 0.000 1403.830 4.000 ;
    END
  END la_data_out[117]
  PIN la_data_out[118]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1412.750 0.000 1413.030 4.000 ;
    END
  END la_data_out[118]
  PIN la_data_out[119]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1421.490 0.000 1421.770 4.000 ;
    END
  END la_data_out[119]
  PIN la_data_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 429.730 0.000 430.010 4.000 ;
    END
  END la_data_out[11]
  PIN la_data_out[120]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1430.690 0.000 1430.970 4.000 ;
    END
  END la_data_out[120]
  PIN la_data_out[121]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1439.890 0.000 1440.170 4.000 ;
    END
  END la_data_out[121]
  PIN la_data_out[122]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1449.090 0.000 1449.370 4.000 ;
    END
  END la_data_out[122]
  PIN la_data_out[123]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1458.290 0.000 1458.570 4.000 ;
    END
  END la_data_out[123]
  PIN la_data_out[124]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1467.490 0.000 1467.770 4.000 ;
    END
  END la_data_out[124]
  PIN la_data_out[125]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1476.690 0.000 1476.970 4.000 ;
    END
  END la_data_out[125]
  PIN la_data_out[126]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1485.890 0.000 1486.170 4.000 ;
    END
  END la_data_out[126]
  PIN la_data_out[127]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1495.090 0.000 1495.370 4.000 ;
    END
  END la_data_out[127]
  PIN la_data_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 438.930 0.000 439.210 4.000 ;
    END
  END la_data_out[12]
  PIN la_data_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 448.130 0.000 448.410 4.000 ;
    END
  END la_data_out[13]
  PIN la_data_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END la_data_out[14]
  PIN la_data_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 466.530 0.000 466.810 4.000 ;
    END
  END la_data_out[15]
  PIN la_data_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 475.730 0.000 476.010 4.000 ;
    END
  END la_data_out[16]
  PIN la_data_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 484.930 0.000 485.210 4.000 ;
    END
  END la_data_out[17]
  PIN la_data_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 494.130 0.000 494.410 4.000 ;
    END
  END la_data_out[18]
  PIN la_data_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 503.330 0.000 503.610 4.000 ;
    END
  END la_data_out[19]
  PIN la_data_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END la_data_out[1]
  PIN la_data_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 512.530 0.000 512.810 4.000 ;
    END
  END la_data_out[20]
  PIN la_data_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 521.730 0.000 522.010 4.000 ;
    END
  END la_data_out[21]
  PIN la_data_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 530.930 0.000 531.210 4.000 ;
    END
  END la_data_out[22]
  PIN la_data_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 540.130 0.000 540.410 4.000 ;
    END
  END la_data_out[23]
  PIN la_data_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 549.330 0.000 549.610 4.000 ;
    END
  END la_data_out[24]
  PIN la_data_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 558.530 0.000 558.810 4.000 ;
    END
  END la_data_out[25]
  PIN la_data_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 567.730 0.000 568.010 4.000 ;
    END
  END la_data_out[26]
  PIN la_data_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 576.930 0.000 577.210 4.000 ;
    END
  END la_data_out[27]
  PIN la_data_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 586.130 0.000 586.410 4.000 ;
    END
  END la_data_out[28]
  PIN la_data_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 595.330 0.000 595.610 4.000 ;
    END
  END la_data_out[29]
  PIN la_data_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 347.390 0.000 347.670 4.000 ;
    END
  END la_data_out[2]
  PIN la_data_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 604.530 0.000 604.810 4.000 ;
    END
  END la_data_out[30]
  PIN la_data_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 613.730 0.000 614.010 4.000 ;
    END
  END la_data_out[31]
  PIN la_data_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 622.470 0.000 622.750 4.000 ;
    END
  END la_data_out[32]
  PIN la_data_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 631.670 0.000 631.950 4.000 ;
    END
  END la_data_out[33]
  PIN la_data_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 640.870 0.000 641.150 4.000 ;
    END
  END la_data_out[34]
  PIN la_data_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 650.070 0.000 650.350 4.000 ;
    END
  END la_data_out[35]
  PIN la_data_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 659.270 0.000 659.550 4.000 ;
    END
  END la_data_out[36]
  PIN la_data_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 668.470 0.000 668.750 4.000 ;
    END
  END la_data_out[37]
  PIN la_data_out[38]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 677.670 0.000 677.950 4.000 ;
    END
  END la_data_out[38]
  PIN la_data_out[39]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 686.870 0.000 687.150 4.000 ;
    END
  END la_data_out[39]
  PIN la_data_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 356.130 0.000 356.410 4.000 ;
    END
  END la_data_out[3]
  PIN la_data_out[40]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 696.070 0.000 696.350 4.000 ;
    END
  END la_data_out[40]
  PIN la_data_out[41]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 705.270 0.000 705.550 4.000 ;
    END
  END la_data_out[41]
  PIN la_data_out[42]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 714.470 0.000 714.750 4.000 ;
    END
  END la_data_out[42]
  PIN la_data_out[43]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 723.670 0.000 723.950 4.000 ;
    END
  END la_data_out[43]
  PIN la_data_out[44]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 732.870 0.000 733.150 4.000 ;
    END
  END la_data_out[44]
  PIN la_data_out[45]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 742.070 0.000 742.350 4.000 ;
    END
  END la_data_out[45]
  PIN la_data_out[46]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 751.270 0.000 751.550 4.000 ;
    END
  END la_data_out[46]
  PIN la_data_out[47]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 760.470 0.000 760.750 4.000 ;
    END
  END la_data_out[47]
  PIN la_data_out[48]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 769.670 0.000 769.950 4.000 ;
    END
  END la_data_out[48]
  PIN la_data_out[49]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 778.870 0.000 779.150 4.000 ;
    END
  END la_data_out[49]
  PIN la_data_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 365.330 0.000 365.610 4.000 ;
    END
  END la_data_out[4]
  PIN la_data_out[50]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 788.070 0.000 788.350 4.000 ;
    END
  END la_data_out[50]
  PIN la_data_out[51]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 797.270 0.000 797.550 4.000 ;
    END
  END la_data_out[51]
  PIN la_data_out[52]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 806.470 0.000 806.750 4.000 ;
    END
  END la_data_out[52]
  PIN la_data_out[53]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 815.670 0.000 815.950 4.000 ;
    END
  END la_data_out[53]
  PIN la_data_out[54]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 824.870 0.000 825.150 4.000 ;
    END
  END la_data_out[54]
  PIN la_data_out[55]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 834.070 0.000 834.350 4.000 ;
    END
  END la_data_out[55]
  PIN la_data_out[56]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 843.270 0.000 843.550 4.000 ;
    END
  END la_data_out[56]
  PIN la_data_out[57]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 852.470 0.000 852.750 4.000 ;
    END
  END la_data_out[57]
  PIN la_data_out[58]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 861.670 0.000 861.950 4.000 ;
    END
  END la_data_out[58]
  PIN la_data_out[59]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 870.870 0.000 871.150 4.000 ;
    END
  END la_data_out[59]
  PIN la_data_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END la_data_out[5]
  PIN la_data_out[60]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 880.070 0.000 880.350 4.000 ;
    END
  END la_data_out[60]
  PIN la_data_out[61]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 888.810 0.000 889.090 4.000 ;
    END
  END la_data_out[61]
  PIN la_data_out[62]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 898.010 0.000 898.290 4.000 ;
    END
  END la_data_out[62]
  PIN la_data_out[63]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 907.210 0.000 907.490 4.000 ;
    END
  END la_data_out[63]
  PIN la_data_out[64]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 916.410 0.000 916.690 4.000 ;
    END
  END la_data_out[64]
  PIN la_data_out[65]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 925.610 0.000 925.890 4.000 ;
    END
  END la_data_out[65]
  PIN la_data_out[66]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 934.810 0.000 935.090 4.000 ;
    END
  END la_data_out[66]
  PIN la_data_out[67]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 944.010 0.000 944.290 4.000 ;
    END
  END la_data_out[67]
  PIN la_data_out[68]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 953.210 0.000 953.490 4.000 ;
    END
  END la_data_out[68]
  PIN la_data_out[69]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 962.410 0.000 962.690 4.000 ;
    END
  END la_data_out[69]
  PIN la_data_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 383.730 0.000 384.010 4.000 ;
    END
  END la_data_out[6]
  PIN la_data_out[70]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 971.610 0.000 971.890 4.000 ;
    END
  END la_data_out[70]
  PIN la_data_out[71]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 980.810 0.000 981.090 4.000 ;
    END
  END la_data_out[71]
  PIN la_data_out[72]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 990.010 0.000 990.290 4.000 ;
    END
  END la_data_out[72]
  PIN la_data_out[73]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 999.210 0.000 999.490 4.000 ;
    END
  END la_data_out[73]
  PIN la_data_out[74]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1008.410 0.000 1008.690 4.000 ;
    END
  END la_data_out[74]
  PIN la_data_out[75]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1017.610 0.000 1017.890 4.000 ;
    END
  END la_data_out[75]
  PIN la_data_out[76]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1026.810 0.000 1027.090 4.000 ;
    END
  END la_data_out[76]
  PIN la_data_out[77]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1036.010 0.000 1036.290 4.000 ;
    END
  END la_data_out[77]
  PIN la_data_out[78]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1045.210 0.000 1045.490 4.000 ;
    END
  END la_data_out[78]
  PIN la_data_out[79]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1054.410 0.000 1054.690 4.000 ;
    END
  END la_data_out[79]
  PIN la_data_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END la_data_out[7]
  PIN la_data_out[80]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1063.610 0.000 1063.890 4.000 ;
    END
  END la_data_out[80]
  PIN la_data_out[81]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1072.810 0.000 1073.090 4.000 ;
    END
  END la_data_out[81]
  PIN la_data_out[82]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1082.010 0.000 1082.290 4.000 ;
    END
  END la_data_out[82]
  PIN la_data_out[83]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1091.210 0.000 1091.490 4.000 ;
    END
  END la_data_out[83]
  PIN la_data_out[84]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1100.410 0.000 1100.690 4.000 ;
    END
  END la_data_out[84]
  PIN la_data_out[85]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1109.610 0.000 1109.890 4.000 ;
    END
  END la_data_out[85]
  PIN la_data_out[86]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1118.810 0.000 1119.090 4.000 ;
    END
  END la_data_out[86]
  PIN la_data_out[87]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1128.010 0.000 1128.290 4.000 ;
    END
  END la_data_out[87]
  PIN la_data_out[88]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1137.210 0.000 1137.490 4.000 ;
    END
  END la_data_out[88]
  PIN la_data_out[89]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1146.410 0.000 1146.690 4.000 ;
    END
  END la_data_out[89]
  PIN la_data_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 402.130 0.000 402.410 4.000 ;
    END
  END la_data_out[8]
  PIN la_data_out[90]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1155.150 0.000 1155.430 4.000 ;
    END
  END la_data_out[90]
  PIN la_data_out[91]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1164.350 0.000 1164.630 4.000 ;
    END
  END la_data_out[91]
  PIN la_data_out[92]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1173.550 0.000 1173.830 4.000 ;
    END
  END la_data_out[92]
  PIN la_data_out[93]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1182.750 0.000 1183.030 4.000 ;
    END
  END la_data_out[93]
  PIN la_data_out[94]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1191.950 0.000 1192.230 4.000 ;
    END
  END la_data_out[94]
  PIN la_data_out[95]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1201.150 0.000 1201.430 4.000 ;
    END
  END la_data_out[95]
  PIN la_data_out[96]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1210.350 0.000 1210.630 4.000 ;
    END
  END la_data_out[96]
  PIN la_data_out[97]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1219.550 0.000 1219.830 4.000 ;
    END
  END la_data_out[97]
  PIN la_data_out[98]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1228.750 0.000 1229.030 4.000 ;
    END
  END la_data_out[98]
  PIN la_data_out[99]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1237.950 0.000 1238.230 4.000 ;
    END
  END la_data_out[99]
  PIN la_data_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 411.330 0.000 411.610 4.000 ;
    END
  END la_data_out[9]
  PIN la_oen[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END la_oen[0]
  PIN la_oen[100]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1250.370 0.000 1250.650 4.000 ;
    END
  END la_oen[100]
  PIN la_oen[101]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1259.570 0.000 1259.850 4.000 ;
    END
  END la_oen[101]
  PIN la_oen[102]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1268.770 0.000 1269.050 4.000 ;
    END
  END la_oen[102]
  PIN la_oen[103]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1277.970 0.000 1278.250 4.000 ;
    END
  END la_oen[103]
  PIN la_oen[104]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1287.170 0.000 1287.450 4.000 ;
    END
  END la_oen[104]
  PIN la_oen[105]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1296.370 0.000 1296.650 4.000 ;
    END
  END la_oen[105]
  PIN la_oen[106]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1305.570 0.000 1305.850 4.000 ;
    END
  END la_oen[106]
  PIN la_oen[107]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1314.770 0.000 1315.050 4.000 ;
    END
  END la_oen[107]
  PIN la_oen[108]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1323.970 0.000 1324.250 4.000 ;
    END
  END la_oen[108]
  PIN la_oen[109]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1332.710 0.000 1332.990 4.000 ;
    END
  END la_oen[109]
  PIN la_oen[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 423.750 0.000 424.030 4.000 ;
    END
  END la_oen[10]
  PIN la_oen[110]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1341.910 0.000 1342.190 4.000 ;
    END
  END la_oen[110]
  PIN la_oen[111]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1351.110 0.000 1351.390 4.000 ;
    END
  END la_oen[111]
  PIN la_oen[112]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1360.310 0.000 1360.590 4.000 ;
    END
  END la_oen[112]
  PIN la_oen[113]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1369.510 0.000 1369.790 4.000 ;
    END
  END la_oen[113]
  PIN la_oen[114]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1378.710 0.000 1378.990 4.000 ;
    END
  END la_oen[114]
  PIN la_oen[115]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1387.910 0.000 1388.190 4.000 ;
    END
  END la_oen[115]
  PIN la_oen[116]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1397.110 0.000 1397.390 4.000 ;
    END
  END la_oen[116]
  PIN la_oen[117]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1406.310 0.000 1406.590 4.000 ;
    END
  END la_oen[117]
  PIN la_oen[118]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1415.510 0.000 1415.790 4.000 ;
    END
  END la_oen[118]
  PIN la_oen[119]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1424.710 0.000 1424.990 4.000 ;
    END
  END la_oen[119]
  PIN la_oen[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 432.950 0.000 433.230 4.000 ;
    END
  END la_oen[11]
  PIN la_oen[120]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1433.910 0.000 1434.190 4.000 ;
    END
  END la_oen[120]
  PIN la_oen[121]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1443.110 0.000 1443.390 4.000 ;
    END
  END la_oen[121]
  PIN la_oen[122]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1452.310 0.000 1452.590 4.000 ;
    END
  END la_oen[122]
  PIN la_oen[123]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1461.510 0.000 1461.790 4.000 ;
    END
  END la_oen[123]
  PIN la_oen[124]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1470.710 0.000 1470.990 4.000 ;
    END
  END la_oen[124]
  PIN la_oen[125]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1479.910 0.000 1480.190 4.000 ;
    END
  END la_oen[125]
  PIN la_oen[126]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1489.110 0.000 1489.390 4.000 ;
    END
  END la_oen[126]
  PIN la_oen[127]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1498.310 0.000 1498.590 4.000 ;
    END
  END la_oen[127]
  PIN la_oen[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 442.150 0.000 442.430 4.000 ;
    END
  END la_oen[12]
  PIN la_oen[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 451.350 0.000 451.630 4.000 ;
    END
  END la_oen[13]
  PIN la_oen[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END la_oen[14]
  PIN la_oen[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 469.750 0.000 470.030 4.000 ;
    END
  END la_oen[15]
  PIN la_oen[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 478.950 0.000 479.230 4.000 ;
    END
  END la_oen[16]
  PIN la_oen[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 488.150 0.000 488.430 4.000 ;
    END
  END la_oen[17]
  PIN la_oen[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 497.350 0.000 497.630 4.000 ;
    END
  END la_oen[18]
  PIN la_oen[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 506.550 0.000 506.830 4.000 ;
    END
  END la_oen[19]
  PIN la_oen[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 340.950 0.000 341.230 4.000 ;
    END
  END la_oen[1]
  PIN la_oen[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 515.750 0.000 516.030 4.000 ;
    END
  END la_oen[20]
  PIN la_oen[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END la_oen[21]
  PIN la_oen[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 533.690 0.000 533.970 4.000 ;
    END
  END la_oen[22]
  PIN la_oen[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 542.890 0.000 543.170 4.000 ;
    END
  END la_oen[23]
  PIN la_oen[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 552.090 0.000 552.370 4.000 ;
    END
  END la_oen[24]
  PIN la_oen[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 561.290 0.000 561.570 4.000 ;
    END
  END la_oen[25]
  PIN la_oen[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 570.490 0.000 570.770 4.000 ;
    END
  END la_oen[26]
  PIN la_oen[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END la_oen[27]
  PIN la_oen[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 588.890 0.000 589.170 4.000 ;
    END
  END la_oen[28]
  PIN la_oen[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 598.090 0.000 598.370 4.000 ;
    END
  END la_oen[29]
  PIN la_oen[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 350.150 0.000 350.430 4.000 ;
    END
  END la_oen[2]
  PIN la_oen[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 607.290 0.000 607.570 4.000 ;
    END
  END la_oen[30]
  PIN la_oen[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 616.490 0.000 616.770 4.000 ;
    END
  END la_oen[31]
  PIN la_oen[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 625.690 0.000 625.970 4.000 ;
    END
  END la_oen[32]
  PIN la_oen[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 634.890 0.000 635.170 4.000 ;
    END
  END la_oen[33]
  PIN la_oen[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 644.090 0.000 644.370 4.000 ;
    END
  END la_oen[34]
  PIN la_oen[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 653.290 0.000 653.570 4.000 ;
    END
  END la_oen[35]
  PIN la_oen[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 662.490 0.000 662.770 4.000 ;
    END
  END la_oen[36]
  PIN la_oen[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 671.690 0.000 671.970 4.000 ;
    END
  END la_oen[37]
  PIN la_oen[38]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 680.890 0.000 681.170 4.000 ;
    END
  END la_oen[38]
  PIN la_oen[39]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 690.090 0.000 690.370 4.000 ;
    END
  END la_oen[39]
  PIN la_oen[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 359.350 0.000 359.630 4.000 ;
    END
  END la_oen[3]
  PIN la_oen[40]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 699.290 0.000 699.570 4.000 ;
    END
  END la_oen[40]
  PIN la_oen[41]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 708.490 0.000 708.770 4.000 ;
    END
  END la_oen[41]
  PIN la_oen[42]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 717.690 0.000 717.970 4.000 ;
    END
  END la_oen[42]
  PIN la_oen[43]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 726.890 0.000 727.170 4.000 ;
    END
  END la_oen[43]
  PIN la_oen[44]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 736.090 0.000 736.370 4.000 ;
    END
  END la_oen[44]
  PIN la_oen[45]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 745.290 0.000 745.570 4.000 ;
    END
  END la_oen[45]
  PIN la_oen[46]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 754.490 0.000 754.770 4.000 ;
    END
  END la_oen[46]
  PIN la_oen[47]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 763.690 0.000 763.970 4.000 ;
    END
  END la_oen[47]
  PIN la_oen[48]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 772.890 0.000 773.170 4.000 ;
    END
  END la_oen[48]
  PIN la_oen[49]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 782.090 0.000 782.370 4.000 ;
    END
  END la_oen[49]
  PIN la_oen[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 368.550 0.000 368.830 4.000 ;
    END
  END la_oen[4]
  PIN la_oen[50]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 791.290 0.000 791.570 4.000 ;
    END
  END la_oen[50]
  PIN la_oen[51]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 800.030 0.000 800.310 4.000 ;
    END
  END la_oen[51]
  PIN la_oen[52]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 809.230 0.000 809.510 4.000 ;
    END
  END la_oen[52]
  PIN la_oen[53]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 818.430 0.000 818.710 4.000 ;
    END
  END la_oen[53]
  PIN la_oen[54]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 827.630 0.000 827.910 4.000 ;
    END
  END la_oen[54]
  PIN la_oen[55]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 836.830 0.000 837.110 4.000 ;
    END
  END la_oen[55]
  PIN la_oen[56]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.030 0.000 846.310 4.000 ;
    END
  END la_oen[56]
  PIN la_oen[57]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 855.230 0.000 855.510 4.000 ;
    END
  END la_oen[57]
  PIN la_oen[58]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 864.430 0.000 864.710 4.000 ;
    END
  END la_oen[58]
  PIN la_oen[59]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 873.630 0.000 873.910 4.000 ;
    END
  END la_oen[59]
  PIN la_oen[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 377.750 0.000 378.030 4.000 ;
    END
  END la_oen[5]
  PIN la_oen[60]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 882.830 0.000 883.110 4.000 ;
    END
  END la_oen[60]
  PIN la_oen[61]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 892.030 0.000 892.310 4.000 ;
    END
  END la_oen[61]
  PIN la_oen[62]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 901.230 0.000 901.510 4.000 ;
    END
  END la_oen[62]
  PIN la_oen[63]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 910.430 0.000 910.710 4.000 ;
    END
  END la_oen[63]
  PIN la_oen[64]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 919.630 0.000 919.910 4.000 ;
    END
  END la_oen[64]
  PIN la_oen[65]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 928.830 0.000 929.110 4.000 ;
    END
  END la_oen[65]
  PIN la_oen[66]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 938.030 0.000 938.310 4.000 ;
    END
  END la_oen[66]
  PIN la_oen[67]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 947.230 0.000 947.510 4.000 ;
    END
  END la_oen[67]
  PIN la_oen[68]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 956.430 0.000 956.710 4.000 ;
    END
  END la_oen[68]
  PIN la_oen[69]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 965.630 0.000 965.910 4.000 ;
    END
  END la_oen[69]
  PIN la_oen[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 386.950 0.000 387.230 4.000 ;
    END
  END la_oen[6]
  PIN la_oen[70]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 974.830 0.000 975.110 4.000 ;
    END
  END la_oen[70]
  PIN la_oen[71]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 984.030 0.000 984.310 4.000 ;
    END
  END la_oen[71]
  PIN la_oen[72]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 993.230 0.000 993.510 4.000 ;
    END
  END la_oen[72]
  PIN la_oen[73]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1002.430 0.000 1002.710 4.000 ;
    END
  END la_oen[73]
  PIN la_oen[74]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1011.630 0.000 1011.910 4.000 ;
    END
  END la_oen[74]
  PIN la_oen[75]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1020.830 0.000 1021.110 4.000 ;
    END
  END la_oen[75]
  PIN la_oen[76]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1030.030 0.000 1030.310 4.000 ;
    END
  END la_oen[76]
  PIN la_oen[77]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1039.230 0.000 1039.510 4.000 ;
    END
  END la_oen[77]
  PIN la_oen[78]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1048.430 0.000 1048.710 4.000 ;
    END
  END la_oen[78]
  PIN la_oen[79]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1057.630 0.000 1057.910 4.000 ;
    END
  END la_oen[79]
  PIN la_oen[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 396.150 0.000 396.430 4.000 ;
    END
  END la_oen[7]
  PIN la_oen[80]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1066.370 0.000 1066.650 4.000 ;
    END
  END la_oen[80]
  PIN la_oen[81]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1075.570 0.000 1075.850 4.000 ;
    END
  END la_oen[81]
  PIN la_oen[82]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1084.770 0.000 1085.050 4.000 ;
    END
  END la_oen[82]
  PIN la_oen[83]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1093.970 0.000 1094.250 4.000 ;
    END
  END la_oen[83]
  PIN la_oen[84]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1103.170 0.000 1103.450 4.000 ;
    END
  END la_oen[84]
  PIN la_oen[85]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1112.370 0.000 1112.650 4.000 ;
    END
  END la_oen[85]
  PIN la_oen[86]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1121.570 0.000 1121.850 4.000 ;
    END
  END la_oen[86]
  PIN la_oen[87]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1130.770 0.000 1131.050 4.000 ;
    END
  END la_oen[87]
  PIN la_oen[88]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1139.970 0.000 1140.250 4.000 ;
    END
  END la_oen[88]
  PIN la_oen[89]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1149.170 0.000 1149.450 4.000 ;
    END
  END la_oen[89]
  PIN la_oen[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 405.350 0.000 405.630 4.000 ;
    END
  END la_oen[8]
  PIN la_oen[90]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1158.370 0.000 1158.650 4.000 ;
    END
  END la_oen[90]
  PIN la_oen[91]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1167.570 0.000 1167.850 4.000 ;
    END
  END la_oen[91]
  PIN la_oen[92]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1176.770 0.000 1177.050 4.000 ;
    END
  END la_oen[92]
  PIN la_oen[93]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.970 0.000 1186.250 4.000 ;
    END
  END la_oen[93]
  PIN la_oen[94]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1195.170 0.000 1195.450 4.000 ;
    END
  END la_oen[94]
  PIN la_oen[95]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1204.370 0.000 1204.650 4.000 ;
    END
  END la_oen[95]
  PIN la_oen[96]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1213.570 0.000 1213.850 4.000 ;
    END
  END la_oen[96]
  PIN la_oen[97]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1222.770 0.000 1223.050 4.000 ;
    END
  END la_oen[97]
  PIN la_oen[98]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1231.970 0.000 1232.250 4.000 ;
    END
  END la_oen[98]
  PIN la_oen[99]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1241.170 0.000 1241.450 4.000 ;
    END
  END la_oen[99]
  PIN la_oen[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 414.550 0.000 414.830 4.000 ;
    END
  END la_oen[9]
  PIN proj0_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 172.590 396.000 172.870 400.000 ;
    END
  END proj0_clk
  PIN proj0_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 179.030 396.000 179.310 400.000 ;
    END
  END proj0_io_in[0]
  PIN proj0_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 222.730 396.000 223.010 400.000 ;
    END
  END proj0_io_in[10]
  PIN proj0_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 226.870 396.000 227.150 400.000 ;
    END
  END proj0_io_in[11]
  PIN proj0_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 231.010 396.000 231.290 400.000 ;
    END
  END proj0_io_in[12]
  PIN proj0_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 235.610 396.000 235.890 400.000 ;
    END
  END proj0_io_in[13]
  PIN proj0_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 239.750 396.000 240.030 400.000 ;
    END
  END proj0_io_in[14]
  PIN proj0_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 244.350 396.000 244.630 400.000 ;
    END
  END proj0_io_in[15]
  PIN proj0_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 248.490 396.000 248.770 400.000 ;
    END
  END proj0_io_in[16]
  PIN proj0_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 253.090 396.000 253.370 400.000 ;
    END
  END proj0_io_in[17]
  PIN proj0_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 257.230 396.000 257.510 400.000 ;
    END
  END proj0_io_in[18]
  PIN proj0_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 261.830 396.000 262.110 400.000 ;
    END
  END proj0_io_in[19]
  PIN proj0_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 183.170 396.000 183.450 400.000 ;
    END
  END proj0_io_in[1]
  PIN proj0_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 265.970 396.000 266.250 400.000 ;
    END
  END proj0_io_in[20]
  PIN proj0_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 270.570 396.000 270.850 400.000 ;
    END
  END proj0_io_in[21]
  PIN proj0_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 274.710 396.000 274.990 400.000 ;
    END
  END proj0_io_in[22]
  PIN proj0_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 278.850 396.000 279.130 400.000 ;
    END
  END proj0_io_in[23]
  PIN proj0_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 283.450 396.000 283.730 400.000 ;
    END
  END proj0_io_in[24]
  PIN proj0_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 287.590 396.000 287.870 400.000 ;
    END
  END proj0_io_in[25]
  PIN proj0_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 292.190 396.000 292.470 400.000 ;
    END
  END proj0_io_in[26]
  PIN proj0_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 296.330 396.000 296.610 400.000 ;
    END
  END proj0_io_in[27]
  PIN proj0_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 300.930 396.000 301.210 400.000 ;
    END
  END proj0_io_in[28]
  PIN proj0_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 305.070 396.000 305.350 400.000 ;
    END
  END proj0_io_in[29]
  PIN proj0_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 187.770 396.000 188.050 400.000 ;
    END
  END proj0_io_in[2]
  PIN proj0_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 309.670 396.000 309.950 400.000 ;
    END
  END proj0_io_in[30]
  PIN proj0_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 313.810 396.000 314.090 400.000 ;
    END
  END proj0_io_in[31]
  PIN proj0_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 318.410 396.000 318.690 400.000 ;
    END
  END proj0_io_in[32]
  PIN proj0_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 322.550 396.000 322.830 400.000 ;
    END
  END proj0_io_in[33]
  PIN proj0_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 326.690 396.000 326.970 400.000 ;
    END
  END proj0_io_in[34]
  PIN proj0_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 331.290 396.000 331.570 400.000 ;
    END
  END proj0_io_in[35]
  PIN proj0_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 335.430 396.000 335.710 400.000 ;
    END
  END proj0_io_in[36]
  PIN proj0_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 340.030 396.000 340.310 400.000 ;
    END
  END proj0_io_in[37]
  PIN proj0_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 191.910 396.000 192.190 400.000 ;
    END
  END proj0_io_in[3]
  PIN proj0_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 196.510 396.000 196.790 400.000 ;
    END
  END proj0_io_in[4]
  PIN proj0_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 200.650 396.000 200.930 400.000 ;
    END
  END proj0_io_in[5]
  PIN proj0_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 205.250 396.000 205.530 400.000 ;
    END
  END proj0_io_in[6]
  PIN proj0_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 209.390 396.000 209.670 400.000 ;
    END
  END proj0_io_in[7]
  PIN proj0_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 213.990 396.000 214.270 400.000 ;
    END
  END proj0_io_in[8]
  PIN proj0_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 218.130 396.000 218.410 400.000 ;
    END
  END proj0_io_in[9]
  PIN proj0_io_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 181.330 396.000 181.610 400.000 ;
    END
  END proj0_io_out[0]
  PIN proj0_io_out[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.570 396.000 224.850 400.000 ;
    END
  END proj0_io_out[10]
  PIN proj0_io_out[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 229.170 396.000 229.450 400.000 ;
    END
  END proj0_io_out[11]
  PIN proj0_io_out[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 233.310 396.000 233.590 400.000 ;
    END
  END proj0_io_out[12]
  PIN proj0_io_out[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 237.910 396.000 238.190 400.000 ;
    END
  END proj0_io_out[13]
  PIN proj0_io_out[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 242.050 396.000 242.330 400.000 ;
    END
  END proj0_io_out[14]
  PIN proj0_io_out[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 246.650 396.000 246.930 400.000 ;
    END
  END proj0_io_out[15]
  PIN proj0_io_out[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 250.790 396.000 251.070 400.000 ;
    END
  END proj0_io_out[16]
  PIN proj0_io_out[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 254.930 396.000 255.210 400.000 ;
    END
  END proj0_io_out[17]
  PIN proj0_io_out[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 259.530 396.000 259.810 400.000 ;
    END
  END proj0_io_out[18]
  PIN proj0_io_out[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 263.670 396.000 263.950 400.000 ;
    END
  END proj0_io_out[19]
  PIN proj0_io_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 185.470 396.000 185.750 400.000 ;
    END
  END proj0_io_out[1]
  PIN proj0_io_out[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 268.270 396.000 268.550 400.000 ;
    END
  END proj0_io_out[20]
  PIN proj0_io_out[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 272.410 396.000 272.690 400.000 ;
    END
  END proj0_io_out[21]
  PIN proj0_io_out[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 277.010 396.000 277.290 400.000 ;
    END
  END proj0_io_out[22]
  PIN proj0_io_out[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 281.150 396.000 281.430 400.000 ;
    END
  END proj0_io_out[23]
  PIN proj0_io_out[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 285.750 396.000 286.030 400.000 ;
    END
  END proj0_io_out[24]
  PIN proj0_io_out[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 289.890 396.000 290.170 400.000 ;
    END
  END proj0_io_out[25]
  PIN proj0_io_out[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 294.490 396.000 294.770 400.000 ;
    END
  END proj0_io_out[26]
  PIN proj0_io_out[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 298.630 396.000 298.910 400.000 ;
    END
  END proj0_io_out[27]
  PIN proj0_io_out[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 302.770 396.000 303.050 400.000 ;
    END
  END proj0_io_out[28]
  PIN proj0_io_out[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 307.370 396.000 307.650 400.000 ;
    END
  END proj0_io_out[29]
  PIN proj0_io_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.070 396.000 190.350 400.000 ;
    END
  END proj0_io_out[2]
  PIN proj0_io_out[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 311.510 396.000 311.790 400.000 ;
    END
  END proj0_io_out[30]
  PIN proj0_io_out[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 316.110 396.000 316.390 400.000 ;
    END
  END proj0_io_out[31]
  PIN proj0_io_out[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 320.250 396.000 320.530 400.000 ;
    END
  END proj0_io_out[32]
  PIN proj0_io_out[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 324.850 396.000 325.130 400.000 ;
    END
  END proj0_io_out[33]
  PIN proj0_io_out[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 328.990 396.000 329.270 400.000 ;
    END
  END proj0_io_out[34]
  PIN proj0_io_out[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 333.590 396.000 333.870 400.000 ;
    END
  END proj0_io_out[35]
  PIN proj0_io_out[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 337.730 396.000 338.010 400.000 ;
    END
  END proj0_io_out[36]
  PIN proj0_io_out[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 341.870 396.000 342.150 400.000 ;
    END
  END proj0_io_out[37]
  PIN proj0_io_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 194.210 396.000 194.490 400.000 ;
    END
  END proj0_io_out[3]
  PIN proj0_io_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 198.810 396.000 199.090 400.000 ;
    END
  END proj0_io_out[4]
  PIN proj0_io_out[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 202.950 396.000 203.230 400.000 ;
    END
  END proj0_io_out[5]
  PIN proj0_io_out[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 207.090 396.000 207.370 400.000 ;
    END
  END proj0_io_out[6]
  PIN proj0_io_out[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 211.690 396.000 211.970 400.000 ;
    END
  END proj0_io_out[7]
  PIN proj0_io_out[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 215.830 396.000 216.110 400.000 ;
    END
  END proj0_io_out[8]
  PIN proj0_io_out[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 220.430 396.000 220.710 400.000 ;
    END
  END proj0_io_out[9]
  PIN proj0_reset
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 174.890 396.000 175.170 400.000 ;
    END
  END proj0_reset
  PIN proj0_wb_update
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 176.730 396.000 177.010 400.000 ;
    END
  END proj0_wb_update
  PIN proj1_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1.010 396.000 1.290 400.000 ;
    END
  END proj1_clk
  PIN proj1_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 7.450 396.000 7.730 400.000 ;
    END
  END proj1_io_in[0]
  PIN proj1_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 50.690 396.000 50.970 400.000 ;
    END
  END proj1_io_in[10]
  PIN proj1_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 55.290 396.000 55.570 400.000 ;
    END
  END proj1_io_in[11]
  PIN proj1_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 59.430 396.000 59.710 400.000 ;
    END
  END proj1_io_in[12]
  PIN proj1_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 64.030 396.000 64.310 400.000 ;
    END
  END proj1_io_in[13]
  PIN proj1_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 68.170 396.000 68.450 400.000 ;
    END
  END proj1_io_in[14]
  PIN proj1_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 72.310 396.000 72.590 400.000 ;
    END
  END proj1_io_in[15]
  PIN proj1_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.910 396.000 77.190 400.000 ;
    END
  END proj1_io_in[16]
  PIN proj1_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 81.050 396.000 81.330 400.000 ;
    END
  END proj1_io_in[17]
  PIN proj1_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 85.650 396.000 85.930 400.000 ;
    END
  END proj1_io_in[18]
  PIN proj1_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 89.790 396.000 90.070 400.000 ;
    END
  END proj1_io_in[19]
  PIN proj1_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 11.590 396.000 11.870 400.000 ;
    END
  END proj1_io_in[1]
  PIN proj1_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 94.390 396.000 94.670 400.000 ;
    END
  END proj1_io_in[20]
  PIN proj1_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.530 396.000 98.810 400.000 ;
    END
  END proj1_io_in[21]
  PIN proj1_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 103.130 396.000 103.410 400.000 ;
    END
  END proj1_io_in[22]
  PIN proj1_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 107.270 396.000 107.550 400.000 ;
    END
  END proj1_io_in[23]
  PIN proj1_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 111.870 396.000 112.150 400.000 ;
    END
  END proj1_io_in[24]
  PIN proj1_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.010 396.000 116.290 400.000 ;
    END
  END proj1_io_in[25]
  PIN proj1_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.150 396.000 120.430 400.000 ;
    END
  END proj1_io_in[26]
  PIN proj1_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 124.750 396.000 125.030 400.000 ;
    END
  END proj1_io_in[27]
  PIN proj1_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 128.890 396.000 129.170 400.000 ;
    END
  END proj1_io_in[28]
  PIN proj1_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 133.490 396.000 133.770 400.000 ;
    END
  END proj1_io_in[29]
  PIN proj1_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 16.190 396.000 16.470 400.000 ;
    END
  END proj1_io_in[2]
  PIN proj1_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 137.630 396.000 137.910 400.000 ;
    END
  END proj1_io_in[30]
  PIN proj1_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 142.230 396.000 142.510 400.000 ;
    END
  END proj1_io_in[31]
  PIN proj1_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 146.370 396.000 146.650 400.000 ;
    END
  END proj1_io_in[32]
  PIN proj1_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 150.970 396.000 151.250 400.000 ;
    END
  END proj1_io_in[33]
  PIN proj1_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 155.110 396.000 155.390 400.000 ;
    END
  END proj1_io_in[34]
  PIN proj1_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 159.710 396.000 159.990 400.000 ;
    END
  END proj1_io_in[35]
  PIN proj1_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 163.850 396.000 164.130 400.000 ;
    END
  END proj1_io_in[36]
  PIN proj1_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 167.990 396.000 168.270 400.000 ;
    END
  END proj1_io_in[37]
  PIN proj1_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 20.330 396.000 20.610 400.000 ;
    END
  END proj1_io_in[3]
  PIN proj1_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.470 396.000 24.750 400.000 ;
    END
  END proj1_io_in[4]
  PIN proj1_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 29.070 396.000 29.350 400.000 ;
    END
  END proj1_io_in[5]
  PIN proj1_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 33.210 396.000 33.490 400.000 ;
    END
  END proj1_io_in[6]
  PIN proj1_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.810 396.000 38.090 400.000 ;
    END
  END proj1_io_in[7]
  PIN proj1_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 41.950 396.000 42.230 400.000 ;
    END
  END proj1_io_in[8]
  PIN proj1_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.550 396.000 46.830 400.000 ;
    END
  END proj1_io_in[9]
  PIN proj1_io_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 9.290 396.000 9.570 400.000 ;
    END
  END proj1_io_out[0]
  PIN proj1_io_out[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 52.990 396.000 53.270 400.000 ;
    END
  END proj1_io_out[10]
  PIN proj1_io_out[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 57.130 396.000 57.410 400.000 ;
    END
  END proj1_io_out[11]
  PIN proj1_io_out[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 61.730 396.000 62.010 400.000 ;
    END
  END proj1_io_out[12]
  PIN proj1_io_out[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.870 396.000 66.150 400.000 ;
    END
  END proj1_io_out[13]
  PIN proj1_io_out[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 70.470 396.000 70.750 400.000 ;
    END
  END proj1_io_out[14]
  PIN proj1_io_out[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 74.610 396.000 74.890 400.000 ;
    END
  END proj1_io_out[15]
  PIN proj1_io_out[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 79.210 396.000 79.490 400.000 ;
    END
  END proj1_io_out[16]
  PIN proj1_io_out[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 83.350 396.000 83.630 400.000 ;
    END
  END proj1_io_out[17]
  PIN proj1_io_out[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.950 396.000 88.230 400.000 ;
    END
  END proj1_io_out[18]
  PIN proj1_io_out[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 92.090 396.000 92.370 400.000 ;
    END
  END proj1_io_out[19]
  PIN proj1_io_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 396.000 14.170 400.000 ;
    END
  END proj1_io_out[1]
  PIN proj1_io_out[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.230 396.000 96.510 400.000 ;
    END
  END proj1_io_out[20]
  PIN proj1_io_out[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 100.830 396.000 101.110 400.000 ;
    END
  END proj1_io_out[21]
  PIN proj1_io_out[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 104.970 396.000 105.250 400.000 ;
    END
  END proj1_io_out[22]
  PIN proj1_io_out[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 109.570 396.000 109.850 400.000 ;
    END
  END proj1_io_out[23]
  PIN proj1_io_out[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 113.710 396.000 113.990 400.000 ;
    END
  END proj1_io_out[24]
  PIN proj1_io_out[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 118.310 396.000 118.590 400.000 ;
    END
  END proj1_io_out[25]
  PIN proj1_io_out[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 122.450 396.000 122.730 400.000 ;
    END
  END proj1_io_out[26]
  PIN proj1_io_out[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 127.050 396.000 127.330 400.000 ;
    END
  END proj1_io_out[27]
  PIN proj1_io_out[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 131.190 396.000 131.470 400.000 ;
    END
  END proj1_io_out[28]
  PIN proj1_io_out[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.790 396.000 136.070 400.000 ;
    END
  END proj1_io_out[29]
  PIN proj1_io_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 18.030 396.000 18.310 400.000 ;
    END
  END proj1_io_out[2]
  PIN proj1_io_out[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 139.930 396.000 140.210 400.000 ;
    END
  END proj1_io_out[30]
  PIN proj1_io_out[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 144.070 396.000 144.350 400.000 ;
    END
  END proj1_io_out[31]
  PIN proj1_io_out[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 148.670 396.000 148.950 400.000 ;
    END
  END proj1_io_out[32]
  PIN proj1_io_out[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 152.810 396.000 153.090 400.000 ;
    END
  END proj1_io_out[33]
  PIN proj1_io_out[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 157.410 396.000 157.690 400.000 ;
    END
  END proj1_io_out[34]
  PIN proj1_io_out[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 161.550 396.000 161.830 400.000 ;
    END
  END proj1_io_out[35]
  PIN proj1_io_out[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 166.150 396.000 166.430 400.000 ;
    END
  END proj1_io_out[36]
  PIN proj1_io_out[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 170.290 396.000 170.570 400.000 ;
    END
  END proj1_io_out[37]
  PIN proj1_io_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.630 396.000 22.910 400.000 ;
    END
  END proj1_io_out[3]
  PIN proj1_io_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 26.770 396.000 27.050 400.000 ;
    END
  END proj1_io_out[4]
  PIN proj1_io_out[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.370 396.000 31.650 400.000 ;
    END
  END proj1_io_out[5]
  PIN proj1_io_out[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.510 396.000 35.790 400.000 ;
    END
  END proj1_io_out[6]
  PIN proj1_io_out[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 40.110 396.000 40.390 400.000 ;
    END
  END proj1_io_out[7]
  PIN proj1_io_out[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 396.000 44.530 400.000 ;
    END
  END proj1_io_out[8]
  PIN proj1_io_out[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 48.390 396.000 48.670 400.000 ;
    END
  END proj1_io_out[9]
  PIN proj1_reset
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 396.000 3.130 400.000 ;
    END
  END proj1_reset
  PIN proj1_wb_update
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 5.150 396.000 5.430 400.000 ;
    END
  END proj1_wb_update
  PIN proj2_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1331.330 396.000 1331.610 400.000 ;
    END
  END proj2_clk
  PIN proj2_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1335.470 396.000 1335.750 400.000 ;
    END
  END proj2_io_in[0]
  PIN proj2_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1379.170 396.000 1379.450 400.000 ;
    END
  END proj2_io_in[10]
  PIN proj2_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1383.310 396.000 1383.590 400.000 ;
    END
  END proj2_io_in[11]
  PIN proj2_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1387.910 396.000 1388.190 400.000 ;
    END
  END proj2_io_in[12]
  PIN proj2_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1392.050 396.000 1392.330 400.000 ;
    END
  END proj2_io_in[13]
  PIN proj2_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1396.650 396.000 1396.930 400.000 ;
    END
  END proj2_io_in[14]
  PIN proj2_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1400.790 396.000 1401.070 400.000 ;
    END
  END proj2_io_in[15]
  PIN proj2_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1405.390 396.000 1405.670 400.000 ;
    END
  END proj2_io_in[16]
  PIN proj2_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1409.530 396.000 1409.810 400.000 ;
    END
  END proj2_io_in[17]
  PIN proj2_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1413.670 396.000 1413.950 400.000 ;
    END
  END proj2_io_in[18]
  PIN proj2_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1418.270 396.000 1418.550 400.000 ;
    END
  END proj2_io_in[19]
  PIN proj2_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1340.070 396.000 1340.350 400.000 ;
    END
  END proj2_io_in[1]
  PIN proj2_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1422.410 396.000 1422.690 400.000 ;
    END
  END proj2_io_in[20]
  PIN proj2_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1427.010 396.000 1427.290 400.000 ;
    END
  END proj2_io_in[21]
  PIN proj2_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1431.150 396.000 1431.430 400.000 ;
    END
  END proj2_io_in[22]
  PIN proj2_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1435.750 396.000 1436.030 400.000 ;
    END
  END proj2_io_in[23]
  PIN proj2_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1439.890 396.000 1440.170 400.000 ;
    END
  END proj2_io_in[24]
  PIN proj2_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1444.490 396.000 1444.770 400.000 ;
    END
  END proj2_io_in[25]
  PIN proj2_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1448.630 396.000 1448.910 400.000 ;
    END
  END proj2_io_in[26]
  PIN proj2_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1453.230 396.000 1453.510 400.000 ;
    END
  END proj2_io_in[27]
  PIN proj2_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1457.370 396.000 1457.650 400.000 ;
    END
  END proj2_io_in[28]
  PIN proj2_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1461.510 396.000 1461.790 400.000 ;
    END
  END proj2_io_in[29]
  PIN proj2_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1344.210 396.000 1344.490 400.000 ;
    END
  END proj2_io_in[2]
  PIN proj2_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1466.110 396.000 1466.390 400.000 ;
    END
  END proj2_io_in[30]
  PIN proj2_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1470.250 396.000 1470.530 400.000 ;
    END
  END proj2_io_in[31]
  PIN proj2_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1474.850 396.000 1475.130 400.000 ;
    END
  END proj2_io_in[32]
  PIN proj2_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1478.990 396.000 1479.270 400.000 ;
    END
  END proj2_io_in[33]
  PIN proj2_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1483.590 396.000 1483.870 400.000 ;
    END
  END proj2_io_in[34]
  PIN proj2_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1487.730 396.000 1488.010 400.000 ;
    END
  END proj2_io_in[35]
  PIN proj2_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1492.330 396.000 1492.610 400.000 ;
    END
  END proj2_io_in[36]
  PIN proj2_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1496.470 396.000 1496.750 400.000 ;
    END
  END proj2_io_in[37]
  PIN proj2_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1348.810 396.000 1349.090 400.000 ;
    END
  END proj2_io_in[3]
  PIN proj2_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1352.950 396.000 1353.230 400.000 ;
    END
  END proj2_io_in[4]
  PIN proj2_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1357.550 396.000 1357.830 400.000 ;
    END
  END proj2_io_in[5]
  PIN proj2_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1361.690 396.000 1361.970 400.000 ;
    END
  END proj2_io_in[6]
  PIN proj2_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1365.830 396.000 1366.110 400.000 ;
    END
  END proj2_io_in[7]
  PIN proj2_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1370.430 396.000 1370.710 400.000 ;
    END
  END proj2_io_in[8]
  PIN proj2_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1374.570 396.000 1374.850 400.000 ;
    END
  END proj2_io_in[9]
  PIN proj2_io_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1337.770 396.000 1338.050 400.000 ;
    END
  END proj2_io_out[0]
  PIN proj2_io_out[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1381.470 396.000 1381.750 400.000 ;
    END
  END proj2_io_out[10]
  PIN proj2_io_out[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1385.610 396.000 1385.890 400.000 ;
    END
  END proj2_io_out[11]
  PIN proj2_io_out[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1389.750 396.000 1390.030 400.000 ;
    END
  END proj2_io_out[12]
  PIN proj2_io_out[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1394.350 396.000 1394.630 400.000 ;
    END
  END proj2_io_out[13]
  PIN proj2_io_out[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1398.490 396.000 1398.770 400.000 ;
    END
  END proj2_io_out[14]
  PIN proj2_io_out[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1403.090 396.000 1403.370 400.000 ;
    END
  END proj2_io_out[15]
  PIN proj2_io_out[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1407.230 396.000 1407.510 400.000 ;
    END
  END proj2_io_out[16]
  PIN proj2_io_out[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1411.830 396.000 1412.110 400.000 ;
    END
  END proj2_io_out[17]
  PIN proj2_io_out[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1415.970 396.000 1416.250 400.000 ;
    END
  END proj2_io_out[18]
  PIN proj2_io_out[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1420.570 396.000 1420.850 400.000 ;
    END
  END proj2_io_out[19]
  PIN proj2_io_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1341.910 396.000 1342.190 400.000 ;
    END
  END proj2_io_out[1]
  PIN proj2_io_out[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1424.710 396.000 1424.990 400.000 ;
    END
  END proj2_io_out[20]
  PIN proj2_io_out[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1429.310 396.000 1429.590 400.000 ;
    END
  END proj2_io_out[21]
  PIN proj2_io_out[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1433.450 396.000 1433.730 400.000 ;
    END
  END proj2_io_out[22]
  PIN proj2_io_out[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1437.590 396.000 1437.870 400.000 ;
    END
  END proj2_io_out[23]
  PIN proj2_io_out[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1442.190 396.000 1442.470 400.000 ;
    END
  END proj2_io_out[24]
  PIN proj2_io_out[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1446.330 396.000 1446.610 400.000 ;
    END
  END proj2_io_out[25]
  PIN proj2_io_out[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1450.930 396.000 1451.210 400.000 ;
    END
  END proj2_io_out[26]
  PIN proj2_io_out[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1455.070 396.000 1455.350 400.000 ;
    END
  END proj2_io_out[27]
  PIN proj2_io_out[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1459.670 396.000 1459.950 400.000 ;
    END
  END proj2_io_out[28]
  PIN proj2_io_out[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1463.810 396.000 1464.090 400.000 ;
    END
  END proj2_io_out[29]
  PIN proj2_io_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1346.510 396.000 1346.790 400.000 ;
    END
  END proj2_io_out[2]
  PIN proj2_io_out[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1468.410 396.000 1468.690 400.000 ;
    END
  END proj2_io_out[30]
  PIN proj2_io_out[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1472.550 396.000 1472.830 400.000 ;
    END
  END proj2_io_out[31]
  PIN proj2_io_out[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1477.150 396.000 1477.430 400.000 ;
    END
  END proj2_io_out[32]
  PIN proj2_io_out[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1481.290 396.000 1481.570 400.000 ;
    END
  END proj2_io_out[33]
  PIN proj2_io_out[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1485.430 396.000 1485.710 400.000 ;
    END
  END proj2_io_out[34]
  PIN proj2_io_out[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1490.030 396.000 1490.310 400.000 ;
    END
  END proj2_io_out[35]
  PIN proj2_io_out[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1494.170 396.000 1494.450 400.000 ;
    END
  END proj2_io_out[36]
  PIN proj2_io_out[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1498.770 396.000 1499.050 400.000 ;
    END
  END proj2_io_out[37]
  PIN proj2_io_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1350.650 396.000 1350.930 400.000 ;
    END
  END proj2_io_out[3]
  PIN proj2_io_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1355.250 396.000 1355.530 400.000 ;
    END
  END proj2_io_out[4]
  PIN proj2_io_out[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1359.390 396.000 1359.670 400.000 ;
    END
  END proj2_io_out[5]
  PIN proj2_io_out[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1363.990 396.000 1364.270 400.000 ;
    END
  END proj2_io_out[6]
  PIN proj2_io_out[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1368.130 396.000 1368.410 400.000 ;
    END
  END proj2_io_out[7]
  PIN proj2_io_out[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1372.730 396.000 1373.010 400.000 ;
    END
  END proj2_io_out[8]
  PIN proj2_io_out[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1376.870 396.000 1377.150 400.000 ;
    END
  END proj2_io_out[9]
  PIN proj2_reset
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1333.630 396.000 1333.910 400.000 ;
    END
  END proj2_reset
  PIN proj3_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 511.610 396.000 511.890 400.000 ;
    END
  END proj3_clk
  PIN proj3_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 516.210 396.000 516.490 400.000 ;
    END
  END proj3_io_in[0]
  PIN proj3_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 559.450 396.000 559.730 400.000 ;
    END
  END proj3_io_in[10]
  PIN proj3_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 564.050 396.000 564.330 400.000 ;
    END
  END proj3_io_in[11]
  PIN proj3_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 568.190 396.000 568.470 400.000 ;
    END
  END proj3_io_in[12]
  PIN proj3_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 572.330 396.000 572.610 400.000 ;
    END
  END proj3_io_in[13]
  PIN proj3_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 576.930 396.000 577.210 400.000 ;
    END
  END proj3_io_in[14]
  PIN proj3_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 581.070 396.000 581.350 400.000 ;
    END
  END proj3_io_in[15]
  PIN proj3_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 585.670 396.000 585.950 400.000 ;
    END
  END proj3_io_in[16]
  PIN proj3_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 589.810 396.000 590.090 400.000 ;
    END
  END proj3_io_in[17]
  PIN proj3_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 594.410 396.000 594.690 400.000 ;
    END
  END proj3_io_in[18]
  PIN proj3_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 598.550 396.000 598.830 400.000 ;
    END
  END proj3_io_in[19]
  PIN proj3_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 520.350 396.000 520.630 400.000 ;
    END
  END proj3_io_in[1]
  PIN proj3_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 603.150 396.000 603.430 400.000 ;
    END
  END proj3_io_in[20]
  PIN proj3_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 607.290 396.000 607.570 400.000 ;
    END
  END proj3_io_in[21]
  PIN proj3_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 611.890 396.000 612.170 400.000 ;
    END
  END proj3_io_in[22]
  PIN proj3_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 616.030 396.000 616.310 400.000 ;
    END
  END proj3_io_in[23]
  PIN proj3_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 620.170 396.000 620.450 400.000 ;
    END
  END proj3_io_in[24]
  PIN proj3_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 624.770 396.000 625.050 400.000 ;
    END
  END proj3_io_in[25]
  PIN proj3_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 628.910 396.000 629.190 400.000 ;
    END
  END proj3_io_in[26]
  PIN proj3_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 633.510 396.000 633.790 400.000 ;
    END
  END proj3_io_in[27]
  PIN proj3_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 637.650 396.000 637.930 400.000 ;
    END
  END proj3_io_in[28]
  PIN proj3_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 642.250 396.000 642.530 400.000 ;
    END
  END proj3_io_in[29]
  PIN proj3_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 524.490 396.000 524.770 400.000 ;
    END
  END proj3_io_in[2]
  PIN proj3_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 646.390 396.000 646.670 400.000 ;
    END
  END proj3_io_in[30]
  PIN proj3_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 650.990 396.000 651.270 400.000 ;
    END
  END proj3_io_in[31]
  PIN proj3_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 655.130 396.000 655.410 400.000 ;
    END
  END proj3_io_in[32]
  PIN proj3_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 659.730 396.000 660.010 400.000 ;
    END
  END proj3_io_in[33]
  PIN proj3_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 663.870 396.000 664.150 400.000 ;
    END
  END proj3_io_in[34]
  PIN proj3_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 668.010 396.000 668.290 400.000 ;
    END
  END proj3_io_in[35]
  PIN proj3_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 672.610 396.000 672.890 400.000 ;
    END
  END proj3_io_in[36]
  PIN proj3_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 676.750 396.000 677.030 400.000 ;
    END
  END proj3_io_in[37]
  PIN proj3_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 529.090 396.000 529.370 400.000 ;
    END
  END proj3_io_in[3]
  PIN proj3_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 533.230 396.000 533.510 400.000 ;
    END
  END proj3_io_in[4]
  PIN proj3_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 537.830 396.000 538.110 400.000 ;
    END
  END proj3_io_in[5]
  PIN proj3_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 541.970 396.000 542.250 400.000 ;
    END
  END proj3_io_in[6]
  PIN proj3_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 546.570 396.000 546.850 400.000 ;
    END
  END proj3_io_in[7]
  PIN proj3_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 550.710 396.000 550.990 400.000 ;
    END
  END proj3_io_in[8]
  PIN proj3_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 555.310 396.000 555.590 400.000 ;
    END
  END proj3_io_in[9]
  PIN proj3_io_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 518.050 396.000 518.330 400.000 ;
    END
  END proj3_io_out[0]
  PIN proj3_io_out[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 561.750 396.000 562.030 400.000 ;
    END
  END proj3_io_out[10]
  PIN proj3_io_out[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 565.890 396.000 566.170 400.000 ;
    END
  END proj3_io_out[11]
  PIN proj3_io_out[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 570.490 396.000 570.770 400.000 ;
    END
  END proj3_io_out[12]
  PIN proj3_io_out[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 574.630 396.000 574.910 400.000 ;
    END
  END proj3_io_out[13]
  PIN proj3_io_out[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 579.230 396.000 579.510 400.000 ;
    END
  END proj3_io_out[14]
  PIN proj3_io_out[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 583.370 396.000 583.650 400.000 ;
    END
  END proj3_io_out[15]
  PIN proj3_io_out[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 587.970 396.000 588.250 400.000 ;
    END
  END proj3_io_out[16]
  PIN proj3_io_out[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 592.110 396.000 592.390 400.000 ;
    END
  END proj3_io_out[17]
  PIN proj3_io_out[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 596.250 396.000 596.530 400.000 ;
    END
  END proj3_io_out[18]
  PIN proj3_io_out[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 600.850 396.000 601.130 400.000 ;
    END
  END proj3_io_out[19]
  PIN proj3_io_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 522.650 396.000 522.930 400.000 ;
    END
  END proj3_io_out[1]
  PIN proj3_io_out[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 604.990 396.000 605.270 400.000 ;
    END
  END proj3_io_out[20]
  PIN proj3_io_out[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 609.590 396.000 609.870 400.000 ;
    END
  END proj3_io_out[21]
  PIN proj3_io_out[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 613.730 396.000 614.010 400.000 ;
    END
  END proj3_io_out[22]
  PIN proj3_io_out[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 618.330 396.000 618.610 400.000 ;
    END
  END proj3_io_out[23]
  PIN proj3_io_out[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 622.470 396.000 622.750 400.000 ;
    END
  END proj3_io_out[24]
  PIN proj3_io_out[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 627.070 396.000 627.350 400.000 ;
    END
  END proj3_io_out[25]
  PIN proj3_io_out[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 631.210 396.000 631.490 400.000 ;
    END
  END proj3_io_out[26]
  PIN proj3_io_out[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 635.810 396.000 636.090 400.000 ;
    END
  END proj3_io_out[27]
  PIN proj3_io_out[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 639.950 396.000 640.230 400.000 ;
    END
  END proj3_io_out[28]
  PIN proj3_io_out[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 644.090 396.000 644.370 400.000 ;
    END
  END proj3_io_out[29]
  PIN proj3_io_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 526.790 396.000 527.070 400.000 ;
    END
  END proj3_io_out[2]
  PIN proj3_io_out[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 648.690 396.000 648.970 400.000 ;
    END
  END proj3_io_out[30]
  PIN proj3_io_out[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 652.830 396.000 653.110 400.000 ;
    END
  END proj3_io_out[31]
  PIN proj3_io_out[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 657.430 396.000 657.710 400.000 ;
    END
  END proj3_io_out[32]
  PIN proj3_io_out[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 661.570 396.000 661.850 400.000 ;
    END
  END proj3_io_out[33]
  PIN proj3_io_out[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 666.170 396.000 666.450 400.000 ;
    END
  END proj3_io_out[34]
  PIN proj3_io_out[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 670.310 396.000 670.590 400.000 ;
    END
  END proj3_io_out[35]
  PIN proj3_io_out[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 674.910 396.000 675.190 400.000 ;
    END
  END proj3_io_out[36]
  PIN proj3_io_out[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 679.050 396.000 679.330 400.000 ;
    END
  END proj3_io_out[37]
  PIN proj3_io_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 531.390 396.000 531.670 400.000 ;
    END
  END proj3_io_out[3]
  PIN proj3_io_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 535.530 396.000 535.810 400.000 ;
    END
  END proj3_io_out[4]
  PIN proj3_io_out[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 540.130 396.000 540.410 400.000 ;
    END
  END proj3_io_out[5]
  PIN proj3_io_out[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 544.270 396.000 544.550 400.000 ;
    END
  END proj3_io_out[6]
  PIN proj3_io_out[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 548.410 396.000 548.690 400.000 ;
    END
  END proj3_io_out[7]
  PIN proj3_io_out[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 553.010 396.000 553.290 400.000 ;
    END
  END proj3_io_out[8]
  PIN proj3_io_out[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 557.150 396.000 557.430 400.000 ;
    END
  END proj3_io_out[9]
  PIN proj3_reset
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 513.910 396.000 514.190 400.000 ;
    END
  END proj3_reset
  PIN proj4_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 681.350 396.000 681.630 400.000 ;
    END
  END proj4_clk
  PIN proj4_cnt[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 687.790 396.000 688.070 400.000 ;
    END
  END proj4_cnt[0]
  PIN proj4_cnt[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 774.730 396.000 775.010 400.000 ;
    END
  END proj4_cnt[10]
  PIN proj4_cnt[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 783.470 396.000 783.750 400.000 ;
    END
  END proj4_cnt[11]
  PIN proj4_cnt[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 792.210 396.000 792.490 400.000 ;
    END
  END proj4_cnt[12]
  PIN proj4_cnt[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 800.950 396.000 801.230 400.000 ;
    END
  END proj4_cnt[13]
  PIN proj4_cnt[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 809.690 396.000 809.970 400.000 ;
    END
  END proj4_cnt[14]
  PIN proj4_cnt[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 818.430 396.000 818.710 400.000 ;
    END
  END proj4_cnt[15]
  PIN proj4_cnt[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 826.710 396.000 826.990 400.000 ;
    END
  END proj4_cnt[16]
  PIN proj4_cnt[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 835.450 396.000 835.730 400.000 ;
    END
  END proj4_cnt[17]
  PIN proj4_cnt[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 844.190 396.000 844.470 400.000 ;
    END
  END proj4_cnt[18]
  PIN proj4_cnt[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 852.930 396.000 853.210 400.000 ;
    END
  END proj4_cnt[19]
  PIN proj4_cnt[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 696.530 396.000 696.810 400.000 ;
    END
  END proj4_cnt[1]
  PIN proj4_cnt[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 861.670 396.000 861.950 400.000 ;
    END
  END proj4_cnt[20]
  PIN proj4_cnt[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 870.410 396.000 870.690 400.000 ;
    END
  END proj4_cnt[21]
  PIN proj4_cnt[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 879.150 396.000 879.430 400.000 ;
    END
  END proj4_cnt[22]
  PIN proj4_cnt[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 887.890 396.000 888.170 400.000 ;
    END
  END proj4_cnt[23]
  PIN proj4_cnt[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 896.630 396.000 896.910 400.000 ;
    END
  END proj4_cnt[24]
  PIN proj4_cnt[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 905.370 396.000 905.650 400.000 ;
    END
  END proj4_cnt[25]
  PIN proj4_cnt[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 913.650 396.000 913.930 400.000 ;
    END
  END proj4_cnt[26]
  PIN proj4_cnt[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 922.390 396.000 922.670 400.000 ;
    END
  END proj4_cnt[27]
  PIN proj4_cnt[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 931.130 396.000 931.410 400.000 ;
    END
  END proj4_cnt[28]
  PIN proj4_cnt[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 939.870 396.000 940.150 400.000 ;
    END
  END proj4_cnt[29]
  PIN proj4_cnt[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 705.270 396.000 705.550 400.000 ;
    END
  END proj4_cnt[2]
  PIN proj4_cnt[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 948.610 396.000 948.890 400.000 ;
    END
  END proj4_cnt[30]
  PIN proj4_cnt[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 957.350 396.000 957.630 400.000 ;
    END
  END proj4_cnt[31]
  PIN proj4_cnt[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 714.010 396.000 714.290 400.000 ;
    END
  END proj4_cnt[3]
  PIN proj4_cnt[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 722.750 396.000 723.030 400.000 ;
    END
  END proj4_cnt[4]
  PIN proj4_cnt[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 731.030 396.000 731.310 400.000 ;
    END
  END proj4_cnt[5]
  PIN proj4_cnt[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 739.770 396.000 740.050 400.000 ;
    END
  END proj4_cnt[6]
  PIN proj4_cnt[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 748.510 396.000 748.790 400.000 ;
    END
  END proj4_cnt[7]
  PIN proj4_cnt[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 757.250 396.000 757.530 400.000 ;
    END
  END proj4_cnt[8]
  PIN proj4_cnt[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 765.990 396.000 766.270 400.000 ;
    END
  END proj4_cnt[9]
  PIN proj4_cnt_cont[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 690.090 396.000 690.370 400.000 ;
    END
  END proj4_cnt_cont[0]
  PIN proj4_cnt_cont[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 777.030 396.000 777.310 400.000 ;
    END
  END proj4_cnt_cont[10]
  PIN proj4_cnt_cont[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 785.770 396.000 786.050 400.000 ;
    END
  END proj4_cnt_cont[11]
  PIN proj4_cnt_cont[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 794.510 396.000 794.790 400.000 ;
    END
  END proj4_cnt_cont[12]
  PIN proj4_cnt_cont[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 802.790 396.000 803.070 400.000 ;
    END
  END proj4_cnt_cont[13]
  PIN proj4_cnt_cont[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 811.530 396.000 811.810 400.000 ;
    END
  END proj4_cnt_cont[14]
  PIN proj4_cnt_cont[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 820.270 396.000 820.550 400.000 ;
    END
  END proj4_cnt_cont[15]
  PIN proj4_cnt_cont[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 829.010 396.000 829.290 400.000 ;
    END
  END proj4_cnt_cont[16]
  PIN proj4_cnt_cont[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 837.750 396.000 838.030 400.000 ;
    END
  END proj4_cnt_cont[17]
  PIN proj4_cnt_cont[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 846.490 396.000 846.770 400.000 ;
    END
  END proj4_cnt_cont[18]
  PIN proj4_cnt_cont[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 855.230 396.000 855.510 400.000 ;
    END
  END proj4_cnt_cont[19]
  PIN proj4_cnt_cont[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 698.830 396.000 699.110 400.000 ;
    END
  END proj4_cnt_cont[1]
  PIN proj4_cnt_cont[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 863.970 396.000 864.250 400.000 ;
    END
  END proj4_cnt_cont[20]
  PIN proj4_cnt_cont[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 872.710 396.000 872.990 400.000 ;
    END
  END proj4_cnt_cont[21]
  PIN proj4_cnt_cont[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 881.450 396.000 881.730 400.000 ;
    END
  END proj4_cnt_cont[22]
  PIN proj4_cnt_cont[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 889.730 396.000 890.010 400.000 ;
    END
  END proj4_cnt_cont[23]
  PIN proj4_cnt_cont[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 898.470 396.000 898.750 400.000 ;
    END
  END proj4_cnt_cont[24]
  PIN proj4_cnt_cont[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 907.210 396.000 907.490 400.000 ;
    END
  END proj4_cnt_cont[25]
  PIN proj4_cnt_cont[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 915.950 396.000 916.230 400.000 ;
    END
  END proj4_cnt_cont[26]
  PIN proj4_cnt_cont[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 924.690 396.000 924.970 400.000 ;
    END
  END proj4_cnt_cont[27]
  PIN proj4_cnt_cont[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 933.430 396.000 933.710 400.000 ;
    END
  END proj4_cnt_cont[28]
  PIN proj4_cnt_cont[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 942.170 396.000 942.450 400.000 ;
    END
  END proj4_cnt_cont[29]
  PIN proj4_cnt_cont[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 707.110 396.000 707.390 400.000 ;
    END
  END proj4_cnt_cont[2]
  PIN proj4_cnt_cont[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 950.910 396.000 951.190 400.000 ;
    END
  END proj4_cnt_cont[30]
  PIN proj4_cnt_cont[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 959.650 396.000 959.930 400.000 ;
    END
  END proj4_cnt_cont[31]
  PIN proj4_cnt_cont[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 715.850 396.000 716.130 400.000 ;
    END
  END proj4_cnt_cont[3]
  PIN proj4_cnt_cont[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 724.590 396.000 724.870 400.000 ;
    END
  END proj4_cnt_cont[4]
  PIN proj4_cnt_cont[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 733.330 396.000 733.610 400.000 ;
    END
  END proj4_cnt_cont[5]
  PIN proj4_cnt_cont[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 742.070 396.000 742.350 400.000 ;
    END
  END proj4_cnt_cont[6]
  PIN proj4_cnt_cont[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 750.810 396.000 751.090 400.000 ;
    END
  END proj4_cnt_cont[7]
  PIN proj4_cnt_cont[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 759.550 396.000 759.830 400.000 ;
    END
  END proj4_cnt_cont[8]
  PIN proj4_cnt_cont[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 768.290 396.000 768.570 400.000 ;
    END
  END proj4_cnt_cont[9]
  PIN proj4_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 691.930 396.000 692.210 400.000 ;
    END
  END proj4_io_in[0]
  PIN proj4_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 778.870 396.000 779.150 400.000 ;
    END
  END proj4_io_in[10]
  PIN proj4_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 787.610 396.000 787.890 400.000 ;
    END
  END proj4_io_in[11]
  PIN proj4_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 796.350 396.000 796.630 400.000 ;
    END
  END proj4_io_in[12]
  PIN proj4_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 805.090 396.000 805.370 400.000 ;
    END
  END proj4_io_in[13]
  PIN proj4_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 813.830 396.000 814.110 400.000 ;
    END
  END proj4_io_in[14]
  PIN proj4_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 822.570 396.000 822.850 400.000 ;
    END
  END proj4_io_in[15]
  PIN proj4_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 831.310 396.000 831.590 400.000 ;
    END
  END proj4_io_in[16]
  PIN proj4_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 840.050 396.000 840.330 400.000 ;
    END
  END proj4_io_in[17]
  PIN proj4_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 848.790 396.000 849.070 400.000 ;
    END
  END proj4_io_in[18]
  PIN proj4_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 857.530 396.000 857.810 400.000 ;
    END
  END proj4_io_in[19]
  PIN proj4_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 700.670 396.000 700.950 400.000 ;
    END
  END proj4_io_in[1]
  PIN proj4_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 865.810 396.000 866.090 400.000 ;
    END
  END proj4_io_in[20]
  PIN proj4_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 874.550 396.000 874.830 400.000 ;
    END
  END proj4_io_in[21]
  PIN proj4_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 883.290 396.000 883.570 400.000 ;
    END
  END proj4_io_in[22]
  PIN proj4_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 892.030 396.000 892.310 400.000 ;
    END
  END proj4_io_in[23]
  PIN proj4_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 900.770 396.000 901.050 400.000 ;
    END
  END proj4_io_in[24]
  PIN proj4_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 909.510 396.000 909.790 400.000 ;
    END
  END proj4_io_in[25]
  PIN proj4_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 918.250 396.000 918.530 400.000 ;
    END
  END proj4_io_in[26]
  PIN proj4_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 926.990 396.000 927.270 400.000 ;
    END
  END proj4_io_in[27]
  PIN proj4_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 935.730 396.000 936.010 400.000 ;
    END
  END proj4_io_in[28]
  PIN proj4_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 944.470 396.000 944.750 400.000 ;
    END
  END proj4_io_in[29]
  PIN proj4_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 709.410 396.000 709.690 400.000 ;
    END
  END proj4_io_in[2]
  PIN proj4_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 953.210 396.000 953.490 400.000 ;
    END
  END proj4_io_in[30]
  PIN proj4_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 961.490 396.000 961.770 400.000 ;
    END
  END proj4_io_in[31]
  PIN proj4_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 966.090 396.000 966.370 400.000 ;
    END
  END proj4_io_in[32]
  PIN proj4_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 970.230 396.000 970.510 400.000 ;
    END
  END proj4_io_in[33]
  PIN proj4_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 974.830 396.000 975.110 400.000 ;
    END
  END proj4_io_in[34]
  PIN proj4_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 978.970 396.000 979.250 400.000 ;
    END
  END proj4_io_in[35]
  PIN proj4_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 983.570 396.000 983.850 400.000 ;
    END
  END proj4_io_in[36]
  PIN proj4_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 987.710 396.000 987.990 400.000 ;
    END
  END proj4_io_in[37]
  PIN proj4_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 718.150 396.000 718.430 400.000 ;
    END
  END proj4_io_in[3]
  PIN proj4_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 726.890 396.000 727.170 400.000 ;
    END
  END proj4_io_in[4]
  PIN proj4_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 735.630 396.000 735.910 400.000 ;
    END
  END proj4_io_in[5]
  PIN proj4_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 744.370 396.000 744.650 400.000 ;
    END
  END proj4_io_in[6]
  PIN proj4_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 753.110 396.000 753.390 400.000 ;
    END
  END proj4_io_in[7]
  PIN proj4_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 761.850 396.000 762.130 400.000 ;
    END
  END proj4_io_in[8]
  PIN proj4_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 770.590 396.000 770.870 400.000 ;
    END
  END proj4_io_in[9]
  PIN proj4_io_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 694.230 396.000 694.510 400.000 ;
    END
  END proj4_io_out[0]
  PIN proj4_io_out[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 781.170 396.000 781.450 400.000 ;
    END
  END proj4_io_out[10]
  PIN proj4_io_out[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 789.910 396.000 790.190 400.000 ;
    END
  END proj4_io_out[11]
  PIN proj4_io_out[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 798.650 396.000 798.930 400.000 ;
    END
  END proj4_io_out[12]
  PIN proj4_io_out[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 807.390 396.000 807.670 400.000 ;
    END
  END proj4_io_out[13]
  PIN proj4_io_out[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 816.130 396.000 816.410 400.000 ;
    END
  END proj4_io_out[14]
  PIN proj4_io_out[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 824.870 396.000 825.150 400.000 ;
    END
  END proj4_io_out[15]
  PIN proj4_io_out[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 833.610 396.000 833.890 400.000 ;
    END
  END proj4_io_out[16]
  PIN proj4_io_out[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 841.890 396.000 842.170 400.000 ;
    END
  END proj4_io_out[17]
  PIN proj4_io_out[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 850.630 396.000 850.910 400.000 ;
    END
  END proj4_io_out[18]
  PIN proj4_io_out[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 859.370 396.000 859.650 400.000 ;
    END
  END proj4_io_out[19]
  PIN proj4_io_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 702.970 396.000 703.250 400.000 ;
    END
  END proj4_io_out[1]
  PIN proj4_io_out[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 868.110 396.000 868.390 400.000 ;
    END
  END proj4_io_out[20]
  PIN proj4_io_out[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 876.850 396.000 877.130 400.000 ;
    END
  END proj4_io_out[21]
  PIN proj4_io_out[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 885.590 396.000 885.870 400.000 ;
    END
  END proj4_io_out[22]
  PIN proj4_io_out[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 894.330 396.000 894.610 400.000 ;
    END
  END proj4_io_out[23]
  PIN proj4_io_out[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 903.070 396.000 903.350 400.000 ;
    END
  END proj4_io_out[24]
  PIN proj4_io_out[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 911.810 396.000 912.090 400.000 ;
    END
  END proj4_io_out[25]
  PIN proj4_io_out[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 920.550 396.000 920.830 400.000 ;
    END
  END proj4_io_out[26]
  PIN proj4_io_out[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 929.290 396.000 929.570 400.000 ;
    END
  END proj4_io_out[27]
  PIN proj4_io_out[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 937.570 396.000 937.850 400.000 ;
    END
  END proj4_io_out[28]
  PIN proj4_io_out[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 946.310 396.000 946.590 400.000 ;
    END
  END proj4_io_out[29]
  PIN proj4_io_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 711.710 396.000 711.990 400.000 ;
    END
  END proj4_io_out[2]
  PIN proj4_io_out[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 955.050 396.000 955.330 400.000 ;
    END
  END proj4_io_out[30]
  PIN proj4_io_out[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 963.790 396.000 964.070 400.000 ;
    END
  END proj4_io_out[31]
  PIN proj4_io_out[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 968.390 396.000 968.670 400.000 ;
    END
  END proj4_io_out[32]
  PIN proj4_io_out[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 972.530 396.000 972.810 400.000 ;
    END
  END proj4_io_out[33]
  PIN proj4_io_out[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 977.130 396.000 977.410 400.000 ;
    END
  END proj4_io_out[34]
  PIN proj4_io_out[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 981.270 396.000 981.550 400.000 ;
    END
  END proj4_io_out[35]
  PIN proj4_io_out[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 985.410 396.000 985.690 400.000 ;
    END
  END proj4_io_out[36]
  PIN proj4_io_out[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 990.010 396.000 990.290 400.000 ;
    END
  END proj4_io_out[37]
  PIN proj4_io_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 720.450 396.000 720.730 400.000 ;
    END
  END proj4_io_out[3]
  PIN proj4_io_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 729.190 396.000 729.470 400.000 ;
    END
  END proj4_io_out[4]
  PIN proj4_io_out[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 737.930 396.000 738.210 400.000 ;
    END
  END proj4_io_out[5]
  PIN proj4_io_out[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 746.670 396.000 746.950 400.000 ;
    END
  END proj4_io_out[6]
  PIN proj4_io_out[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 754.950 396.000 755.230 400.000 ;
    END
  END proj4_io_out[7]
  PIN proj4_io_out[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 763.690 396.000 763.970 400.000 ;
    END
  END proj4_io_out[8]
  PIN proj4_io_out[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 772.430 396.000 772.710 400.000 ;
    END
  END proj4_io_out[9]
  PIN proj4_reset
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 683.190 396.000 683.470 400.000 ;
    END
  END proj4_reset
  PIN proj4_wb_update
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 685.490 396.000 685.770 400.000 ;
    END
  END proj4_wb_update
  PIN proj5_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 992.310 396.000 992.590 400.000 ;
    END
  END proj5_clk
  PIN proj5_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 998.750 396.000 999.030 400.000 ;
    END
  END proj5_io_in[0]
  PIN proj5_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1041.990 396.000 1042.270 400.000 ;
    END
  END proj5_io_in[10]
  PIN proj5_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1046.590 396.000 1046.870 400.000 ;
    END
  END proj5_io_in[11]
  PIN proj5_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1050.730 396.000 1051.010 400.000 ;
    END
  END proj5_io_in[12]
  PIN proj5_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1055.330 396.000 1055.610 400.000 ;
    END
  END proj5_io_in[13]
  PIN proj5_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1059.470 396.000 1059.750 400.000 ;
    END
  END proj5_io_in[14]
  PIN proj5_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1064.070 396.000 1064.350 400.000 ;
    END
  END proj5_io_in[15]
  PIN proj5_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1068.210 396.000 1068.490 400.000 ;
    END
  END proj5_io_in[16]
  PIN proj5_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1072.350 396.000 1072.630 400.000 ;
    END
  END proj5_io_in[17]
  PIN proj5_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1076.950 396.000 1077.230 400.000 ;
    END
  END proj5_io_in[18]
  PIN proj5_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1081.090 396.000 1081.370 400.000 ;
    END
  END proj5_io_in[19]
  PIN proj5_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1002.890 396.000 1003.170 400.000 ;
    END
  END proj5_io_in[1]
  PIN proj5_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1085.690 396.000 1085.970 400.000 ;
    END
  END proj5_io_in[20]
  PIN proj5_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1089.830 396.000 1090.110 400.000 ;
    END
  END proj5_io_in[21]
  PIN proj5_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1094.430 396.000 1094.710 400.000 ;
    END
  END proj5_io_in[22]
  PIN proj5_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1098.570 396.000 1098.850 400.000 ;
    END
  END proj5_io_in[23]
  PIN proj5_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1103.170 396.000 1103.450 400.000 ;
    END
  END proj5_io_in[24]
  PIN proj5_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1107.310 396.000 1107.590 400.000 ;
    END
  END proj5_io_in[25]
  PIN proj5_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1111.910 396.000 1112.190 400.000 ;
    END
  END proj5_io_in[26]
  PIN proj5_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1116.050 396.000 1116.330 400.000 ;
    END
  END proj5_io_in[27]
  PIN proj5_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1120.190 396.000 1120.470 400.000 ;
    END
  END proj5_io_in[28]
  PIN proj5_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1124.790 396.000 1125.070 400.000 ;
    END
  END proj5_io_in[29]
  PIN proj5_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1007.490 396.000 1007.770 400.000 ;
    END
  END proj5_io_in[2]
  PIN proj5_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1128.930 396.000 1129.210 400.000 ;
    END
  END proj5_io_in[30]
  PIN proj5_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1133.530 396.000 1133.810 400.000 ;
    END
  END proj5_io_in[31]
  PIN proj5_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1137.670 396.000 1137.950 400.000 ;
    END
  END proj5_io_in[32]
  PIN proj5_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1142.270 396.000 1142.550 400.000 ;
    END
  END proj5_io_in[33]
  PIN proj5_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1146.410 396.000 1146.690 400.000 ;
    END
  END proj5_io_in[34]
  PIN proj5_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1151.010 396.000 1151.290 400.000 ;
    END
  END proj5_io_in[35]
  PIN proj5_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1155.150 396.000 1155.430 400.000 ;
    END
  END proj5_io_in[36]
  PIN proj5_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1159.750 396.000 1160.030 400.000 ;
    END
  END proj5_io_in[37]
  PIN proj5_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1011.630 396.000 1011.910 400.000 ;
    END
  END proj5_io_in[3]
  PIN proj5_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1016.230 396.000 1016.510 400.000 ;
    END
  END proj5_io_in[4]
  PIN proj5_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1020.370 396.000 1020.650 400.000 ;
    END
  END proj5_io_in[5]
  PIN proj5_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1024.510 396.000 1024.790 400.000 ;
    END
  END proj5_io_in[6]
  PIN proj5_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1029.110 396.000 1029.390 400.000 ;
    END
  END proj5_io_in[7]
  PIN proj5_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1033.250 396.000 1033.530 400.000 ;
    END
  END proj5_io_in[8]
  PIN proj5_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1037.850 396.000 1038.130 400.000 ;
    END
  END proj5_io_in[9]
  PIN proj5_io_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1001.050 396.000 1001.330 400.000 ;
    END
  END proj5_io_out[0]
  PIN proj5_io_out[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1044.290 396.000 1044.570 400.000 ;
    END
  END proj5_io_out[10]
  PIN proj5_io_out[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1048.430 396.000 1048.710 400.000 ;
    END
  END proj5_io_out[11]
  PIN proj5_io_out[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1053.030 396.000 1053.310 400.000 ;
    END
  END proj5_io_out[12]
  PIN proj5_io_out[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1057.170 396.000 1057.450 400.000 ;
    END
  END proj5_io_out[13]
  PIN proj5_io_out[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1061.770 396.000 1062.050 400.000 ;
    END
  END proj5_io_out[14]
  PIN proj5_io_out[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1065.910 396.000 1066.190 400.000 ;
    END
  END proj5_io_out[15]
  PIN proj5_io_out[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1070.510 396.000 1070.790 400.000 ;
    END
  END proj5_io_out[16]
  PIN proj5_io_out[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1074.650 396.000 1074.930 400.000 ;
    END
  END proj5_io_out[17]
  PIN proj5_io_out[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1079.250 396.000 1079.530 400.000 ;
    END
  END proj5_io_out[18]
  PIN proj5_io_out[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1083.390 396.000 1083.670 400.000 ;
    END
  END proj5_io_out[19]
  PIN proj5_io_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1005.190 396.000 1005.470 400.000 ;
    END
  END proj5_io_out[1]
  PIN proj5_io_out[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1087.990 396.000 1088.270 400.000 ;
    END
  END proj5_io_out[20]
  PIN proj5_io_out[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1092.130 396.000 1092.410 400.000 ;
    END
  END proj5_io_out[21]
  PIN proj5_io_out[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1096.270 396.000 1096.550 400.000 ;
    END
  END proj5_io_out[22]
  PIN proj5_io_out[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1100.870 396.000 1101.150 400.000 ;
    END
  END proj5_io_out[23]
  PIN proj5_io_out[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1105.010 396.000 1105.290 400.000 ;
    END
  END proj5_io_out[24]
  PIN proj5_io_out[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1109.610 396.000 1109.890 400.000 ;
    END
  END proj5_io_out[25]
  PIN proj5_io_out[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1113.750 396.000 1114.030 400.000 ;
    END
  END proj5_io_out[26]
  PIN proj5_io_out[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1118.350 396.000 1118.630 400.000 ;
    END
  END proj5_io_out[27]
  PIN proj5_io_out[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1122.490 396.000 1122.770 400.000 ;
    END
  END proj5_io_out[28]
  PIN proj5_io_out[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1127.090 396.000 1127.370 400.000 ;
    END
  END proj5_io_out[29]
  PIN proj5_io_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1009.330 396.000 1009.610 400.000 ;
    END
  END proj5_io_out[2]
  PIN proj5_io_out[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1131.230 396.000 1131.510 400.000 ;
    END
  END proj5_io_out[30]
  PIN proj5_io_out[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1135.830 396.000 1136.110 400.000 ;
    END
  END proj5_io_out[31]
  PIN proj5_io_out[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1139.970 396.000 1140.250 400.000 ;
    END
  END proj5_io_out[32]
  PIN proj5_io_out[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1144.110 396.000 1144.390 400.000 ;
    END
  END proj5_io_out[33]
  PIN proj5_io_out[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1148.710 396.000 1148.990 400.000 ;
    END
  END proj5_io_out[34]
  PIN proj5_io_out[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1152.850 396.000 1153.130 400.000 ;
    END
  END proj5_io_out[35]
  PIN proj5_io_out[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1157.450 396.000 1157.730 400.000 ;
    END
  END proj5_io_out[36]
  PIN proj5_io_out[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1161.590 396.000 1161.870 400.000 ;
    END
  END proj5_io_out[37]
  PIN proj5_io_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1013.930 396.000 1014.210 400.000 ;
    END
  END proj5_io_out[3]
  PIN proj5_io_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1018.070 396.000 1018.350 400.000 ;
    END
  END proj5_io_out[4]
  PIN proj5_io_out[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1022.670 396.000 1022.950 400.000 ;
    END
  END proj5_io_out[5]
  PIN proj5_io_out[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1026.810 396.000 1027.090 400.000 ;
    END
  END proj5_io_out[6]
  PIN proj5_io_out[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1031.410 396.000 1031.690 400.000 ;
    END
  END proj5_io_out[7]
  PIN proj5_io_out[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1035.550 396.000 1035.830 400.000 ;
    END
  END proj5_io_out[8]
  PIN proj5_io_out[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1040.150 396.000 1040.430 400.000 ;
    END
  END proj5_io_out[9]
  PIN proj5_reset
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 994.150 396.000 994.430 400.000 ;
    END
  END proj5_reset
  PIN proj5_wb_update
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 996.450 396.000 996.730 400.000 ;
    END
  END proj5_wb_update
  PIN proj6_clk
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1163.890 396.000 1164.170 400.000 ;
    END
  END proj6_clk
  PIN proj6_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1166.190 396.000 1166.470 400.000 ;
    END
  END proj6_io_in[0]
  PIN proj6_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1209.430 396.000 1209.710 400.000 ;
    END
  END proj6_io_in[10]
  PIN proj6_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1214.030 396.000 1214.310 400.000 ;
    END
  END proj6_io_in[11]
  PIN proj6_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1218.170 396.000 1218.450 400.000 ;
    END
  END proj6_io_in[12]
  PIN proj6_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1222.770 396.000 1223.050 400.000 ;
    END
  END proj6_io_in[13]
  PIN proj6_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1226.910 396.000 1227.190 400.000 ;
    END
  END proj6_io_in[14]
  PIN proj6_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1231.050 396.000 1231.330 400.000 ;
    END
  END proj6_io_in[15]
  PIN proj6_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1235.650 396.000 1235.930 400.000 ;
    END
  END proj6_io_in[16]
  PIN proj6_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1239.790 396.000 1240.070 400.000 ;
    END
  END proj6_io_in[17]
  PIN proj6_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1244.390 396.000 1244.670 400.000 ;
    END
  END proj6_io_in[18]
  PIN proj6_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1248.530 396.000 1248.810 400.000 ;
    END
  END proj6_io_in[19]
  PIN proj6_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1170.330 396.000 1170.610 400.000 ;
    END
  END proj6_io_in[1]
  PIN proj6_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1253.130 396.000 1253.410 400.000 ;
    END
  END proj6_io_in[20]
  PIN proj6_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1257.270 396.000 1257.550 400.000 ;
    END
  END proj6_io_in[21]
  PIN proj6_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1261.870 396.000 1262.150 400.000 ;
    END
  END proj6_io_in[22]
  PIN proj6_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1266.010 396.000 1266.290 400.000 ;
    END
  END proj6_io_in[23]
  PIN proj6_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1270.610 396.000 1270.890 400.000 ;
    END
  END proj6_io_in[24]
  PIN proj6_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1274.750 396.000 1275.030 400.000 ;
    END
  END proj6_io_in[25]
  PIN proj6_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1278.890 396.000 1279.170 400.000 ;
    END
  END proj6_io_in[26]
  PIN proj6_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1283.490 396.000 1283.770 400.000 ;
    END
  END proj6_io_in[27]
  PIN proj6_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1287.630 396.000 1287.910 400.000 ;
    END
  END proj6_io_in[28]
  PIN proj6_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1292.230 396.000 1292.510 400.000 ;
    END
  END proj6_io_in[29]
  PIN proj6_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1174.930 396.000 1175.210 400.000 ;
    END
  END proj6_io_in[2]
  PIN proj6_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1296.370 396.000 1296.650 400.000 ;
    END
  END proj6_io_in[30]
  PIN proj6_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1300.970 396.000 1301.250 400.000 ;
    END
  END proj6_io_in[31]
  PIN proj6_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1305.110 396.000 1305.390 400.000 ;
    END
  END proj6_io_in[32]
  PIN proj6_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1309.710 396.000 1309.990 400.000 ;
    END
  END proj6_io_in[33]
  PIN proj6_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1313.850 396.000 1314.130 400.000 ;
    END
  END proj6_io_in[34]
  PIN proj6_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1318.450 396.000 1318.730 400.000 ;
    END
  END proj6_io_in[35]
  PIN proj6_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1322.590 396.000 1322.870 400.000 ;
    END
  END proj6_io_in[36]
  PIN proj6_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1326.730 396.000 1327.010 400.000 ;
    END
  END proj6_io_in[37]
  PIN proj6_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1179.070 396.000 1179.350 400.000 ;
    END
  END proj6_io_in[3]
  PIN proj6_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1183.210 396.000 1183.490 400.000 ;
    END
  END proj6_io_in[4]
  PIN proj6_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1187.810 396.000 1188.090 400.000 ;
    END
  END proj6_io_in[5]
  PIN proj6_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1191.950 396.000 1192.230 400.000 ;
    END
  END proj6_io_in[6]
  PIN proj6_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1196.550 396.000 1196.830 400.000 ;
    END
  END proj6_io_in[7]
  PIN proj6_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1200.690 396.000 1200.970 400.000 ;
    END
  END proj6_io_in[8]
  PIN proj6_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 1205.290 396.000 1205.570 400.000 ;
    END
  END proj6_io_in[9]
  PIN proj6_io_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1168.030 396.000 1168.310 400.000 ;
    END
  END proj6_io_out[0]
  PIN proj6_io_out[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1211.730 396.000 1212.010 400.000 ;
    END
  END proj6_io_out[10]
  PIN proj6_io_out[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1215.870 396.000 1216.150 400.000 ;
    END
  END proj6_io_out[11]
  PIN proj6_io_out[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1220.470 396.000 1220.750 400.000 ;
    END
  END proj6_io_out[12]
  PIN proj6_io_out[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1224.610 396.000 1224.890 400.000 ;
    END
  END proj6_io_out[13]
  PIN proj6_io_out[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1229.210 396.000 1229.490 400.000 ;
    END
  END proj6_io_out[14]
  PIN proj6_io_out[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1233.350 396.000 1233.630 400.000 ;
    END
  END proj6_io_out[15]
  PIN proj6_io_out[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1237.950 396.000 1238.230 400.000 ;
    END
  END proj6_io_out[16]
  PIN proj6_io_out[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1242.090 396.000 1242.370 400.000 ;
    END
  END proj6_io_out[17]
  PIN proj6_io_out[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1246.690 396.000 1246.970 400.000 ;
    END
  END proj6_io_out[18]
  PIN proj6_io_out[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1250.830 396.000 1251.110 400.000 ;
    END
  END proj6_io_out[19]
  PIN proj6_io_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1172.630 396.000 1172.910 400.000 ;
    END
  END proj6_io_out[1]
  PIN proj6_io_out[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1254.970 396.000 1255.250 400.000 ;
    END
  END proj6_io_out[20]
  PIN proj6_io_out[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1259.570 396.000 1259.850 400.000 ;
    END
  END proj6_io_out[21]
  PIN proj6_io_out[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1263.710 396.000 1263.990 400.000 ;
    END
  END proj6_io_out[22]
  PIN proj6_io_out[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1268.310 396.000 1268.590 400.000 ;
    END
  END proj6_io_out[23]
  PIN proj6_io_out[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1272.450 396.000 1272.730 400.000 ;
    END
  END proj6_io_out[24]
  PIN proj6_io_out[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1277.050 396.000 1277.330 400.000 ;
    END
  END proj6_io_out[25]
  PIN proj6_io_out[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1281.190 396.000 1281.470 400.000 ;
    END
  END proj6_io_out[26]
  PIN proj6_io_out[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1285.790 396.000 1286.070 400.000 ;
    END
  END proj6_io_out[27]
  PIN proj6_io_out[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1289.930 396.000 1290.210 400.000 ;
    END
  END proj6_io_out[28]
  PIN proj6_io_out[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1294.530 396.000 1294.810 400.000 ;
    END
  END proj6_io_out[29]
  PIN proj6_io_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1176.770 396.000 1177.050 400.000 ;
    END
  END proj6_io_out[2]
  PIN proj6_io_out[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1298.670 396.000 1298.950 400.000 ;
    END
  END proj6_io_out[30]
  PIN proj6_io_out[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1302.810 396.000 1303.090 400.000 ;
    END
  END proj6_io_out[31]
  PIN proj6_io_out[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1307.410 396.000 1307.690 400.000 ;
    END
  END proj6_io_out[32]
  PIN proj6_io_out[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1311.550 396.000 1311.830 400.000 ;
    END
  END proj6_io_out[33]
  PIN proj6_io_out[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1316.150 396.000 1316.430 400.000 ;
    END
  END proj6_io_out[34]
  PIN proj6_io_out[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1320.290 396.000 1320.570 400.000 ;
    END
  END proj6_io_out[35]
  PIN proj6_io_out[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1324.890 396.000 1325.170 400.000 ;
    END
  END proj6_io_out[36]
  PIN proj6_io_out[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1329.030 396.000 1329.310 400.000 ;
    END
  END proj6_io_out[37]
  PIN proj6_io_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1181.370 396.000 1181.650 400.000 ;
    END
  END proj6_io_out[3]
  PIN proj6_io_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1185.510 396.000 1185.790 400.000 ;
    END
  END proj6_io_out[4]
  PIN proj6_io_out[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1190.110 396.000 1190.390 400.000 ;
    END
  END proj6_io_out[5]
  PIN proj6_io_out[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1194.250 396.000 1194.530 400.000 ;
    END
  END proj6_io_out[6]
  PIN proj6_io_out[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1198.850 396.000 1199.130 400.000 ;
    END
  END proj6_io_out[7]
  PIN proj6_io_out[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1202.990 396.000 1203.270 400.000 ;
    END
  END proj6_io_out[8]
  PIN proj6_io_out[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1207.130 396.000 1207.410 400.000 ;
    END
  END proj6_io_out[9]
  PIN proj7_io_in[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 346.470 396.000 346.750 400.000 ;
    END
  END proj7_io_in[0]
  PIN proj7_io_in[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 389.710 396.000 389.990 400.000 ;
    END
  END proj7_io_in[10]
  PIN proj7_io_in[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 394.310 396.000 394.590 400.000 ;
    END
  END proj7_io_in[11]
  PIN proj7_io_in[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 398.450 396.000 398.730 400.000 ;
    END
  END proj7_io_in[12]
  PIN proj7_io_in[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 403.050 396.000 403.330 400.000 ;
    END
  END proj7_io_in[13]
  PIN proj7_io_in[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 407.190 396.000 407.470 400.000 ;
    END
  END proj7_io_in[14]
  PIN proj7_io_in[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 411.790 396.000 412.070 400.000 ;
    END
  END proj7_io_in[15]
  PIN proj7_io_in[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 415.930 396.000 416.210 400.000 ;
    END
  END proj7_io_in[16]
  PIN proj7_io_in[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 420.530 396.000 420.810 400.000 ;
    END
  END proj7_io_in[17]
  PIN proj7_io_in[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 424.670 396.000 424.950 400.000 ;
    END
  END proj7_io_in[18]
  PIN proj7_io_in[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 429.270 396.000 429.550 400.000 ;
    END
  END proj7_io_in[19]
  PIN proj7_io_in[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 350.610 396.000 350.890 400.000 ;
    END
  END proj7_io_in[1]
  PIN proj7_io_in[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 433.410 396.000 433.690 400.000 ;
    END
  END proj7_io_in[20]
  PIN proj7_io_in[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 437.550 396.000 437.830 400.000 ;
    END
  END proj7_io_in[21]
  PIN proj7_io_in[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 442.150 396.000 442.430 400.000 ;
    END
  END proj7_io_in[22]
  PIN proj7_io_in[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 446.290 396.000 446.570 400.000 ;
    END
  END proj7_io_in[23]
  PIN proj7_io_in[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 450.890 396.000 451.170 400.000 ;
    END
  END proj7_io_in[24]
  PIN proj7_io_in[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 455.030 396.000 455.310 400.000 ;
    END
  END proj7_io_in[25]
  PIN proj7_io_in[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 459.630 396.000 459.910 400.000 ;
    END
  END proj7_io_in[26]
  PIN proj7_io_in[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 463.770 396.000 464.050 400.000 ;
    END
  END proj7_io_in[27]
  PIN proj7_io_in[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 468.370 396.000 468.650 400.000 ;
    END
  END proj7_io_in[28]
  PIN proj7_io_in[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 472.510 396.000 472.790 400.000 ;
    END
  END proj7_io_in[29]
  PIN proj7_io_in[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 355.210 396.000 355.490 400.000 ;
    END
  END proj7_io_in[2]
  PIN proj7_io_in[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 477.110 396.000 477.390 400.000 ;
    END
  END proj7_io_in[30]
  PIN proj7_io_in[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 481.250 396.000 481.530 400.000 ;
    END
  END proj7_io_in[31]
  PIN proj7_io_in[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 485.390 396.000 485.670 400.000 ;
    END
  END proj7_io_in[32]
  PIN proj7_io_in[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 489.990 396.000 490.270 400.000 ;
    END
  END proj7_io_in[33]
  PIN proj7_io_in[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 494.130 396.000 494.410 400.000 ;
    END
  END proj7_io_in[34]
  PIN proj7_io_in[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 498.730 396.000 499.010 400.000 ;
    END
  END proj7_io_in[35]
  PIN proj7_io_in[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 502.870 396.000 503.150 400.000 ;
    END
  END proj7_io_in[36]
  PIN proj7_io_in[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 507.470 396.000 507.750 400.000 ;
    END
  END proj7_io_in[37]
  PIN proj7_io_in[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 359.350 396.000 359.630 400.000 ;
    END
  END proj7_io_in[3]
  PIN proj7_io_in[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 363.950 396.000 364.230 400.000 ;
    END
  END proj7_io_in[4]
  PIN proj7_io_in[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 368.090 396.000 368.370 400.000 ;
    END
  END proj7_io_in[5]
  PIN proj7_io_in[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 372.690 396.000 372.970 400.000 ;
    END
  END proj7_io_in[6]
  PIN proj7_io_in[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 376.830 396.000 377.110 400.000 ;
    END
  END proj7_io_in[7]
  PIN proj7_io_in[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 381.430 396.000 381.710 400.000 ;
    END
  END proj7_io_in[8]
  PIN proj7_io_in[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 385.570 396.000 385.850 400.000 ;
    END
  END proj7_io_in[9]
  PIN proj7_io_out[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 348.770 396.000 349.050 400.000 ;
    END
  END proj7_io_out[0]
  PIN proj7_io_out[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 392.010 396.000 392.290 400.000 ;
    END
  END proj7_io_out[10]
  PIN proj7_io_out[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 396.610 396.000 396.890 400.000 ;
    END
  END proj7_io_out[11]
  PIN proj7_io_out[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 400.750 396.000 401.030 400.000 ;
    END
  END proj7_io_out[12]
  PIN proj7_io_out[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 405.350 396.000 405.630 400.000 ;
    END
  END proj7_io_out[13]
  PIN proj7_io_out[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 409.490 396.000 409.770 400.000 ;
    END
  END proj7_io_out[14]
  PIN proj7_io_out[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 413.630 396.000 413.910 400.000 ;
    END
  END proj7_io_out[15]
  PIN proj7_io_out[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 418.230 396.000 418.510 400.000 ;
    END
  END proj7_io_out[16]
  PIN proj7_io_out[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 422.370 396.000 422.650 400.000 ;
    END
  END proj7_io_out[17]
  PIN proj7_io_out[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 426.970 396.000 427.250 400.000 ;
    END
  END proj7_io_out[18]
  PIN proj7_io_out[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 431.110 396.000 431.390 400.000 ;
    END
  END proj7_io_out[19]
  PIN proj7_io_out[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 352.910 396.000 353.190 400.000 ;
    END
  END proj7_io_out[1]
  PIN proj7_io_out[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 435.710 396.000 435.990 400.000 ;
    END
  END proj7_io_out[20]
  PIN proj7_io_out[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 439.850 396.000 440.130 400.000 ;
    END
  END proj7_io_out[21]
  PIN proj7_io_out[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 444.450 396.000 444.730 400.000 ;
    END
  END proj7_io_out[22]
  PIN proj7_io_out[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 448.590 396.000 448.870 400.000 ;
    END
  END proj7_io_out[23]
  PIN proj7_io_out[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 453.190 396.000 453.470 400.000 ;
    END
  END proj7_io_out[24]
  PIN proj7_io_out[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 457.330 396.000 457.610 400.000 ;
    END
  END proj7_io_out[25]
  PIN proj7_io_out[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 461.470 396.000 461.750 400.000 ;
    END
  END proj7_io_out[26]
  PIN proj7_io_out[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 466.070 396.000 466.350 400.000 ;
    END
  END proj7_io_out[27]
  PIN proj7_io_out[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 470.210 396.000 470.490 400.000 ;
    END
  END proj7_io_out[28]
  PIN proj7_io_out[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 474.810 396.000 475.090 400.000 ;
    END
  END proj7_io_out[29]
  PIN proj7_io_out[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 357.510 396.000 357.790 400.000 ;
    END
  END proj7_io_out[2]
  PIN proj7_io_out[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 478.950 396.000 479.230 400.000 ;
    END
  END proj7_io_out[30]
  PIN proj7_io_out[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 483.550 396.000 483.830 400.000 ;
    END
  END proj7_io_out[31]
  PIN proj7_io_out[32]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 487.690 396.000 487.970 400.000 ;
    END
  END proj7_io_out[32]
  PIN proj7_io_out[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 492.290 396.000 492.570 400.000 ;
    END
  END proj7_io_out[33]
  PIN proj7_io_out[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 496.430 396.000 496.710 400.000 ;
    END
  END proj7_io_out[34]
  PIN proj7_io_out[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 501.030 396.000 501.310 400.000 ;
    END
  END proj7_io_out[35]
  PIN proj7_io_out[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 505.170 396.000 505.450 400.000 ;
    END
  END proj7_io_out[36]
  PIN proj7_io_out[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 509.310 396.000 509.590 400.000 ;
    END
  END proj7_io_out[37]
  PIN proj7_io_out[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 361.650 396.000 361.930 400.000 ;
    END
  END proj7_io_out[3]
  PIN proj7_io_out[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 365.790 396.000 366.070 400.000 ;
    END
  END proj7_io_out[4]
  PIN proj7_io_out[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 370.390 396.000 370.670 400.000 ;
    END
  END proj7_io_out[5]
  PIN proj7_io_out[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 374.530 396.000 374.810 400.000 ;
    END
  END proj7_io_out[6]
  PIN proj7_io_out[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 379.130 396.000 379.410 400.000 ;
    END
  END proj7_io_out[7]
  PIN proj7_io_out[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 383.270 396.000 383.550 400.000 ;
    END
  END proj7_io_out[8]
  PIN proj7_io_out[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 387.870 396.000 388.150 400.000 ;
    END
  END proj7_io_out[9]
  PIN proj7_reset
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 344.170 396.000 344.450 400.000 ;
    END
  END proj7_reset
  PIN wb_clk_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 1.470 0.000 1.750 4.000 ;
    END
  END wb_clk_i
  PIN wb_rst_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 4.230 0.000 4.510 4.000 ;
    END
  END wb_rst_i
  PIN wbs_ack_o
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 7.450 0.000 7.730 4.000 ;
    END
  END wbs_ack_o
  PIN wbs_adr_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 19.410 0.000 19.690 4.000 ;
    END
  END wbs_adr_i[0]
  PIN wbs_adr_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 123.830 0.000 124.110 4.000 ;
    END
  END wbs_adr_i[10]
  PIN wbs_adr_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 133.030 0.000 133.310 4.000 ;
    END
  END wbs_adr_i[11]
  PIN wbs_adr_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 142.230 0.000 142.510 4.000 ;
    END
  END wbs_adr_i[12]
  PIN wbs_adr_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END wbs_adr_i[13]
  PIN wbs_adr_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 160.630 0.000 160.910 4.000 ;
    END
  END wbs_adr_i[14]
  PIN wbs_adr_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 169.830 0.000 170.110 4.000 ;
    END
  END wbs_adr_i[15]
  PIN wbs_adr_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 178.570 0.000 178.850 4.000 ;
    END
  END wbs_adr_i[16]
  PIN wbs_adr_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END wbs_adr_i[17]
  PIN wbs_adr_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 196.970 0.000 197.250 4.000 ;
    END
  END wbs_adr_i[18]
  PIN wbs_adr_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END wbs_adr_i[19]
  PIN wbs_adr_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.830 0.000 32.110 4.000 ;
    END
  END wbs_adr_i[1]
  PIN wbs_adr_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END wbs_adr_i[20]
  PIN wbs_adr_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 224.570 0.000 224.850 4.000 ;
    END
  END wbs_adr_i[21]
  PIN wbs_adr_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 233.770 0.000 234.050 4.000 ;
    END
  END wbs_adr_i[22]
  PIN wbs_adr_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 242.970 0.000 243.250 4.000 ;
    END
  END wbs_adr_i[23]
  PIN wbs_adr_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 252.170 0.000 252.450 4.000 ;
    END
  END wbs_adr_i[24]
  PIN wbs_adr_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 261.370 0.000 261.650 4.000 ;
    END
  END wbs_adr_i[25]
  PIN wbs_adr_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END wbs_adr_i[26]
  PIN wbs_adr_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 279.770 0.000 280.050 4.000 ;
    END
  END wbs_adr_i[27]
  PIN wbs_adr_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 288.970 0.000 289.250 4.000 ;
    END
  END wbs_adr_i[28]
  PIN wbs_adr_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 298.170 0.000 298.450 4.000 ;
    END
  END wbs_adr_i[29]
  PIN wbs_adr_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 44.250 0.000 44.530 4.000 ;
    END
  END wbs_adr_i[2]
  PIN wbs_adr_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 307.370 0.000 307.650 4.000 ;
    END
  END wbs_adr_i[30]
  PIN wbs_adr_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 316.570 0.000 316.850 4.000 ;
    END
  END wbs_adr_i[31]
  PIN wbs_adr_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.210 0.000 56.490 4.000 ;
    END
  END wbs_adr_i[3]
  PIN wbs_adr_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 68.630 0.000 68.910 4.000 ;
    END
  END wbs_adr_i[4]
  PIN wbs_adr_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.830 0.000 78.110 4.000 ;
    END
  END wbs_adr_i[5]
  PIN wbs_adr_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 87.030 0.000 87.310 4.000 ;
    END
  END wbs_adr_i[6]
  PIN wbs_adr_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 96.230 0.000 96.510 4.000 ;
    END
  END wbs_adr_i[7]
  PIN wbs_adr_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 105.430 0.000 105.710 4.000 ;
    END
  END wbs_adr_i[8]
  PIN wbs_adr_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 114.630 0.000 114.910 4.000 ;
    END
  END wbs_adr_i[9]
  PIN wbs_cyc_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 10.210 0.000 10.490 4.000 ;
    END
  END wbs_cyc_i
  PIN wbs_dat_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END wbs_dat_i[0]
  PIN wbs_dat_i[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 126.590 0.000 126.870 4.000 ;
    END
  END wbs_dat_i[10]
  PIN wbs_dat_i[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 135.790 0.000 136.070 4.000 ;
    END
  END wbs_dat_i[11]
  PIN wbs_dat_i[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END wbs_dat_i[12]
  PIN wbs_dat_i[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 154.190 0.000 154.470 4.000 ;
    END
  END wbs_dat_i[13]
  PIN wbs_dat_i[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 163.390 0.000 163.670 4.000 ;
    END
  END wbs_dat_i[14]
  PIN wbs_dat_i[15]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 172.590 0.000 172.870 4.000 ;
    END
  END wbs_dat_i[15]
  PIN wbs_dat_i[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 181.790 0.000 182.070 4.000 ;
    END
  END wbs_dat_i[16]
  PIN wbs_dat_i[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 190.990 0.000 191.270 4.000 ;
    END
  END wbs_dat_i[17]
  PIN wbs_dat_i[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 200.190 0.000 200.470 4.000 ;
    END
  END wbs_dat_i[18]
  PIN wbs_dat_i[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 209.390 0.000 209.670 4.000 ;
    END
  END wbs_dat_i[19]
  PIN wbs_dat_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.050 0.000 35.330 4.000 ;
    END
  END wbs_dat_i[1]
  PIN wbs_dat_i[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 218.590 0.000 218.870 4.000 ;
    END
  END wbs_dat_i[20]
  PIN wbs_dat_i[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 227.790 0.000 228.070 4.000 ;
    END
  END wbs_dat_i[21]
  PIN wbs_dat_i[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.990 0.000 237.270 4.000 ;
    END
  END wbs_dat_i[22]
  PIN wbs_dat_i[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 246.190 0.000 246.470 4.000 ;
    END
  END wbs_dat_i[23]
  PIN wbs_dat_i[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 255.390 0.000 255.670 4.000 ;
    END
  END wbs_dat_i[24]
  PIN wbs_dat_i[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 264.590 0.000 264.870 4.000 ;
    END
  END wbs_dat_i[25]
  PIN wbs_dat_i[26]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END wbs_dat_i[26]
  PIN wbs_dat_i[27]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 282.990 0.000 283.270 4.000 ;
    END
  END wbs_dat_i[27]
  PIN wbs_dat_i[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 292.190 0.000 292.470 4.000 ;
    END
  END wbs_dat_i[28]
  PIN wbs_dat_i[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 301.390 0.000 301.670 4.000 ;
    END
  END wbs_dat_i[29]
  PIN wbs_dat_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 47.010 0.000 47.290 4.000 ;
    END
  END wbs_dat_i[2]
  PIN wbs_dat_i[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 310.590 0.000 310.870 4.000 ;
    END
  END wbs_dat_i[30]
  PIN wbs_dat_i[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 319.790 0.000 320.070 4.000 ;
    END
  END wbs_dat_i[31]
  PIN wbs_dat_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.430 0.000 59.710 4.000 ;
    END
  END wbs_dat_i[3]
  PIN wbs_dat_i[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 71.850 0.000 72.130 4.000 ;
    END
  END wbs_dat_i[4]
  PIN wbs_dat_i[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 81.050 0.000 81.330 4.000 ;
    END
  END wbs_dat_i[5]
  PIN wbs_dat_i[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 89.790 0.000 90.070 4.000 ;
    END
  END wbs_dat_i[6]
  PIN wbs_dat_i[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.990 0.000 99.270 4.000 ;
    END
  END wbs_dat_i[7]
  PIN wbs_dat_i[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 108.190 0.000 108.470 4.000 ;
    END
  END wbs_dat_i[8]
  PIN wbs_dat_i[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 117.390 0.000 117.670 4.000 ;
    END
  END wbs_dat_i[9]
  PIN wbs_dat_o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END wbs_dat_o[0]
  PIN wbs_dat_o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END wbs_dat_o[10]
  PIN wbs_dat_o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 139.010 0.000 139.290 4.000 ;
    END
  END wbs_dat_o[11]
  PIN wbs_dat_o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 148.210 0.000 148.490 4.000 ;
    END
  END wbs_dat_o[12]
  PIN wbs_dat_o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 157.410 0.000 157.690 4.000 ;
    END
  END wbs_dat_o[13]
  PIN wbs_dat_o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 166.610 0.000 166.890 4.000 ;
    END
  END wbs_dat_o[14]
  PIN wbs_dat_o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 175.810 0.000 176.090 4.000 ;
    END
  END wbs_dat_o[15]
  PIN wbs_dat_o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 185.010 0.000 185.290 4.000 ;
    END
  END wbs_dat_o[16]
  PIN wbs_dat_o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END wbs_dat_o[17]
  PIN wbs_dat_o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 203.410 0.000 203.690 4.000 ;
    END
  END wbs_dat_o[18]
  PIN wbs_dat_o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END wbs_dat_o[19]
  PIN wbs_dat_o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 37.810 0.000 38.090 4.000 ;
    END
  END wbs_dat_o[1]
  PIN wbs_dat_o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 221.810 0.000 222.090 4.000 ;
    END
  END wbs_dat_o[20]
  PIN wbs_dat_o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 231.010 0.000 231.290 4.000 ;
    END
  END wbs_dat_o[21]
  PIN wbs_dat_o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 240.210 0.000 240.490 4.000 ;
    END
  END wbs_dat_o[22]
  PIN wbs_dat_o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 249.410 0.000 249.690 4.000 ;
    END
  END wbs_dat_o[23]
  PIN wbs_dat_o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END wbs_dat_o[24]
  PIN wbs_dat_o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 267.350 0.000 267.630 4.000 ;
    END
  END wbs_dat_o[25]
  PIN wbs_dat_o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 276.550 0.000 276.830 4.000 ;
    END
  END wbs_dat_o[26]
  PIN wbs_dat_o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 285.750 0.000 286.030 4.000 ;
    END
  END wbs_dat_o[27]
  PIN wbs_dat_o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 294.950 0.000 295.230 4.000 ;
    END
  END wbs_dat_o[28]
  PIN wbs_dat_o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 304.150 0.000 304.430 4.000 ;
    END
  END wbs_dat_o[29]
  PIN wbs_dat_o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 50.230 0.000 50.510 4.000 ;
    END
  END wbs_dat_o[2]
  PIN wbs_dat_o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 313.350 0.000 313.630 4.000 ;
    END
  END wbs_dat_o[30]
  PIN wbs_dat_o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 322.550 0.000 322.830 4.000 ;
    END
  END wbs_dat_o[31]
  PIN wbs_dat_o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 62.650 0.000 62.930 4.000 ;
    END
  END wbs_dat_o[3]
  PIN wbs_dat_o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 74.610 0.000 74.890 4.000 ;
    END
  END wbs_dat_o[4]
  PIN wbs_dat_o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END wbs_dat_o[5]
  PIN wbs_dat_o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 93.010 0.000 93.290 4.000 ;
    END
  END wbs_dat_o[6]
  PIN wbs_dat_o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END wbs_dat_o[7]
  PIN wbs_dat_o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 111.410 0.000 111.690 4.000 ;
    END
  END wbs_dat_o[8]
  PIN wbs_dat_o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 120.610 0.000 120.890 4.000 ;
    END
  END wbs_dat_o[9]
  PIN wbs_sel_i[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 28.610 0.000 28.890 4.000 ;
    END
  END wbs_sel_i[0]
  PIN wbs_sel_i[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 41.030 0.000 41.310 4.000 ;
    END
  END wbs_sel_i[1]
  PIN wbs_sel_i[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 53.450 0.000 53.730 4.000 ;
    END
  END wbs_sel_i[2]
  PIN wbs_sel_i[3]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 65.410 0.000 65.690 4.000 ;
    END
  END wbs_sel_i[3]
  PIN wbs_stb_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.430 0.000 13.710 4.000 ;
    END
  END wbs_stb_i
  PIN wbs_we_i
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END wbs_we_i
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 389.200 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 389.200 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 1494.080 398.055 ;
      LAYER met1 ;
        RECT 0.990 4.460 1499.070 398.780 ;
      LAYER met2 ;
        RECT 1.570 395.720 2.570 398.810 ;
        RECT 3.410 395.720 4.870 398.810 ;
        RECT 5.710 395.720 7.170 398.810 ;
        RECT 8.010 395.720 9.010 398.810 ;
        RECT 9.850 395.720 11.310 398.810 ;
        RECT 12.150 395.720 13.610 398.810 ;
        RECT 14.450 395.720 15.910 398.810 ;
        RECT 16.750 395.720 17.750 398.810 ;
        RECT 18.590 395.720 20.050 398.810 ;
        RECT 20.890 395.720 22.350 398.810 ;
        RECT 23.190 395.720 24.190 398.810 ;
        RECT 25.030 395.720 26.490 398.810 ;
        RECT 27.330 395.720 28.790 398.810 ;
        RECT 29.630 395.720 31.090 398.810 ;
        RECT 31.930 395.720 32.930 398.810 ;
        RECT 33.770 395.720 35.230 398.810 ;
        RECT 36.070 395.720 37.530 398.810 ;
        RECT 38.370 395.720 39.830 398.810 ;
        RECT 40.670 395.720 41.670 398.810 ;
        RECT 42.510 395.720 43.970 398.810 ;
        RECT 44.810 395.720 46.270 398.810 ;
        RECT 47.110 395.720 48.110 398.810 ;
        RECT 48.950 395.720 50.410 398.810 ;
        RECT 51.250 395.720 52.710 398.810 ;
        RECT 53.550 395.720 55.010 398.810 ;
        RECT 55.850 395.720 56.850 398.810 ;
        RECT 57.690 395.720 59.150 398.810 ;
        RECT 59.990 395.720 61.450 398.810 ;
        RECT 62.290 395.720 63.750 398.810 ;
        RECT 64.590 395.720 65.590 398.810 ;
        RECT 66.430 395.720 67.890 398.810 ;
        RECT 68.730 395.720 70.190 398.810 ;
        RECT 71.030 395.720 72.030 398.810 ;
        RECT 72.870 395.720 74.330 398.810 ;
        RECT 75.170 395.720 76.630 398.810 ;
        RECT 77.470 395.720 78.930 398.810 ;
        RECT 79.770 395.720 80.770 398.810 ;
        RECT 81.610 395.720 83.070 398.810 ;
        RECT 83.910 395.720 85.370 398.810 ;
        RECT 86.210 395.720 87.670 398.810 ;
        RECT 88.510 395.720 89.510 398.810 ;
        RECT 90.350 395.720 91.810 398.810 ;
        RECT 92.650 395.720 94.110 398.810 ;
        RECT 94.950 395.720 95.950 398.810 ;
        RECT 96.790 395.720 98.250 398.810 ;
        RECT 99.090 395.720 100.550 398.810 ;
        RECT 101.390 395.720 102.850 398.810 ;
        RECT 103.690 395.720 104.690 398.810 ;
        RECT 105.530 395.720 106.990 398.810 ;
        RECT 107.830 395.720 109.290 398.810 ;
        RECT 110.130 395.720 111.590 398.810 ;
        RECT 112.430 395.720 113.430 398.810 ;
        RECT 114.270 395.720 115.730 398.810 ;
        RECT 116.570 395.720 118.030 398.810 ;
        RECT 118.870 395.720 119.870 398.810 ;
        RECT 120.710 395.720 122.170 398.810 ;
        RECT 123.010 395.720 124.470 398.810 ;
        RECT 125.310 395.720 126.770 398.810 ;
        RECT 127.610 395.720 128.610 398.810 ;
        RECT 129.450 395.720 130.910 398.810 ;
        RECT 131.750 395.720 133.210 398.810 ;
        RECT 134.050 395.720 135.510 398.810 ;
        RECT 136.350 395.720 137.350 398.810 ;
        RECT 138.190 395.720 139.650 398.810 ;
        RECT 140.490 395.720 141.950 398.810 ;
        RECT 142.790 395.720 143.790 398.810 ;
        RECT 144.630 395.720 146.090 398.810 ;
        RECT 146.930 395.720 148.390 398.810 ;
        RECT 149.230 395.720 150.690 398.810 ;
        RECT 151.530 395.720 152.530 398.810 ;
        RECT 153.370 395.720 154.830 398.810 ;
        RECT 155.670 395.720 157.130 398.810 ;
        RECT 157.970 395.720 159.430 398.810 ;
        RECT 160.270 395.720 161.270 398.810 ;
        RECT 162.110 395.720 163.570 398.810 ;
        RECT 164.410 395.720 165.870 398.810 ;
        RECT 166.710 395.720 167.710 398.810 ;
        RECT 168.550 395.720 170.010 398.810 ;
        RECT 170.850 395.720 172.310 398.810 ;
        RECT 173.150 395.720 174.610 398.810 ;
        RECT 175.450 395.720 176.450 398.810 ;
        RECT 177.290 395.720 178.750 398.810 ;
        RECT 179.590 395.720 181.050 398.810 ;
        RECT 181.890 395.720 182.890 398.810 ;
        RECT 183.730 395.720 185.190 398.810 ;
        RECT 186.030 395.720 187.490 398.810 ;
        RECT 188.330 395.720 189.790 398.810 ;
        RECT 190.630 395.720 191.630 398.810 ;
        RECT 192.470 395.720 193.930 398.810 ;
        RECT 194.770 395.720 196.230 398.810 ;
        RECT 197.070 395.720 198.530 398.810 ;
        RECT 199.370 395.720 200.370 398.810 ;
        RECT 201.210 395.720 202.670 398.810 ;
        RECT 203.510 395.720 204.970 398.810 ;
        RECT 205.810 395.720 206.810 398.810 ;
        RECT 207.650 395.720 209.110 398.810 ;
        RECT 209.950 395.720 211.410 398.810 ;
        RECT 212.250 395.720 213.710 398.810 ;
        RECT 214.550 395.720 215.550 398.810 ;
        RECT 216.390 395.720 217.850 398.810 ;
        RECT 218.690 395.720 220.150 398.810 ;
        RECT 220.990 395.720 222.450 398.810 ;
        RECT 223.290 395.720 224.290 398.810 ;
        RECT 225.130 395.720 226.590 398.810 ;
        RECT 227.430 395.720 228.890 398.810 ;
        RECT 229.730 395.720 230.730 398.810 ;
        RECT 231.570 395.720 233.030 398.810 ;
        RECT 233.870 395.720 235.330 398.810 ;
        RECT 236.170 395.720 237.630 398.810 ;
        RECT 238.470 395.720 239.470 398.810 ;
        RECT 240.310 395.720 241.770 398.810 ;
        RECT 242.610 395.720 244.070 398.810 ;
        RECT 244.910 395.720 246.370 398.810 ;
        RECT 247.210 395.720 248.210 398.810 ;
        RECT 249.050 395.720 250.510 398.810 ;
        RECT 251.350 395.720 252.810 398.810 ;
        RECT 253.650 395.720 254.650 398.810 ;
        RECT 255.490 395.720 256.950 398.810 ;
        RECT 257.790 395.720 259.250 398.810 ;
        RECT 260.090 395.720 261.550 398.810 ;
        RECT 262.390 395.720 263.390 398.810 ;
        RECT 264.230 395.720 265.690 398.810 ;
        RECT 266.530 395.720 267.990 398.810 ;
        RECT 268.830 395.720 270.290 398.810 ;
        RECT 271.130 395.720 272.130 398.810 ;
        RECT 272.970 395.720 274.430 398.810 ;
        RECT 275.270 395.720 276.730 398.810 ;
        RECT 277.570 395.720 278.570 398.810 ;
        RECT 279.410 395.720 280.870 398.810 ;
        RECT 281.710 395.720 283.170 398.810 ;
        RECT 284.010 395.720 285.470 398.810 ;
        RECT 286.310 395.720 287.310 398.810 ;
        RECT 288.150 395.720 289.610 398.810 ;
        RECT 290.450 395.720 291.910 398.810 ;
        RECT 292.750 395.720 294.210 398.810 ;
        RECT 295.050 395.720 296.050 398.810 ;
        RECT 296.890 395.720 298.350 398.810 ;
        RECT 299.190 395.720 300.650 398.810 ;
        RECT 301.490 395.720 302.490 398.810 ;
        RECT 303.330 395.720 304.790 398.810 ;
        RECT 305.630 395.720 307.090 398.810 ;
        RECT 307.930 395.720 309.390 398.810 ;
        RECT 310.230 395.720 311.230 398.810 ;
        RECT 312.070 395.720 313.530 398.810 ;
        RECT 314.370 395.720 315.830 398.810 ;
        RECT 316.670 395.720 318.130 398.810 ;
        RECT 318.970 395.720 319.970 398.810 ;
        RECT 320.810 395.720 322.270 398.810 ;
        RECT 323.110 395.720 324.570 398.810 ;
        RECT 325.410 395.720 326.410 398.810 ;
        RECT 327.250 395.720 328.710 398.810 ;
        RECT 329.550 395.720 331.010 398.810 ;
        RECT 331.850 395.720 333.310 398.810 ;
        RECT 334.150 395.720 335.150 398.810 ;
        RECT 335.990 395.720 337.450 398.810 ;
        RECT 338.290 395.720 339.750 398.810 ;
        RECT 340.590 395.720 341.590 398.810 ;
        RECT 342.430 395.720 343.890 398.810 ;
        RECT 344.730 395.720 346.190 398.810 ;
        RECT 347.030 395.720 348.490 398.810 ;
        RECT 349.330 395.720 350.330 398.810 ;
        RECT 351.170 395.720 352.630 398.810 ;
        RECT 353.470 395.720 354.930 398.810 ;
        RECT 355.770 395.720 357.230 398.810 ;
        RECT 358.070 395.720 359.070 398.810 ;
        RECT 359.910 395.720 361.370 398.810 ;
        RECT 362.210 395.720 363.670 398.810 ;
        RECT 364.510 395.720 365.510 398.810 ;
        RECT 366.350 395.720 367.810 398.810 ;
        RECT 368.650 395.720 370.110 398.810 ;
        RECT 370.950 395.720 372.410 398.810 ;
        RECT 373.250 395.720 374.250 398.810 ;
        RECT 375.090 395.720 376.550 398.810 ;
        RECT 377.390 395.720 378.850 398.810 ;
        RECT 379.690 395.720 381.150 398.810 ;
        RECT 381.990 395.720 382.990 398.810 ;
        RECT 383.830 395.720 385.290 398.810 ;
        RECT 386.130 395.720 387.590 398.810 ;
        RECT 388.430 395.720 389.430 398.810 ;
        RECT 390.270 395.720 391.730 398.810 ;
        RECT 392.570 395.720 394.030 398.810 ;
        RECT 394.870 395.720 396.330 398.810 ;
        RECT 397.170 395.720 398.170 398.810 ;
        RECT 399.010 395.720 400.470 398.810 ;
        RECT 401.310 395.720 402.770 398.810 ;
        RECT 403.610 395.720 405.070 398.810 ;
        RECT 405.910 395.720 406.910 398.810 ;
        RECT 407.750 395.720 409.210 398.810 ;
        RECT 410.050 395.720 411.510 398.810 ;
        RECT 412.350 395.720 413.350 398.810 ;
        RECT 414.190 395.720 415.650 398.810 ;
        RECT 416.490 395.720 417.950 398.810 ;
        RECT 418.790 395.720 420.250 398.810 ;
        RECT 421.090 395.720 422.090 398.810 ;
        RECT 422.930 395.720 424.390 398.810 ;
        RECT 425.230 395.720 426.690 398.810 ;
        RECT 427.530 395.720 428.990 398.810 ;
        RECT 429.830 395.720 430.830 398.810 ;
        RECT 431.670 395.720 433.130 398.810 ;
        RECT 433.970 395.720 435.430 398.810 ;
        RECT 436.270 395.720 437.270 398.810 ;
        RECT 438.110 395.720 439.570 398.810 ;
        RECT 440.410 395.720 441.870 398.810 ;
        RECT 442.710 395.720 444.170 398.810 ;
        RECT 445.010 395.720 446.010 398.810 ;
        RECT 446.850 395.720 448.310 398.810 ;
        RECT 449.150 395.720 450.610 398.810 ;
        RECT 451.450 395.720 452.910 398.810 ;
        RECT 453.750 395.720 454.750 398.810 ;
        RECT 455.590 395.720 457.050 398.810 ;
        RECT 457.890 395.720 459.350 398.810 ;
        RECT 460.190 395.720 461.190 398.810 ;
        RECT 462.030 395.720 463.490 398.810 ;
        RECT 464.330 395.720 465.790 398.810 ;
        RECT 466.630 395.720 468.090 398.810 ;
        RECT 468.930 395.720 469.930 398.810 ;
        RECT 470.770 395.720 472.230 398.810 ;
        RECT 473.070 395.720 474.530 398.810 ;
        RECT 475.370 395.720 476.830 398.810 ;
        RECT 477.670 395.720 478.670 398.810 ;
        RECT 479.510 395.720 480.970 398.810 ;
        RECT 481.810 395.720 483.270 398.810 ;
        RECT 484.110 395.720 485.110 398.810 ;
        RECT 485.950 395.720 487.410 398.810 ;
        RECT 488.250 395.720 489.710 398.810 ;
        RECT 490.550 395.720 492.010 398.810 ;
        RECT 492.850 395.720 493.850 398.810 ;
        RECT 494.690 395.720 496.150 398.810 ;
        RECT 496.990 395.720 498.450 398.810 ;
        RECT 499.290 395.720 500.750 398.810 ;
        RECT 501.590 395.720 502.590 398.810 ;
        RECT 503.430 395.720 504.890 398.810 ;
        RECT 505.730 395.720 507.190 398.810 ;
        RECT 508.030 395.720 509.030 398.810 ;
        RECT 509.870 395.720 511.330 398.810 ;
        RECT 512.170 395.720 513.630 398.810 ;
        RECT 514.470 395.720 515.930 398.810 ;
        RECT 516.770 395.720 517.770 398.810 ;
        RECT 518.610 395.720 520.070 398.810 ;
        RECT 520.910 395.720 522.370 398.810 ;
        RECT 523.210 395.720 524.210 398.810 ;
        RECT 525.050 395.720 526.510 398.810 ;
        RECT 527.350 395.720 528.810 398.810 ;
        RECT 529.650 395.720 531.110 398.810 ;
        RECT 531.950 395.720 532.950 398.810 ;
        RECT 533.790 395.720 535.250 398.810 ;
        RECT 536.090 395.720 537.550 398.810 ;
        RECT 538.390 395.720 539.850 398.810 ;
        RECT 540.690 395.720 541.690 398.810 ;
        RECT 542.530 395.720 543.990 398.810 ;
        RECT 544.830 395.720 546.290 398.810 ;
        RECT 547.130 395.720 548.130 398.810 ;
        RECT 548.970 395.720 550.430 398.810 ;
        RECT 551.270 395.720 552.730 398.810 ;
        RECT 553.570 395.720 555.030 398.810 ;
        RECT 555.870 395.720 556.870 398.810 ;
        RECT 557.710 395.720 559.170 398.810 ;
        RECT 560.010 395.720 561.470 398.810 ;
        RECT 562.310 395.720 563.770 398.810 ;
        RECT 564.610 395.720 565.610 398.810 ;
        RECT 566.450 395.720 567.910 398.810 ;
        RECT 568.750 395.720 570.210 398.810 ;
        RECT 571.050 395.720 572.050 398.810 ;
        RECT 572.890 395.720 574.350 398.810 ;
        RECT 575.190 395.720 576.650 398.810 ;
        RECT 577.490 395.720 578.950 398.810 ;
        RECT 579.790 395.720 580.790 398.810 ;
        RECT 581.630 395.720 583.090 398.810 ;
        RECT 583.930 395.720 585.390 398.810 ;
        RECT 586.230 395.720 587.690 398.810 ;
        RECT 588.530 395.720 589.530 398.810 ;
        RECT 590.370 395.720 591.830 398.810 ;
        RECT 592.670 395.720 594.130 398.810 ;
        RECT 594.970 395.720 595.970 398.810 ;
        RECT 596.810 395.720 598.270 398.810 ;
        RECT 599.110 395.720 600.570 398.810 ;
        RECT 601.410 395.720 602.870 398.810 ;
        RECT 603.710 395.720 604.710 398.810 ;
        RECT 605.550 395.720 607.010 398.810 ;
        RECT 607.850 395.720 609.310 398.810 ;
        RECT 610.150 395.720 611.610 398.810 ;
        RECT 612.450 395.720 613.450 398.810 ;
        RECT 614.290 395.720 615.750 398.810 ;
        RECT 616.590 395.720 618.050 398.810 ;
        RECT 618.890 395.720 619.890 398.810 ;
        RECT 620.730 395.720 622.190 398.810 ;
        RECT 623.030 395.720 624.490 398.810 ;
        RECT 625.330 395.720 626.790 398.810 ;
        RECT 627.630 395.720 628.630 398.810 ;
        RECT 629.470 395.720 630.930 398.810 ;
        RECT 631.770 395.720 633.230 398.810 ;
        RECT 634.070 395.720 635.530 398.810 ;
        RECT 636.370 395.720 637.370 398.810 ;
        RECT 638.210 395.720 639.670 398.810 ;
        RECT 640.510 395.720 641.970 398.810 ;
        RECT 642.810 395.720 643.810 398.810 ;
        RECT 644.650 395.720 646.110 398.810 ;
        RECT 646.950 395.720 648.410 398.810 ;
        RECT 649.250 395.720 650.710 398.810 ;
        RECT 651.550 395.720 652.550 398.810 ;
        RECT 653.390 395.720 654.850 398.810 ;
        RECT 655.690 395.720 657.150 398.810 ;
        RECT 657.990 395.720 659.450 398.810 ;
        RECT 660.290 395.720 661.290 398.810 ;
        RECT 662.130 395.720 663.590 398.810 ;
        RECT 664.430 395.720 665.890 398.810 ;
        RECT 666.730 395.720 667.730 398.810 ;
        RECT 668.570 395.720 670.030 398.810 ;
        RECT 670.870 395.720 672.330 398.810 ;
        RECT 673.170 395.720 674.630 398.810 ;
        RECT 675.470 395.720 676.470 398.810 ;
        RECT 677.310 395.720 678.770 398.810 ;
        RECT 679.610 395.720 681.070 398.810 ;
        RECT 681.910 395.720 682.910 398.810 ;
        RECT 683.750 395.720 685.210 398.810 ;
        RECT 686.050 395.720 687.510 398.810 ;
        RECT 688.350 395.720 689.810 398.810 ;
        RECT 690.650 395.720 691.650 398.810 ;
        RECT 692.490 395.720 693.950 398.810 ;
        RECT 694.790 395.720 696.250 398.810 ;
        RECT 697.090 395.720 698.550 398.810 ;
        RECT 699.390 395.720 700.390 398.810 ;
        RECT 701.230 395.720 702.690 398.810 ;
        RECT 703.530 395.720 704.990 398.810 ;
        RECT 705.830 395.720 706.830 398.810 ;
        RECT 707.670 395.720 709.130 398.810 ;
        RECT 709.970 395.720 711.430 398.810 ;
        RECT 712.270 395.720 713.730 398.810 ;
        RECT 714.570 395.720 715.570 398.810 ;
        RECT 716.410 395.720 717.870 398.810 ;
        RECT 718.710 395.720 720.170 398.810 ;
        RECT 721.010 395.720 722.470 398.810 ;
        RECT 723.310 395.720 724.310 398.810 ;
        RECT 725.150 395.720 726.610 398.810 ;
        RECT 727.450 395.720 728.910 398.810 ;
        RECT 729.750 395.720 730.750 398.810 ;
        RECT 731.590 395.720 733.050 398.810 ;
        RECT 733.890 395.720 735.350 398.810 ;
        RECT 736.190 395.720 737.650 398.810 ;
        RECT 738.490 395.720 739.490 398.810 ;
        RECT 740.330 395.720 741.790 398.810 ;
        RECT 742.630 395.720 744.090 398.810 ;
        RECT 744.930 395.720 746.390 398.810 ;
        RECT 747.230 395.720 748.230 398.810 ;
        RECT 749.070 395.720 750.530 398.810 ;
        RECT 751.370 395.720 752.830 398.810 ;
        RECT 753.670 395.720 754.670 398.810 ;
        RECT 755.510 395.720 756.970 398.810 ;
        RECT 757.810 395.720 759.270 398.810 ;
        RECT 760.110 395.720 761.570 398.810 ;
        RECT 762.410 395.720 763.410 398.810 ;
        RECT 764.250 395.720 765.710 398.810 ;
        RECT 766.550 395.720 768.010 398.810 ;
        RECT 768.850 395.720 770.310 398.810 ;
        RECT 771.150 395.720 772.150 398.810 ;
        RECT 772.990 395.720 774.450 398.810 ;
        RECT 775.290 395.720 776.750 398.810 ;
        RECT 777.590 395.720 778.590 398.810 ;
        RECT 779.430 395.720 780.890 398.810 ;
        RECT 781.730 395.720 783.190 398.810 ;
        RECT 784.030 395.720 785.490 398.810 ;
        RECT 786.330 395.720 787.330 398.810 ;
        RECT 788.170 395.720 789.630 398.810 ;
        RECT 790.470 395.720 791.930 398.810 ;
        RECT 792.770 395.720 794.230 398.810 ;
        RECT 795.070 395.720 796.070 398.810 ;
        RECT 796.910 395.720 798.370 398.810 ;
        RECT 799.210 395.720 800.670 398.810 ;
        RECT 801.510 395.720 802.510 398.810 ;
        RECT 803.350 395.720 804.810 398.810 ;
        RECT 805.650 395.720 807.110 398.810 ;
        RECT 807.950 395.720 809.410 398.810 ;
        RECT 810.250 395.720 811.250 398.810 ;
        RECT 812.090 395.720 813.550 398.810 ;
        RECT 814.390 395.720 815.850 398.810 ;
        RECT 816.690 395.720 818.150 398.810 ;
        RECT 818.990 395.720 819.990 398.810 ;
        RECT 820.830 395.720 822.290 398.810 ;
        RECT 823.130 395.720 824.590 398.810 ;
        RECT 825.430 395.720 826.430 398.810 ;
        RECT 827.270 395.720 828.730 398.810 ;
        RECT 829.570 395.720 831.030 398.810 ;
        RECT 831.870 395.720 833.330 398.810 ;
        RECT 834.170 395.720 835.170 398.810 ;
        RECT 836.010 395.720 837.470 398.810 ;
        RECT 838.310 395.720 839.770 398.810 ;
        RECT 840.610 395.720 841.610 398.810 ;
        RECT 842.450 395.720 843.910 398.810 ;
        RECT 844.750 395.720 846.210 398.810 ;
        RECT 847.050 395.720 848.510 398.810 ;
        RECT 849.350 395.720 850.350 398.810 ;
        RECT 851.190 395.720 852.650 398.810 ;
        RECT 853.490 395.720 854.950 398.810 ;
        RECT 855.790 395.720 857.250 398.810 ;
        RECT 858.090 395.720 859.090 398.810 ;
        RECT 859.930 395.720 861.390 398.810 ;
        RECT 862.230 395.720 863.690 398.810 ;
        RECT 864.530 395.720 865.530 398.810 ;
        RECT 866.370 395.720 867.830 398.810 ;
        RECT 868.670 395.720 870.130 398.810 ;
        RECT 870.970 395.720 872.430 398.810 ;
        RECT 873.270 395.720 874.270 398.810 ;
        RECT 875.110 395.720 876.570 398.810 ;
        RECT 877.410 395.720 878.870 398.810 ;
        RECT 879.710 395.720 881.170 398.810 ;
        RECT 882.010 395.720 883.010 398.810 ;
        RECT 883.850 395.720 885.310 398.810 ;
        RECT 886.150 395.720 887.610 398.810 ;
        RECT 888.450 395.720 889.450 398.810 ;
        RECT 890.290 395.720 891.750 398.810 ;
        RECT 892.590 395.720 894.050 398.810 ;
        RECT 894.890 395.720 896.350 398.810 ;
        RECT 897.190 395.720 898.190 398.810 ;
        RECT 899.030 395.720 900.490 398.810 ;
        RECT 901.330 395.720 902.790 398.810 ;
        RECT 903.630 395.720 905.090 398.810 ;
        RECT 905.930 395.720 906.930 398.810 ;
        RECT 907.770 395.720 909.230 398.810 ;
        RECT 910.070 395.720 911.530 398.810 ;
        RECT 912.370 395.720 913.370 398.810 ;
        RECT 914.210 395.720 915.670 398.810 ;
        RECT 916.510 395.720 917.970 398.810 ;
        RECT 918.810 395.720 920.270 398.810 ;
        RECT 921.110 395.720 922.110 398.810 ;
        RECT 922.950 395.720 924.410 398.810 ;
        RECT 925.250 395.720 926.710 398.810 ;
        RECT 927.550 395.720 929.010 398.810 ;
        RECT 929.850 395.720 930.850 398.810 ;
        RECT 931.690 395.720 933.150 398.810 ;
        RECT 933.990 395.720 935.450 398.810 ;
        RECT 936.290 395.720 937.290 398.810 ;
        RECT 938.130 395.720 939.590 398.810 ;
        RECT 940.430 395.720 941.890 398.810 ;
        RECT 942.730 395.720 944.190 398.810 ;
        RECT 945.030 395.720 946.030 398.810 ;
        RECT 946.870 395.720 948.330 398.810 ;
        RECT 949.170 395.720 950.630 398.810 ;
        RECT 951.470 395.720 952.930 398.810 ;
        RECT 953.770 395.720 954.770 398.810 ;
        RECT 955.610 395.720 957.070 398.810 ;
        RECT 957.910 395.720 959.370 398.810 ;
        RECT 960.210 395.720 961.210 398.810 ;
        RECT 962.050 395.720 963.510 398.810 ;
        RECT 964.350 395.720 965.810 398.810 ;
        RECT 966.650 395.720 968.110 398.810 ;
        RECT 968.950 395.720 969.950 398.810 ;
        RECT 970.790 395.720 972.250 398.810 ;
        RECT 973.090 395.720 974.550 398.810 ;
        RECT 975.390 395.720 976.850 398.810 ;
        RECT 977.690 395.720 978.690 398.810 ;
        RECT 979.530 395.720 980.990 398.810 ;
        RECT 981.830 395.720 983.290 398.810 ;
        RECT 984.130 395.720 985.130 398.810 ;
        RECT 985.970 395.720 987.430 398.810 ;
        RECT 988.270 395.720 989.730 398.810 ;
        RECT 990.570 395.720 992.030 398.810 ;
        RECT 992.870 395.720 993.870 398.810 ;
        RECT 994.710 395.720 996.170 398.810 ;
        RECT 997.010 395.720 998.470 398.810 ;
        RECT 999.310 395.720 1000.770 398.810 ;
        RECT 1001.610 395.720 1002.610 398.810 ;
        RECT 1003.450 395.720 1004.910 398.810 ;
        RECT 1005.750 395.720 1007.210 398.810 ;
        RECT 1008.050 395.720 1009.050 398.810 ;
        RECT 1009.890 395.720 1011.350 398.810 ;
        RECT 1012.190 395.720 1013.650 398.810 ;
        RECT 1014.490 395.720 1015.950 398.810 ;
        RECT 1016.790 395.720 1017.790 398.810 ;
        RECT 1018.630 395.720 1020.090 398.810 ;
        RECT 1020.930 395.720 1022.390 398.810 ;
        RECT 1023.230 395.720 1024.230 398.810 ;
        RECT 1025.070 395.720 1026.530 398.810 ;
        RECT 1027.370 395.720 1028.830 398.810 ;
        RECT 1029.670 395.720 1031.130 398.810 ;
        RECT 1031.970 395.720 1032.970 398.810 ;
        RECT 1033.810 395.720 1035.270 398.810 ;
        RECT 1036.110 395.720 1037.570 398.810 ;
        RECT 1038.410 395.720 1039.870 398.810 ;
        RECT 1040.710 395.720 1041.710 398.810 ;
        RECT 1042.550 395.720 1044.010 398.810 ;
        RECT 1044.850 395.720 1046.310 398.810 ;
        RECT 1047.150 395.720 1048.150 398.810 ;
        RECT 1048.990 395.720 1050.450 398.810 ;
        RECT 1051.290 395.720 1052.750 398.810 ;
        RECT 1053.590 395.720 1055.050 398.810 ;
        RECT 1055.890 395.720 1056.890 398.810 ;
        RECT 1057.730 395.720 1059.190 398.810 ;
        RECT 1060.030 395.720 1061.490 398.810 ;
        RECT 1062.330 395.720 1063.790 398.810 ;
        RECT 1064.630 395.720 1065.630 398.810 ;
        RECT 1066.470 395.720 1067.930 398.810 ;
        RECT 1068.770 395.720 1070.230 398.810 ;
        RECT 1071.070 395.720 1072.070 398.810 ;
        RECT 1072.910 395.720 1074.370 398.810 ;
        RECT 1075.210 395.720 1076.670 398.810 ;
        RECT 1077.510 395.720 1078.970 398.810 ;
        RECT 1079.810 395.720 1080.810 398.810 ;
        RECT 1081.650 395.720 1083.110 398.810 ;
        RECT 1083.950 395.720 1085.410 398.810 ;
        RECT 1086.250 395.720 1087.710 398.810 ;
        RECT 1088.550 395.720 1089.550 398.810 ;
        RECT 1090.390 395.720 1091.850 398.810 ;
        RECT 1092.690 395.720 1094.150 398.810 ;
        RECT 1094.990 395.720 1095.990 398.810 ;
        RECT 1096.830 395.720 1098.290 398.810 ;
        RECT 1099.130 395.720 1100.590 398.810 ;
        RECT 1101.430 395.720 1102.890 398.810 ;
        RECT 1103.730 395.720 1104.730 398.810 ;
        RECT 1105.570 395.720 1107.030 398.810 ;
        RECT 1107.870 395.720 1109.330 398.810 ;
        RECT 1110.170 395.720 1111.630 398.810 ;
        RECT 1112.470 395.720 1113.470 398.810 ;
        RECT 1114.310 395.720 1115.770 398.810 ;
        RECT 1116.610 395.720 1118.070 398.810 ;
        RECT 1118.910 395.720 1119.910 398.810 ;
        RECT 1120.750 395.720 1122.210 398.810 ;
        RECT 1123.050 395.720 1124.510 398.810 ;
        RECT 1125.350 395.720 1126.810 398.810 ;
        RECT 1127.650 395.720 1128.650 398.810 ;
        RECT 1129.490 395.720 1130.950 398.810 ;
        RECT 1131.790 395.720 1133.250 398.810 ;
        RECT 1134.090 395.720 1135.550 398.810 ;
        RECT 1136.390 395.720 1137.390 398.810 ;
        RECT 1138.230 395.720 1139.690 398.810 ;
        RECT 1140.530 395.720 1141.990 398.810 ;
        RECT 1142.830 395.720 1143.830 398.810 ;
        RECT 1144.670 395.720 1146.130 398.810 ;
        RECT 1146.970 395.720 1148.430 398.810 ;
        RECT 1149.270 395.720 1150.730 398.810 ;
        RECT 1151.570 395.720 1152.570 398.810 ;
        RECT 1153.410 395.720 1154.870 398.810 ;
        RECT 1155.710 395.720 1157.170 398.810 ;
        RECT 1158.010 395.720 1159.470 398.810 ;
        RECT 1160.310 395.720 1161.310 398.810 ;
        RECT 1162.150 395.720 1163.610 398.810 ;
        RECT 1164.450 395.720 1165.910 398.810 ;
        RECT 1166.750 395.720 1167.750 398.810 ;
        RECT 1168.590 395.720 1170.050 398.810 ;
        RECT 1170.890 395.720 1172.350 398.810 ;
        RECT 1173.190 395.720 1174.650 398.810 ;
        RECT 1175.490 395.720 1176.490 398.810 ;
        RECT 1177.330 395.720 1178.790 398.810 ;
        RECT 1179.630 395.720 1181.090 398.810 ;
        RECT 1181.930 395.720 1182.930 398.810 ;
        RECT 1183.770 395.720 1185.230 398.810 ;
        RECT 1186.070 395.720 1187.530 398.810 ;
        RECT 1188.370 395.720 1189.830 398.810 ;
        RECT 1190.670 395.720 1191.670 398.810 ;
        RECT 1192.510 395.720 1193.970 398.810 ;
        RECT 1194.810 395.720 1196.270 398.810 ;
        RECT 1197.110 395.720 1198.570 398.810 ;
        RECT 1199.410 395.720 1200.410 398.810 ;
        RECT 1201.250 395.720 1202.710 398.810 ;
        RECT 1203.550 395.720 1205.010 398.810 ;
        RECT 1205.850 395.720 1206.850 398.810 ;
        RECT 1207.690 395.720 1209.150 398.810 ;
        RECT 1209.990 395.720 1211.450 398.810 ;
        RECT 1212.290 395.720 1213.750 398.810 ;
        RECT 1214.590 395.720 1215.590 398.810 ;
        RECT 1216.430 395.720 1217.890 398.810 ;
        RECT 1218.730 395.720 1220.190 398.810 ;
        RECT 1221.030 395.720 1222.490 398.810 ;
        RECT 1223.330 395.720 1224.330 398.810 ;
        RECT 1225.170 395.720 1226.630 398.810 ;
        RECT 1227.470 395.720 1228.930 398.810 ;
        RECT 1229.770 395.720 1230.770 398.810 ;
        RECT 1231.610 395.720 1233.070 398.810 ;
        RECT 1233.910 395.720 1235.370 398.810 ;
        RECT 1236.210 395.720 1237.670 398.810 ;
        RECT 1238.510 395.720 1239.510 398.810 ;
        RECT 1240.350 395.720 1241.810 398.810 ;
        RECT 1242.650 395.720 1244.110 398.810 ;
        RECT 1244.950 395.720 1246.410 398.810 ;
        RECT 1247.250 395.720 1248.250 398.810 ;
        RECT 1249.090 395.720 1250.550 398.810 ;
        RECT 1251.390 395.720 1252.850 398.810 ;
        RECT 1253.690 395.720 1254.690 398.810 ;
        RECT 1255.530 395.720 1256.990 398.810 ;
        RECT 1257.830 395.720 1259.290 398.810 ;
        RECT 1260.130 395.720 1261.590 398.810 ;
        RECT 1262.430 395.720 1263.430 398.810 ;
        RECT 1264.270 395.720 1265.730 398.810 ;
        RECT 1266.570 395.720 1268.030 398.810 ;
        RECT 1268.870 395.720 1270.330 398.810 ;
        RECT 1271.170 395.720 1272.170 398.810 ;
        RECT 1273.010 395.720 1274.470 398.810 ;
        RECT 1275.310 395.720 1276.770 398.810 ;
        RECT 1277.610 395.720 1278.610 398.810 ;
        RECT 1279.450 395.720 1280.910 398.810 ;
        RECT 1281.750 395.720 1283.210 398.810 ;
        RECT 1284.050 395.720 1285.510 398.810 ;
        RECT 1286.350 395.720 1287.350 398.810 ;
        RECT 1288.190 395.720 1289.650 398.810 ;
        RECT 1290.490 395.720 1291.950 398.810 ;
        RECT 1292.790 395.720 1294.250 398.810 ;
        RECT 1295.090 395.720 1296.090 398.810 ;
        RECT 1296.930 395.720 1298.390 398.810 ;
        RECT 1299.230 395.720 1300.690 398.810 ;
        RECT 1301.530 395.720 1302.530 398.810 ;
        RECT 1303.370 395.720 1304.830 398.810 ;
        RECT 1305.670 395.720 1307.130 398.810 ;
        RECT 1307.970 395.720 1309.430 398.810 ;
        RECT 1310.270 395.720 1311.270 398.810 ;
        RECT 1312.110 395.720 1313.570 398.810 ;
        RECT 1314.410 395.720 1315.870 398.810 ;
        RECT 1316.710 395.720 1318.170 398.810 ;
        RECT 1319.010 395.720 1320.010 398.810 ;
        RECT 1320.850 395.720 1322.310 398.810 ;
        RECT 1323.150 395.720 1324.610 398.810 ;
        RECT 1325.450 395.720 1326.450 398.810 ;
        RECT 1327.290 395.720 1328.750 398.810 ;
        RECT 1329.590 395.720 1331.050 398.810 ;
        RECT 1331.890 395.720 1333.350 398.810 ;
        RECT 1334.190 395.720 1335.190 398.810 ;
        RECT 1336.030 395.720 1337.490 398.810 ;
        RECT 1338.330 395.720 1339.790 398.810 ;
        RECT 1340.630 395.720 1341.630 398.810 ;
        RECT 1342.470 395.720 1343.930 398.810 ;
        RECT 1344.770 395.720 1346.230 398.810 ;
        RECT 1347.070 395.720 1348.530 398.810 ;
        RECT 1349.370 395.720 1350.370 398.810 ;
        RECT 1351.210 395.720 1352.670 398.810 ;
        RECT 1353.510 395.720 1354.970 398.810 ;
        RECT 1355.810 395.720 1357.270 398.810 ;
        RECT 1358.110 395.720 1359.110 398.810 ;
        RECT 1359.950 395.720 1361.410 398.810 ;
        RECT 1362.250 395.720 1363.710 398.810 ;
        RECT 1364.550 395.720 1365.550 398.810 ;
        RECT 1366.390 395.720 1367.850 398.810 ;
        RECT 1368.690 395.720 1370.150 398.810 ;
        RECT 1370.990 395.720 1372.450 398.810 ;
        RECT 1373.290 395.720 1374.290 398.810 ;
        RECT 1375.130 395.720 1376.590 398.810 ;
        RECT 1377.430 395.720 1378.890 398.810 ;
        RECT 1379.730 395.720 1381.190 398.810 ;
        RECT 1382.030 395.720 1383.030 398.810 ;
        RECT 1383.870 395.720 1385.330 398.810 ;
        RECT 1386.170 395.720 1387.630 398.810 ;
        RECT 1388.470 395.720 1389.470 398.810 ;
        RECT 1390.310 395.720 1391.770 398.810 ;
        RECT 1392.610 395.720 1394.070 398.810 ;
        RECT 1394.910 395.720 1396.370 398.810 ;
        RECT 1397.210 395.720 1398.210 398.810 ;
        RECT 1399.050 395.720 1400.510 398.810 ;
        RECT 1401.350 395.720 1402.810 398.810 ;
        RECT 1403.650 395.720 1405.110 398.810 ;
        RECT 1405.950 395.720 1406.950 398.810 ;
        RECT 1407.790 395.720 1409.250 398.810 ;
        RECT 1410.090 395.720 1411.550 398.810 ;
        RECT 1412.390 395.720 1413.390 398.810 ;
        RECT 1414.230 395.720 1415.690 398.810 ;
        RECT 1416.530 395.720 1417.990 398.810 ;
        RECT 1418.830 395.720 1420.290 398.810 ;
        RECT 1421.130 395.720 1422.130 398.810 ;
        RECT 1422.970 395.720 1424.430 398.810 ;
        RECT 1425.270 395.720 1426.730 398.810 ;
        RECT 1427.570 395.720 1429.030 398.810 ;
        RECT 1429.870 395.720 1430.870 398.810 ;
        RECT 1431.710 395.720 1433.170 398.810 ;
        RECT 1434.010 395.720 1435.470 398.810 ;
        RECT 1436.310 395.720 1437.310 398.810 ;
        RECT 1438.150 395.720 1439.610 398.810 ;
        RECT 1440.450 395.720 1441.910 398.810 ;
        RECT 1442.750 395.720 1444.210 398.810 ;
        RECT 1445.050 395.720 1446.050 398.810 ;
        RECT 1446.890 395.720 1448.350 398.810 ;
        RECT 1449.190 395.720 1450.650 398.810 ;
        RECT 1451.490 395.720 1452.950 398.810 ;
        RECT 1453.790 395.720 1454.790 398.810 ;
        RECT 1455.630 395.720 1457.090 398.810 ;
        RECT 1457.930 395.720 1459.390 398.810 ;
        RECT 1460.230 395.720 1461.230 398.810 ;
        RECT 1462.070 395.720 1463.530 398.810 ;
        RECT 1464.370 395.720 1465.830 398.810 ;
        RECT 1466.670 395.720 1468.130 398.810 ;
        RECT 1468.970 395.720 1469.970 398.810 ;
        RECT 1470.810 395.720 1472.270 398.810 ;
        RECT 1473.110 395.720 1474.570 398.810 ;
        RECT 1475.410 395.720 1476.870 398.810 ;
        RECT 1477.710 395.720 1478.710 398.810 ;
        RECT 1479.550 395.720 1481.010 398.810 ;
        RECT 1481.850 395.720 1483.310 398.810 ;
        RECT 1484.150 395.720 1485.150 398.810 ;
        RECT 1485.990 395.720 1487.450 398.810 ;
        RECT 1488.290 395.720 1489.750 398.810 ;
        RECT 1490.590 395.720 1492.050 398.810 ;
        RECT 1492.890 395.720 1493.890 398.810 ;
        RECT 1494.730 395.720 1496.190 398.810 ;
        RECT 1497.030 395.720 1498.490 398.810 ;
        RECT 1.020 4.280 1499.040 395.720 ;
        RECT 1.020 2.195 1.190 4.280 ;
        RECT 2.030 2.195 3.950 4.280 ;
        RECT 4.790 2.195 7.170 4.280 ;
        RECT 8.010 2.195 9.930 4.280 ;
        RECT 10.770 2.195 13.150 4.280 ;
        RECT 13.990 2.195 16.370 4.280 ;
        RECT 17.210 2.195 19.130 4.280 ;
        RECT 19.970 2.195 22.350 4.280 ;
        RECT 23.190 2.195 25.570 4.280 ;
        RECT 26.410 2.195 28.330 4.280 ;
        RECT 29.170 2.195 31.550 4.280 ;
        RECT 32.390 2.195 34.770 4.280 ;
        RECT 35.610 2.195 37.530 4.280 ;
        RECT 38.370 2.195 40.750 4.280 ;
        RECT 41.590 2.195 43.970 4.280 ;
        RECT 44.810 2.195 46.730 4.280 ;
        RECT 47.570 2.195 49.950 4.280 ;
        RECT 50.790 2.195 53.170 4.280 ;
        RECT 54.010 2.195 55.930 4.280 ;
        RECT 56.770 2.195 59.150 4.280 ;
        RECT 59.990 2.195 62.370 4.280 ;
        RECT 63.210 2.195 65.130 4.280 ;
        RECT 65.970 2.195 68.350 4.280 ;
        RECT 69.190 2.195 71.570 4.280 ;
        RECT 72.410 2.195 74.330 4.280 ;
        RECT 75.170 2.195 77.550 4.280 ;
        RECT 78.390 2.195 80.770 4.280 ;
        RECT 81.610 2.195 83.530 4.280 ;
        RECT 84.370 2.195 86.750 4.280 ;
        RECT 87.590 2.195 89.510 4.280 ;
        RECT 90.350 2.195 92.730 4.280 ;
        RECT 93.570 2.195 95.950 4.280 ;
        RECT 96.790 2.195 98.710 4.280 ;
        RECT 99.550 2.195 101.930 4.280 ;
        RECT 102.770 2.195 105.150 4.280 ;
        RECT 105.990 2.195 107.910 4.280 ;
        RECT 108.750 2.195 111.130 4.280 ;
        RECT 111.970 2.195 114.350 4.280 ;
        RECT 115.190 2.195 117.110 4.280 ;
        RECT 117.950 2.195 120.330 4.280 ;
        RECT 121.170 2.195 123.550 4.280 ;
        RECT 124.390 2.195 126.310 4.280 ;
        RECT 127.150 2.195 129.530 4.280 ;
        RECT 130.370 2.195 132.750 4.280 ;
        RECT 133.590 2.195 135.510 4.280 ;
        RECT 136.350 2.195 138.730 4.280 ;
        RECT 139.570 2.195 141.950 4.280 ;
        RECT 142.790 2.195 144.710 4.280 ;
        RECT 145.550 2.195 147.930 4.280 ;
        RECT 148.770 2.195 151.150 4.280 ;
        RECT 151.990 2.195 153.910 4.280 ;
        RECT 154.750 2.195 157.130 4.280 ;
        RECT 157.970 2.195 160.350 4.280 ;
        RECT 161.190 2.195 163.110 4.280 ;
        RECT 163.950 2.195 166.330 4.280 ;
        RECT 167.170 2.195 169.550 4.280 ;
        RECT 170.390 2.195 172.310 4.280 ;
        RECT 173.150 2.195 175.530 4.280 ;
        RECT 176.370 2.195 178.290 4.280 ;
        RECT 179.130 2.195 181.510 4.280 ;
        RECT 182.350 2.195 184.730 4.280 ;
        RECT 185.570 2.195 187.490 4.280 ;
        RECT 188.330 2.195 190.710 4.280 ;
        RECT 191.550 2.195 193.930 4.280 ;
        RECT 194.770 2.195 196.690 4.280 ;
        RECT 197.530 2.195 199.910 4.280 ;
        RECT 200.750 2.195 203.130 4.280 ;
        RECT 203.970 2.195 205.890 4.280 ;
        RECT 206.730 2.195 209.110 4.280 ;
        RECT 209.950 2.195 212.330 4.280 ;
        RECT 213.170 2.195 215.090 4.280 ;
        RECT 215.930 2.195 218.310 4.280 ;
        RECT 219.150 2.195 221.530 4.280 ;
        RECT 222.370 2.195 224.290 4.280 ;
        RECT 225.130 2.195 227.510 4.280 ;
        RECT 228.350 2.195 230.730 4.280 ;
        RECT 231.570 2.195 233.490 4.280 ;
        RECT 234.330 2.195 236.710 4.280 ;
        RECT 237.550 2.195 239.930 4.280 ;
        RECT 240.770 2.195 242.690 4.280 ;
        RECT 243.530 2.195 245.910 4.280 ;
        RECT 246.750 2.195 249.130 4.280 ;
        RECT 249.970 2.195 251.890 4.280 ;
        RECT 252.730 2.195 255.110 4.280 ;
        RECT 255.950 2.195 258.330 4.280 ;
        RECT 259.170 2.195 261.090 4.280 ;
        RECT 261.930 2.195 264.310 4.280 ;
        RECT 265.150 2.195 267.070 4.280 ;
        RECT 267.910 2.195 270.290 4.280 ;
        RECT 271.130 2.195 273.510 4.280 ;
        RECT 274.350 2.195 276.270 4.280 ;
        RECT 277.110 2.195 279.490 4.280 ;
        RECT 280.330 2.195 282.710 4.280 ;
        RECT 283.550 2.195 285.470 4.280 ;
        RECT 286.310 2.195 288.690 4.280 ;
        RECT 289.530 2.195 291.910 4.280 ;
        RECT 292.750 2.195 294.670 4.280 ;
        RECT 295.510 2.195 297.890 4.280 ;
        RECT 298.730 2.195 301.110 4.280 ;
        RECT 301.950 2.195 303.870 4.280 ;
        RECT 304.710 2.195 307.090 4.280 ;
        RECT 307.930 2.195 310.310 4.280 ;
        RECT 311.150 2.195 313.070 4.280 ;
        RECT 313.910 2.195 316.290 4.280 ;
        RECT 317.130 2.195 319.510 4.280 ;
        RECT 320.350 2.195 322.270 4.280 ;
        RECT 323.110 2.195 325.490 4.280 ;
        RECT 326.330 2.195 328.710 4.280 ;
        RECT 329.550 2.195 331.470 4.280 ;
        RECT 332.310 2.195 334.690 4.280 ;
        RECT 335.530 2.195 337.910 4.280 ;
        RECT 338.750 2.195 340.670 4.280 ;
        RECT 341.510 2.195 343.890 4.280 ;
        RECT 344.730 2.195 347.110 4.280 ;
        RECT 347.950 2.195 349.870 4.280 ;
        RECT 350.710 2.195 353.090 4.280 ;
        RECT 353.930 2.195 355.850 4.280 ;
        RECT 356.690 2.195 359.070 4.280 ;
        RECT 359.910 2.195 362.290 4.280 ;
        RECT 363.130 2.195 365.050 4.280 ;
        RECT 365.890 2.195 368.270 4.280 ;
        RECT 369.110 2.195 371.490 4.280 ;
        RECT 372.330 2.195 374.250 4.280 ;
        RECT 375.090 2.195 377.470 4.280 ;
        RECT 378.310 2.195 380.690 4.280 ;
        RECT 381.530 2.195 383.450 4.280 ;
        RECT 384.290 2.195 386.670 4.280 ;
        RECT 387.510 2.195 389.890 4.280 ;
        RECT 390.730 2.195 392.650 4.280 ;
        RECT 393.490 2.195 395.870 4.280 ;
        RECT 396.710 2.195 399.090 4.280 ;
        RECT 399.930 2.195 401.850 4.280 ;
        RECT 402.690 2.195 405.070 4.280 ;
        RECT 405.910 2.195 408.290 4.280 ;
        RECT 409.130 2.195 411.050 4.280 ;
        RECT 411.890 2.195 414.270 4.280 ;
        RECT 415.110 2.195 417.490 4.280 ;
        RECT 418.330 2.195 420.250 4.280 ;
        RECT 421.090 2.195 423.470 4.280 ;
        RECT 424.310 2.195 426.690 4.280 ;
        RECT 427.530 2.195 429.450 4.280 ;
        RECT 430.290 2.195 432.670 4.280 ;
        RECT 433.510 2.195 435.890 4.280 ;
        RECT 436.730 2.195 438.650 4.280 ;
        RECT 439.490 2.195 441.870 4.280 ;
        RECT 442.710 2.195 444.630 4.280 ;
        RECT 445.470 2.195 447.850 4.280 ;
        RECT 448.690 2.195 451.070 4.280 ;
        RECT 451.910 2.195 453.830 4.280 ;
        RECT 454.670 2.195 457.050 4.280 ;
        RECT 457.890 2.195 460.270 4.280 ;
        RECT 461.110 2.195 463.030 4.280 ;
        RECT 463.870 2.195 466.250 4.280 ;
        RECT 467.090 2.195 469.470 4.280 ;
        RECT 470.310 2.195 472.230 4.280 ;
        RECT 473.070 2.195 475.450 4.280 ;
        RECT 476.290 2.195 478.670 4.280 ;
        RECT 479.510 2.195 481.430 4.280 ;
        RECT 482.270 2.195 484.650 4.280 ;
        RECT 485.490 2.195 487.870 4.280 ;
        RECT 488.710 2.195 490.630 4.280 ;
        RECT 491.470 2.195 493.850 4.280 ;
        RECT 494.690 2.195 497.070 4.280 ;
        RECT 497.910 2.195 499.830 4.280 ;
        RECT 500.670 2.195 503.050 4.280 ;
        RECT 503.890 2.195 506.270 4.280 ;
        RECT 507.110 2.195 509.030 4.280 ;
        RECT 509.870 2.195 512.250 4.280 ;
        RECT 513.090 2.195 515.470 4.280 ;
        RECT 516.310 2.195 518.230 4.280 ;
        RECT 519.070 2.195 521.450 4.280 ;
        RECT 522.290 2.195 524.670 4.280 ;
        RECT 525.510 2.195 527.430 4.280 ;
        RECT 528.270 2.195 530.650 4.280 ;
        RECT 531.490 2.195 533.410 4.280 ;
        RECT 534.250 2.195 536.630 4.280 ;
        RECT 537.470 2.195 539.850 4.280 ;
        RECT 540.690 2.195 542.610 4.280 ;
        RECT 543.450 2.195 545.830 4.280 ;
        RECT 546.670 2.195 549.050 4.280 ;
        RECT 549.890 2.195 551.810 4.280 ;
        RECT 552.650 2.195 555.030 4.280 ;
        RECT 555.870 2.195 558.250 4.280 ;
        RECT 559.090 2.195 561.010 4.280 ;
        RECT 561.850 2.195 564.230 4.280 ;
        RECT 565.070 2.195 567.450 4.280 ;
        RECT 568.290 2.195 570.210 4.280 ;
        RECT 571.050 2.195 573.430 4.280 ;
        RECT 574.270 2.195 576.650 4.280 ;
        RECT 577.490 2.195 579.410 4.280 ;
        RECT 580.250 2.195 582.630 4.280 ;
        RECT 583.470 2.195 585.850 4.280 ;
        RECT 586.690 2.195 588.610 4.280 ;
        RECT 589.450 2.195 591.830 4.280 ;
        RECT 592.670 2.195 595.050 4.280 ;
        RECT 595.890 2.195 597.810 4.280 ;
        RECT 598.650 2.195 601.030 4.280 ;
        RECT 601.870 2.195 604.250 4.280 ;
        RECT 605.090 2.195 607.010 4.280 ;
        RECT 607.850 2.195 610.230 4.280 ;
        RECT 611.070 2.195 613.450 4.280 ;
        RECT 614.290 2.195 616.210 4.280 ;
        RECT 617.050 2.195 619.430 4.280 ;
        RECT 620.270 2.195 622.190 4.280 ;
        RECT 623.030 2.195 625.410 4.280 ;
        RECT 626.250 2.195 628.630 4.280 ;
        RECT 629.470 2.195 631.390 4.280 ;
        RECT 632.230 2.195 634.610 4.280 ;
        RECT 635.450 2.195 637.830 4.280 ;
        RECT 638.670 2.195 640.590 4.280 ;
        RECT 641.430 2.195 643.810 4.280 ;
        RECT 644.650 2.195 647.030 4.280 ;
        RECT 647.870 2.195 649.790 4.280 ;
        RECT 650.630 2.195 653.010 4.280 ;
        RECT 653.850 2.195 656.230 4.280 ;
        RECT 657.070 2.195 658.990 4.280 ;
        RECT 659.830 2.195 662.210 4.280 ;
        RECT 663.050 2.195 665.430 4.280 ;
        RECT 666.270 2.195 668.190 4.280 ;
        RECT 669.030 2.195 671.410 4.280 ;
        RECT 672.250 2.195 674.630 4.280 ;
        RECT 675.470 2.195 677.390 4.280 ;
        RECT 678.230 2.195 680.610 4.280 ;
        RECT 681.450 2.195 683.830 4.280 ;
        RECT 684.670 2.195 686.590 4.280 ;
        RECT 687.430 2.195 689.810 4.280 ;
        RECT 690.650 2.195 693.030 4.280 ;
        RECT 693.870 2.195 695.790 4.280 ;
        RECT 696.630 2.195 699.010 4.280 ;
        RECT 699.850 2.195 702.230 4.280 ;
        RECT 703.070 2.195 704.990 4.280 ;
        RECT 705.830 2.195 708.210 4.280 ;
        RECT 709.050 2.195 710.970 4.280 ;
        RECT 711.810 2.195 714.190 4.280 ;
        RECT 715.030 2.195 717.410 4.280 ;
        RECT 718.250 2.195 720.170 4.280 ;
        RECT 721.010 2.195 723.390 4.280 ;
        RECT 724.230 2.195 726.610 4.280 ;
        RECT 727.450 2.195 729.370 4.280 ;
        RECT 730.210 2.195 732.590 4.280 ;
        RECT 733.430 2.195 735.810 4.280 ;
        RECT 736.650 2.195 738.570 4.280 ;
        RECT 739.410 2.195 741.790 4.280 ;
        RECT 742.630 2.195 745.010 4.280 ;
        RECT 745.850 2.195 747.770 4.280 ;
        RECT 748.610 2.195 750.990 4.280 ;
        RECT 751.830 2.195 754.210 4.280 ;
        RECT 755.050 2.195 756.970 4.280 ;
        RECT 757.810 2.195 760.190 4.280 ;
        RECT 761.030 2.195 763.410 4.280 ;
        RECT 764.250 2.195 766.170 4.280 ;
        RECT 767.010 2.195 769.390 4.280 ;
        RECT 770.230 2.195 772.610 4.280 ;
        RECT 773.450 2.195 775.370 4.280 ;
        RECT 776.210 2.195 778.590 4.280 ;
        RECT 779.430 2.195 781.810 4.280 ;
        RECT 782.650 2.195 784.570 4.280 ;
        RECT 785.410 2.195 787.790 4.280 ;
        RECT 788.630 2.195 791.010 4.280 ;
        RECT 791.850 2.195 793.770 4.280 ;
        RECT 794.610 2.195 796.990 4.280 ;
        RECT 797.830 2.195 799.750 4.280 ;
        RECT 800.590 2.195 802.970 4.280 ;
        RECT 803.810 2.195 806.190 4.280 ;
        RECT 807.030 2.195 808.950 4.280 ;
        RECT 809.790 2.195 812.170 4.280 ;
        RECT 813.010 2.195 815.390 4.280 ;
        RECT 816.230 2.195 818.150 4.280 ;
        RECT 818.990 2.195 821.370 4.280 ;
        RECT 822.210 2.195 824.590 4.280 ;
        RECT 825.430 2.195 827.350 4.280 ;
        RECT 828.190 2.195 830.570 4.280 ;
        RECT 831.410 2.195 833.790 4.280 ;
        RECT 834.630 2.195 836.550 4.280 ;
        RECT 837.390 2.195 839.770 4.280 ;
        RECT 840.610 2.195 842.990 4.280 ;
        RECT 843.830 2.195 845.750 4.280 ;
        RECT 846.590 2.195 848.970 4.280 ;
        RECT 849.810 2.195 852.190 4.280 ;
        RECT 853.030 2.195 854.950 4.280 ;
        RECT 855.790 2.195 858.170 4.280 ;
        RECT 859.010 2.195 861.390 4.280 ;
        RECT 862.230 2.195 864.150 4.280 ;
        RECT 864.990 2.195 867.370 4.280 ;
        RECT 868.210 2.195 870.590 4.280 ;
        RECT 871.430 2.195 873.350 4.280 ;
        RECT 874.190 2.195 876.570 4.280 ;
        RECT 877.410 2.195 879.790 4.280 ;
        RECT 880.630 2.195 882.550 4.280 ;
        RECT 883.390 2.195 885.770 4.280 ;
        RECT 886.610 2.195 888.530 4.280 ;
        RECT 889.370 2.195 891.750 4.280 ;
        RECT 892.590 2.195 894.970 4.280 ;
        RECT 895.810 2.195 897.730 4.280 ;
        RECT 898.570 2.195 900.950 4.280 ;
        RECT 901.790 2.195 904.170 4.280 ;
        RECT 905.010 2.195 906.930 4.280 ;
        RECT 907.770 2.195 910.150 4.280 ;
        RECT 910.990 2.195 913.370 4.280 ;
        RECT 914.210 2.195 916.130 4.280 ;
        RECT 916.970 2.195 919.350 4.280 ;
        RECT 920.190 2.195 922.570 4.280 ;
        RECT 923.410 2.195 925.330 4.280 ;
        RECT 926.170 2.195 928.550 4.280 ;
        RECT 929.390 2.195 931.770 4.280 ;
        RECT 932.610 2.195 934.530 4.280 ;
        RECT 935.370 2.195 937.750 4.280 ;
        RECT 938.590 2.195 940.970 4.280 ;
        RECT 941.810 2.195 943.730 4.280 ;
        RECT 944.570 2.195 946.950 4.280 ;
        RECT 947.790 2.195 950.170 4.280 ;
        RECT 951.010 2.195 952.930 4.280 ;
        RECT 953.770 2.195 956.150 4.280 ;
        RECT 956.990 2.195 959.370 4.280 ;
        RECT 960.210 2.195 962.130 4.280 ;
        RECT 962.970 2.195 965.350 4.280 ;
        RECT 966.190 2.195 968.570 4.280 ;
        RECT 969.410 2.195 971.330 4.280 ;
        RECT 972.170 2.195 974.550 4.280 ;
        RECT 975.390 2.195 977.310 4.280 ;
        RECT 978.150 2.195 980.530 4.280 ;
        RECT 981.370 2.195 983.750 4.280 ;
        RECT 984.590 2.195 986.510 4.280 ;
        RECT 987.350 2.195 989.730 4.280 ;
        RECT 990.570 2.195 992.950 4.280 ;
        RECT 993.790 2.195 995.710 4.280 ;
        RECT 996.550 2.195 998.930 4.280 ;
        RECT 999.770 2.195 1002.150 4.280 ;
        RECT 1002.990 2.195 1004.910 4.280 ;
        RECT 1005.750 2.195 1008.130 4.280 ;
        RECT 1008.970 2.195 1011.350 4.280 ;
        RECT 1012.190 2.195 1014.110 4.280 ;
        RECT 1014.950 2.195 1017.330 4.280 ;
        RECT 1018.170 2.195 1020.550 4.280 ;
        RECT 1021.390 2.195 1023.310 4.280 ;
        RECT 1024.150 2.195 1026.530 4.280 ;
        RECT 1027.370 2.195 1029.750 4.280 ;
        RECT 1030.590 2.195 1032.510 4.280 ;
        RECT 1033.350 2.195 1035.730 4.280 ;
        RECT 1036.570 2.195 1038.950 4.280 ;
        RECT 1039.790 2.195 1041.710 4.280 ;
        RECT 1042.550 2.195 1044.930 4.280 ;
        RECT 1045.770 2.195 1048.150 4.280 ;
        RECT 1048.990 2.195 1050.910 4.280 ;
        RECT 1051.750 2.195 1054.130 4.280 ;
        RECT 1054.970 2.195 1057.350 4.280 ;
        RECT 1058.190 2.195 1060.110 4.280 ;
        RECT 1060.950 2.195 1063.330 4.280 ;
        RECT 1064.170 2.195 1066.090 4.280 ;
        RECT 1066.930 2.195 1069.310 4.280 ;
        RECT 1070.150 2.195 1072.530 4.280 ;
        RECT 1073.370 2.195 1075.290 4.280 ;
        RECT 1076.130 2.195 1078.510 4.280 ;
        RECT 1079.350 2.195 1081.730 4.280 ;
        RECT 1082.570 2.195 1084.490 4.280 ;
        RECT 1085.330 2.195 1087.710 4.280 ;
        RECT 1088.550 2.195 1090.930 4.280 ;
        RECT 1091.770 2.195 1093.690 4.280 ;
        RECT 1094.530 2.195 1096.910 4.280 ;
        RECT 1097.750 2.195 1100.130 4.280 ;
        RECT 1100.970 2.195 1102.890 4.280 ;
        RECT 1103.730 2.195 1106.110 4.280 ;
        RECT 1106.950 2.195 1109.330 4.280 ;
        RECT 1110.170 2.195 1112.090 4.280 ;
        RECT 1112.930 2.195 1115.310 4.280 ;
        RECT 1116.150 2.195 1118.530 4.280 ;
        RECT 1119.370 2.195 1121.290 4.280 ;
        RECT 1122.130 2.195 1124.510 4.280 ;
        RECT 1125.350 2.195 1127.730 4.280 ;
        RECT 1128.570 2.195 1130.490 4.280 ;
        RECT 1131.330 2.195 1133.710 4.280 ;
        RECT 1134.550 2.195 1136.930 4.280 ;
        RECT 1137.770 2.195 1139.690 4.280 ;
        RECT 1140.530 2.195 1142.910 4.280 ;
        RECT 1143.750 2.195 1146.130 4.280 ;
        RECT 1146.970 2.195 1148.890 4.280 ;
        RECT 1149.730 2.195 1152.110 4.280 ;
        RECT 1152.950 2.195 1154.870 4.280 ;
        RECT 1155.710 2.195 1158.090 4.280 ;
        RECT 1158.930 2.195 1161.310 4.280 ;
        RECT 1162.150 2.195 1164.070 4.280 ;
        RECT 1164.910 2.195 1167.290 4.280 ;
        RECT 1168.130 2.195 1170.510 4.280 ;
        RECT 1171.350 2.195 1173.270 4.280 ;
        RECT 1174.110 2.195 1176.490 4.280 ;
        RECT 1177.330 2.195 1179.710 4.280 ;
        RECT 1180.550 2.195 1182.470 4.280 ;
        RECT 1183.310 2.195 1185.690 4.280 ;
        RECT 1186.530 2.195 1188.910 4.280 ;
        RECT 1189.750 2.195 1191.670 4.280 ;
        RECT 1192.510 2.195 1194.890 4.280 ;
        RECT 1195.730 2.195 1198.110 4.280 ;
        RECT 1198.950 2.195 1200.870 4.280 ;
        RECT 1201.710 2.195 1204.090 4.280 ;
        RECT 1204.930 2.195 1207.310 4.280 ;
        RECT 1208.150 2.195 1210.070 4.280 ;
        RECT 1210.910 2.195 1213.290 4.280 ;
        RECT 1214.130 2.195 1216.510 4.280 ;
        RECT 1217.350 2.195 1219.270 4.280 ;
        RECT 1220.110 2.195 1222.490 4.280 ;
        RECT 1223.330 2.195 1225.710 4.280 ;
        RECT 1226.550 2.195 1228.470 4.280 ;
        RECT 1229.310 2.195 1231.690 4.280 ;
        RECT 1232.530 2.195 1234.910 4.280 ;
        RECT 1235.750 2.195 1237.670 4.280 ;
        RECT 1238.510 2.195 1240.890 4.280 ;
        RECT 1241.730 2.195 1243.650 4.280 ;
        RECT 1244.490 2.195 1246.870 4.280 ;
        RECT 1247.710 2.195 1250.090 4.280 ;
        RECT 1250.930 2.195 1252.850 4.280 ;
        RECT 1253.690 2.195 1256.070 4.280 ;
        RECT 1256.910 2.195 1259.290 4.280 ;
        RECT 1260.130 2.195 1262.050 4.280 ;
        RECT 1262.890 2.195 1265.270 4.280 ;
        RECT 1266.110 2.195 1268.490 4.280 ;
        RECT 1269.330 2.195 1271.250 4.280 ;
        RECT 1272.090 2.195 1274.470 4.280 ;
        RECT 1275.310 2.195 1277.690 4.280 ;
        RECT 1278.530 2.195 1280.450 4.280 ;
        RECT 1281.290 2.195 1283.670 4.280 ;
        RECT 1284.510 2.195 1286.890 4.280 ;
        RECT 1287.730 2.195 1289.650 4.280 ;
        RECT 1290.490 2.195 1292.870 4.280 ;
        RECT 1293.710 2.195 1296.090 4.280 ;
        RECT 1296.930 2.195 1298.850 4.280 ;
        RECT 1299.690 2.195 1302.070 4.280 ;
        RECT 1302.910 2.195 1305.290 4.280 ;
        RECT 1306.130 2.195 1308.050 4.280 ;
        RECT 1308.890 2.195 1311.270 4.280 ;
        RECT 1312.110 2.195 1314.490 4.280 ;
        RECT 1315.330 2.195 1317.250 4.280 ;
        RECT 1318.090 2.195 1320.470 4.280 ;
        RECT 1321.310 2.195 1323.690 4.280 ;
        RECT 1324.530 2.195 1326.450 4.280 ;
        RECT 1327.290 2.195 1329.670 4.280 ;
        RECT 1330.510 2.195 1332.430 4.280 ;
        RECT 1333.270 2.195 1335.650 4.280 ;
        RECT 1336.490 2.195 1338.870 4.280 ;
        RECT 1339.710 2.195 1341.630 4.280 ;
        RECT 1342.470 2.195 1344.850 4.280 ;
        RECT 1345.690 2.195 1348.070 4.280 ;
        RECT 1348.910 2.195 1350.830 4.280 ;
        RECT 1351.670 2.195 1354.050 4.280 ;
        RECT 1354.890 2.195 1357.270 4.280 ;
        RECT 1358.110 2.195 1360.030 4.280 ;
        RECT 1360.870 2.195 1363.250 4.280 ;
        RECT 1364.090 2.195 1366.470 4.280 ;
        RECT 1367.310 2.195 1369.230 4.280 ;
        RECT 1370.070 2.195 1372.450 4.280 ;
        RECT 1373.290 2.195 1375.670 4.280 ;
        RECT 1376.510 2.195 1378.430 4.280 ;
        RECT 1379.270 2.195 1381.650 4.280 ;
        RECT 1382.490 2.195 1384.870 4.280 ;
        RECT 1385.710 2.195 1387.630 4.280 ;
        RECT 1388.470 2.195 1390.850 4.280 ;
        RECT 1391.690 2.195 1394.070 4.280 ;
        RECT 1394.910 2.195 1396.830 4.280 ;
        RECT 1397.670 2.195 1400.050 4.280 ;
        RECT 1400.890 2.195 1403.270 4.280 ;
        RECT 1404.110 2.195 1406.030 4.280 ;
        RECT 1406.870 2.195 1409.250 4.280 ;
        RECT 1410.090 2.195 1412.470 4.280 ;
        RECT 1413.310 2.195 1415.230 4.280 ;
        RECT 1416.070 2.195 1418.450 4.280 ;
        RECT 1419.290 2.195 1421.210 4.280 ;
        RECT 1422.050 2.195 1424.430 4.280 ;
        RECT 1425.270 2.195 1427.650 4.280 ;
        RECT 1428.490 2.195 1430.410 4.280 ;
        RECT 1431.250 2.195 1433.630 4.280 ;
        RECT 1434.470 2.195 1436.850 4.280 ;
        RECT 1437.690 2.195 1439.610 4.280 ;
        RECT 1440.450 2.195 1442.830 4.280 ;
        RECT 1443.670 2.195 1446.050 4.280 ;
        RECT 1446.890 2.195 1448.810 4.280 ;
        RECT 1449.650 2.195 1452.030 4.280 ;
        RECT 1452.870 2.195 1455.250 4.280 ;
        RECT 1456.090 2.195 1458.010 4.280 ;
        RECT 1458.850 2.195 1461.230 4.280 ;
        RECT 1462.070 2.195 1464.450 4.280 ;
        RECT 1465.290 2.195 1467.210 4.280 ;
        RECT 1468.050 2.195 1470.430 4.280 ;
        RECT 1471.270 2.195 1473.650 4.280 ;
        RECT 1474.490 2.195 1476.410 4.280 ;
        RECT 1477.250 2.195 1479.630 4.280 ;
        RECT 1480.470 2.195 1482.850 4.280 ;
        RECT 1483.690 2.195 1485.610 4.280 ;
        RECT 1486.450 2.195 1488.830 4.280 ;
        RECT 1489.670 2.195 1492.050 4.280 ;
        RECT 1492.890 2.195 1494.810 4.280 ;
        RECT 1495.650 2.195 1498.030 4.280 ;
        RECT 1498.870 2.195 1499.040 4.280 ;
      LAYER met3 ;
        RECT 4.400 396.080 1496.000 396.945 ;
        RECT 4.000 394.760 1496.000 396.080 ;
        RECT 4.000 393.360 1495.600 394.760 ;
        RECT 4.000 392.040 1496.000 393.360 ;
        RECT 4.400 390.640 1496.000 392.040 ;
        RECT 4.000 386.600 1496.000 390.640 ;
        RECT 4.400 385.200 1496.000 386.600 ;
        RECT 4.000 384.560 1496.000 385.200 ;
        RECT 4.000 383.160 1495.600 384.560 ;
        RECT 4.000 381.840 1496.000 383.160 ;
        RECT 4.400 380.440 1496.000 381.840 ;
        RECT 4.000 376.400 1496.000 380.440 ;
        RECT 4.400 375.000 1496.000 376.400 ;
        RECT 4.000 373.680 1496.000 375.000 ;
        RECT 4.000 372.280 1495.600 373.680 ;
        RECT 4.000 370.960 1496.000 372.280 ;
        RECT 4.400 369.560 1496.000 370.960 ;
        RECT 4.000 365.520 1496.000 369.560 ;
        RECT 4.400 364.120 1496.000 365.520 ;
        RECT 4.000 363.480 1496.000 364.120 ;
        RECT 4.000 362.080 1495.600 363.480 ;
        RECT 4.000 360.760 1496.000 362.080 ;
        RECT 4.400 359.360 1496.000 360.760 ;
        RECT 4.000 355.320 1496.000 359.360 ;
        RECT 4.400 353.920 1496.000 355.320 ;
        RECT 4.000 352.600 1496.000 353.920 ;
        RECT 4.000 351.200 1495.600 352.600 ;
        RECT 4.000 349.880 1496.000 351.200 ;
        RECT 4.400 348.480 1496.000 349.880 ;
        RECT 4.000 344.440 1496.000 348.480 ;
        RECT 4.400 343.040 1496.000 344.440 ;
        RECT 4.000 342.400 1496.000 343.040 ;
        RECT 4.000 341.000 1495.600 342.400 ;
        RECT 4.000 339.680 1496.000 341.000 ;
        RECT 4.400 338.280 1496.000 339.680 ;
        RECT 4.000 334.240 1496.000 338.280 ;
        RECT 4.400 332.840 1496.000 334.240 ;
        RECT 4.000 331.520 1496.000 332.840 ;
        RECT 4.000 330.120 1495.600 331.520 ;
        RECT 4.000 328.800 1496.000 330.120 ;
        RECT 4.400 327.400 1496.000 328.800 ;
        RECT 4.000 323.360 1496.000 327.400 ;
        RECT 4.400 321.960 1496.000 323.360 ;
        RECT 4.000 321.320 1496.000 321.960 ;
        RECT 4.000 319.920 1495.600 321.320 ;
        RECT 4.000 318.600 1496.000 319.920 ;
        RECT 4.400 317.200 1496.000 318.600 ;
        RECT 4.000 313.160 1496.000 317.200 ;
        RECT 4.400 311.760 1496.000 313.160 ;
        RECT 4.000 310.440 1496.000 311.760 ;
        RECT 4.000 309.040 1495.600 310.440 ;
        RECT 4.000 307.720 1496.000 309.040 ;
        RECT 4.400 306.320 1496.000 307.720 ;
        RECT 4.000 302.960 1496.000 306.320 ;
        RECT 4.400 301.560 1496.000 302.960 ;
        RECT 4.000 300.240 1496.000 301.560 ;
        RECT 4.000 298.840 1495.600 300.240 ;
        RECT 4.000 297.520 1496.000 298.840 ;
        RECT 4.400 296.120 1496.000 297.520 ;
        RECT 4.000 292.080 1496.000 296.120 ;
        RECT 4.400 290.680 1496.000 292.080 ;
        RECT 4.000 289.360 1496.000 290.680 ;
        RECT 4.000 287.960 1495.600 289.360 ;
        RECT 4.000 286.640 1496.000 287.960 ;
        RECT 4.400 285.240 1496.000 286.640 ;
        RECT 4.000 281.880 1496.000 285.240 ;
        RECT 4.400 280.480 1496.000 281.880 ;
        RECT 4.000 279.160 1496.000 280.480 ;
        RECT 4.000 277.760 1495.600 279.160 ;
        RECT 4.000 276.440 1496.000 277.760 ;
        RECT 4.400 275.040 1496.000 276.440 ;
        RECT 4.000 271.000 1496.000 275.040 ;
        RECT 4.400 269.600 1496.000 271.000 ;
        RECT 4.000 268.280 1496.000 269.600 ;
        RECT 4.000 266.880 1495.600 268.280 ;
        RECT 4.000 265.560 1496.000 266.880 ;
        RECT 4.400 264.160 1496.000 265.560 ;
        RECT 4.000 260.800 1496.000 264.160 ;
        RECT 4.400 259.400 1496.000 260.800 ;
        RECT 4.000 258.080 1496.000 259.400 ;
        RECT 4.000 256.680 1495.600 258.080 ;
        RECT 4.000 255.360 1496.000 256.680 ;
        RECT 4.400 253.960 1496.000 255.360 ;
        RECT 4.000 249.920 1496.000 253.960 ;
        RECT 4.400 248.520 1496.000 249.920 ;
        RECT 4.000 247.200 1496.000 248.520 ;
        RECT 4.000 245.800 1495.600 247.200 ;
        RECT 4.000 244.480 1496.000 245.800 ;
        RECT 4.400 243.080 1496.000 244.480 ;
        RECT 4.000 239.720 1496.000 243.080 ;
        RECT 4.400 238.320 1496.000 239.720 ;
        RECT 4.000 237.000 1496.000 238.320 ;
        RECT 4.000 235.600 1495.600 237.000 ;
        RECT 4.000 234.280 1496.000 235.600 ;
        RECT 4.400 232.880 1496.000 234.280 ;
        RECT 4.000 228.840 1496.000 232.880 ;
        RECT 4.400 227.440 1496.000 228.840 ;
        RECT 4.000 226.120 1496.000 227.440 ;
        RECT 4.000 224.720 1495.600 226.120 ;
        RECT 4.000 223.400 1496.000 224.720 ;
        RECT 4.400 222.000 1496.000 223.400 ;
        RECT 4.000 218.640 1496.000 222.000 ;
        RECT 4.400 217.240 1496.000 218.640 ;
        RECT 4.000 215.920 1496.000 217.240 ;
        RECT 4.000 214.520 1495.600 215.920 ;
        RECT 4.000 213.200 1496.000 214.520 ;
        RECT 4.400 211.800 1496.000 213.200 ;
        RECT 4.000 207.760 1496.000 211.800 ;
        RECT 4.400 206.360 1496.000 207.760 ;
        RECT 4.000 205.720 1496.000 206.360 ;
        RECT 4.000 204.320 1495.600 205.720 ;
        RECT 4.000 203.000 1496.000 204.320 ;
        RECT 4.400 201.600 1496.000 203.000 ;
        RECT 4.000 197.560 1496.000 201.600 ;
        RECT 4.400 196.160 1496.000 197.560 ;
        RECT 4.000 194.840 1496.000 196.160 ;
        RECT 4.000 193.440 1495.600 194.840 ;
        RECT 4.000 192.120 1496.000 193.440 ;
        RECT 4.400 190.720 1496.000 192.120 ;
        RECT 4.000 186.680 1496.000 190.720 ;
        RECT 4.400 185.280 1496.000 186.680 ;
        RECT 4.000 184.640 1496.000 185.280 ;
        RECT 4.000 183.240 1495.600 184.640 ;
        RECT 4.000 181.920 1496.000 183.240 ;
        RECT 4.400 180.520 1496.000 181.920 ;
        RECT 4.000 176.480 1496.000 180.520 ;
        RECT 4.400 175.080 1496.000 176.480 ;
        RECT 4.000 173.760 1496.000 175.080 ;
        RECT 4.000 172.360 1495.600 173.760 ;
        RECT 4.000 171.040 1496.000 172.360 ;
        RECT 4.400 169.640 1496.000 171.040 ;
        RECT 4.000 165.600 1496.000 169.640 ;
        RECT 4.400 164.200 1496.000 165.600 ;
        RECT 4.000 163.560 1496.000 164.200 ;
        RECT 4.000 162.160 1495.600 163.560 ;
        RECT 4.000 160.840 1496.000 162.160 ;
        RECT 4.400 159.440 1496.000 160.840 ;
        RECT 4.000 155.400 1496.000 159.440 ;
        RECT 4.400 154.000 1496.000 155.400 ;
        RECT 4.000 152.680 1496.000 154.000 ;
        RECT 4.000 151.280 1495.600 152.680 ;
        RECT 4.000 149.960 1496.000 151.280 ;
        RECT 4.400 148.560 1496.000 149.960 ;
        RECT 4.000 144.520 1496.000 148.560 ;
        RECT 4.400 143.120 1496.000 144.520 ;
        RECT 4.000 142.480 1496.000 143.120 ;
        RECT 4.000 141.080 1495.600 142.480 ;
        RECT 4.000 139.760 1496.000 141.080 ;
        RECT 4.400 138.360 1496.000 139.760 ;
        RECT 4.000 134.320 1496.000 138.360 ;
        RECT 4.400 132.920 1496.000 134.320 ;
        RECT 4.000 131.600 1496.000 132.920 ;
        RECT 4.000 130.200 1495.600 131.600 ;
        RECT 4.000 128.880 1496.000 130.200 ;
        RECT 4.400 127.480 1496.000 128.880 ;
        RECT 4.000 123.440 1496.000 127.480 ;
        RECT 4.400 122.040 1496.000 123.440 ;
        RECT 4.000 121.400 1496.000 122.040 ;
        RECT 4.000 120.000 1495.600 121.400 ;
        RECT 4.000 118.680 1496.000 120.000 ;
        RECT 4.400 117.280 1496.000 118.680 ;
        RECT 4.000 113.240 1496.000 117.280 ;
        RECT 4.400 111.840 1496.000 113.240 ;
        RECT 4.000 110.520 1496.000 111.840 ;
        RECT 4.000 109.120 1495.600 110.520 ;
        RECT 4.000 107.800 1496.000 109.120 ;
        RECT 4.400 106.400 1496.000 107.800 ;
        RECT 4.000 103.040 1496.000 106.400 ;
        RECT 4.400 101.640 1496.000 103.040 ;
        RECT 4.000 100.320 1496.000 101.640 ;
        RECT 4.000 98.920 1495.600 100.320 ;
        RECT 4.000 97.600 1496.000 98.920 ;
        RECT 4.400 96.200 1496.000 97.600 ;
        RECT 4.000 92.160 1496.000 96.200 ;
        RECT 4.400 90.760 1496.000 92.160 ;
        RECT 4.000 89.440 1496.000 90.760 ;
        RECT 4.000 88.040 1495.600 89.440 ;
        RECT 4.000 86.720 1496.000 88.040 ;
        RECT 4.400 85.320 1496.000 86.720 ;
        RECT 4.000 81.960 1496.000 85.320 ;
        RECT 4.400 80.560 1496.000 81.960 ;
        RECT 4.000 79.240 1496.000 80.560 ;
        RECT 4.000 77.840 1495.600 79.240 ;
        RECT 4.000 76.520 1496.000 77.840 ;
        RECT 4.400 75.120 1496.000 76.520 ;
        RECT 4.000 71.080 1496.000 75.120 ;
        RECT 4.400 69.680 1496.000 71.080 ;
        RECT 4.000 68.360 1496.000 69.680 ;
        RECT 4.000 66.960 1495.600 68.360 ;
        RECT 4.000 65.640 1496.000 66.960 ;
        RECT 4.400 64.240 1496.000 65.640 ;
        RECT 4.000 60.880 1496.000 64.240 ;
        RECT 4.400 59.480 1496.000 60.880 ;
        RECT 4.000 58.160 1496.000 59.480 ;
        RECT 4.000 56.760 1495.600 58.160 ;
        RECT 4.000 55.440 1496.000 56.760 ;
        RECT 4.400 54.040 1496.000 55.440 ;
        RECT 4.000 50.000 1496.000 54.040 ;
        RECT 4.400 48.600 1496.000 50.000 ;
        RECT 4.000 47.280 1496.000 48.600 ;
        RECT 4.000 45.880 1495.600 47.280 ;
        RECT 4.000 44.560 1496.000 45.880 ;
        RECT 4.400 43.160 1496.000 44.560 ;
        RECT 4.000 39.800 1496.000 43.160 ;
        RECT 4.400 38.400 1496.000 39.800 ;
        RECT 4.000 37.080 1496.000 38.400 ;
        RECT 4.000 35.680 1495.600 37.080 ;
        RECT 4.000 34.360 1496.000 35.680 ;
        RECT 4.400 32.960 1496.000 34.360 ;
        RECT 4.000 28.920 1496.000 32.960 ;
        RECT 4.400 27.520 1496.000 28.920 ;
        RECT 4.000 26.200 1496.000 27.520 ;
        RECT 4.000 24.800 1495.600 26.200 ;
        RECT 4.000 23.480 1496.000 24.800 ;
        RECT 4.400 22.080 1496.000 23.480 ;
        RECT 4.000 18.720 1496.000 22.080 ;
        RECT 4.400 17.320 1496.000 18.720 ;
        RECT 4.000 16.000 1496.000 17.320 ;
        RECT 4.000 14.600 1495.600 16.000 ;
        RECT 4.000 13.280 1496.000 14.600 ;
        RECT 4.400 11.880 1496.000 13.280 ;
        RECT 4.000 7.840 1496.000 11.880 ;
        RECT 4.400 6.440 1496.000 7.840 ;
        RECT 4.000 5.800 1496.000 6.440 ;
        RECT 4.000 4.400 1495.600 5.800 ;
        RECT 4.000 3.080 1496.000 4.400 ;
        RECT 4.400 2.215 1496.000 3.080 ;
      LAYER met4 ;
        RECT 48.135 389.600 1481.840 395.585 ;
        RECT 48.135 10.640 97.440 389.600 ;
        RECT 99.840 10.640 1481.840 389.600 ;
      LAYER met5 ;
        RECT 185.500 344.300 1191.740 383.300 ;
  END
END multi_project_harness
END LIBRARY

