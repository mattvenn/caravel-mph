magic
tech sky130A
magscale 1 2
timestamp 1608298212
<< metal1 >>
rect 133874 700952 133880 701004
rect 133932 700992 133938 701004
rect 218974 700992 218980 701004
rect 133932 700964 218980 700992
rect 133932 700952 133938 700964
rect 218974 700952 218980 700964
rect 219032 700952 219038 701004
rect 235166 700952 235172 701004
rect 235224 700992 235230 701004
rect 434070 700992 434076 701004
rect 235224 700964 434076 700992
rect 235224 700952 235230 700964
rect 434070 700952 434076 700964
rect 434128 700952 434134 701004
rect 133598 700884 133604 700936
rect 133656 700924 133662 700936
rect 348786 700924 348792 700936
rect 133656 700896 348792 700924
rect 133656 700884 133662 700896
rect 348786 700884 348792 700896
rect 348844 700884 348850 700936
rect 364978 700884 364984 700936
rect 365036 700924 365042 700936
rect 433978 700924 433984 700936
rect 365036 700896 433984 700924
rect 365036 700884 365042 700896
rect 433978 700884 433984 700896
rect 434036 700884 434042 700936
rect 133230 700816 133236 700868
rect 133288 700856 133294 700868
rect 397454 700856 397460 700868
rect 133288 700828 397460 700856
rect 133288 700816 133294 700828
rect 397454 700816 397460 700828
rect 397512 700816 397518 700868
rect 132218 700748 132224 700800
rect 132276 700788 132282 700800
rect 154114 700788 154120 700800
rect 132276 700760 154120 700788
rect 132276 700748 132282 700760
rect 154114 700748 154120 700760
rect 154172 700748 154178 700800
rect 170306 700748 170312 700800
rect 170364 700788 170370 700800
rect 434162 700788 434168 700800
rect 170364 700760 434168 700788
rect 170364 700748 170370 700760
rect 434162 700748 434168 700760
rect 434220 700748 434226 700800
rect 131114 700680 131120 700732
rect 131172 700720 131178 700732
rect 413646 700720 413652 700732
rect 131172 700692 413652 700720
rect 131172 700680 131178 700692
rect 413646 700680 413652 700692
rect 413704 700680 413710 700732
rect 105446 700612 105452 700664
rect 105504 700652 105510 700664
rect 434346 700652 434352 700664
rect 105504 700624 434352 700652
rect 105504 700612 105510 700624
rect 434346 700612 434352 700624
rect 434404 700612 434410 700664
rect 438118 700612 438124 700664
rect 438176 700652 438182 700664
rect 494790 700652 494796 700664
rect 438176 700624 494796 700652
rect 438176 700612 438182 700624
rect 494790 700612 494796 700624
rect 494848 700612 494854 700664
rect 133414 700544 133420 700596
rect 133472 700584 133478 700596
rect 462314 700584 462320 700596
rect 133472 700556 462320 700584
rect 133472 700544 133478 700556
rect 462314 700544 462320 700556
rect 462372 700544 462378 700596
rect 133690 700476 133696 700528
rect 133748 700516 133754 700528
rect 478506 700516 478512 700528
rect 133748 700488 478512 700516
rect 133748 700476 133754 700488
rect 478506 700476 478512 700488
rect 478564 700476 478570 700528
rect 40494 700408 40500 700460
rect 40552 700448 40558 700460
rect 434438 700448 434444 700460
rect 40552 700420 434444 700448
rect 40552 700408 40558 700420
rect 434438 700408 434444 700420
rect 434496 700408 434502 700460
rect 442258 700408 442264 700460
rect 442316 700448 442322 700460
rect 559650 700448 559656 700460
rect 442316 700420 559656 700448
rect 442316 700408 442322 700420
rect 559650 700408 559656 700420
rect 559708 700408 559714 700460
rect 132586 700340 132592 700392
rect 132644 700380 132650 700392
rect 527174 700380 527180 700392
rect 132644 700352 527180 700380
rect 132644 700340 132650 700352
rect 527174 700340 527180 700352
rect 527232 700340 527238 700392
rect 132494 700272 132500 700324
rect 132552 700312 132558 700324
rect 543458 700312 543464 700324
rect 132552 700284 543464 700312
rect 132552 700272 132558 700284
rect 543458 700272 543464 700284
rect 543516 700272 543522 700324
rect 133322 700204 133328 700256
rect 133380 700244 133386 700256
rect 332502 700244 332508 700256
rect 133380 700216 332508 700244
rect 133380 700204 133386 700216
rect 332502 700204 332508 700216
rect 332560 700204 332566 700256
rect 132310 700136 132316 700188
rect 132368 700176 132374 700188
rect 283834 700176 283840 700188
rect 132368 700148 283840 700176
rect 132368 700136 132374 700148
rect 283834 700136 283840 700148
rect 283892 700136 283898 700188
rect 300118 700136 300124 700188
rect 300176 700176 300182 700188
rect 436094 700176 436100 700188
rect 300176 700148 436100 700176
rect 300176 700136 300182 700148
rect 436094 700136 436100 700148
rect 436152 700136 436158 700188
rect 132034 700068 132040 700120
rect 132092 700108 132098 700120
rect 267642 700108 267648 700120
rect 132092 700080 267648 700108
rect 132092 700068 132098 700080
rect 267642 700068 267648 700080
rect 267700 700068 267706 700120
rect 133138 700000 133144 700052
rect 133196 700040 133202 700052
rect 202782 700040 202788 700052
rect 133196 700012 202788 700040
rect 133196 700000 133202 700012
rect 202782 700000 202788 700012
rect 202840 700000 202846 700052
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 72418 699660 72424 699712
rect 72476 699700 72482 699712
rect 72970 699700 72976 699712
rect 72476 699672 72976 699700
rect 72476 699660 72482 699672
rect 72970 699660 72976 699672
rect 73028 699660 73034 699712
rect 89162 699660 89168 699712
rect 89220 699700 89226 699712
rect 89622 699700 89628 699712
rect 89220 699672 89628 699700
rect 89220 699660 89226 699672
rect 89622 699660 89628 699672
rect 89680 699660 89686 699712
rect 133046 699660 133052 699712
rect 133104 699700 133110 699712
rect 137830 699700 137836 699712
rect 133104 699672 137836 699700
rect 133104 699660 133110 699672
rect 137830 699660 137836 699672
rect 137888 699660 137894 699712
rect 429838 699660 429844 699712
rect 429896 699700 429902 699712
rect 433886 699700 433892 699712
rect 429896 699672 433892 699700
rect 429896 699660 429902 699672
rect 433886 699660 433892 699672
rect 433944 699660 433950 699712
rect 8018 698232 8024 698284
rect 8076 698272 8082 698284
rect 8202 698272 8208 698284
rect 8076 698244 8208 698272
rect 8076 698232 8082 698244
rect 8202 698232 8208 698244
rect 8260 698232 8266 698284
rect 129642 696940 129648 696992
rect 129700 696980 129706 696992
rect 580166 696980 580172 696992
rect 129700 696952 580172 696980
rect 129700 696940 129706 696952
rect 580166 696940 580172 696952
rect 580224 696940 580230 696992
rect 7926 695444 7932 695496
rect 7984 695484 7990 695496
rect 8202 695484 8208 695496
rect 7984 695456 8208 695484
rect 7984 695444 7990 695456
rect 8202 695444 8208 695456
rect 8260 695444 8266 695496
rect 7926 685856 7932 685908
rect 7984 685896 7990 685908
rect 8110 685896 8116 685908
rect 7984 685868 8116 685896
rect 7984 685856 7990 685868
rect 8110 685856 8116 685868
rect 8168 685856 8174 685908
rect 132126 685856 132132 685908
rect 132184 685896 132190 685908
rect 580166 685896 580172 685908
rect 132184 685868 580172 685896
rect 132184 685856 132190 685868
rect 580166 685856 580172 685868
rect 580224 685856 580230 685908
rect 3786 681708 3792 681760
rect 3844 681748 3850 681760
rect 434530 681748 434536 681760
rect 3844 681720 434536 681748
rect 3844 681708 3850 681720
rect 434530 681708 434536 681720
rect 434588 681708 434594 681760
rect 8110 679028 8116 679040
rect 8036 679000 8116 679028
rect 8036 678972 8064 679000
rect 8110 678988 8116 679000
rect 8168 678988 8174 679040
rect 8018 678920 8024 678972
rect 8076 678920 8082 678972
rect 8018 673480 8024 673532
rect 8076 673520 8082 673532
rect 8202 673520 8208 673532
rect 8076 673492 8208 673520
rect 8076 673480 8082 673492
rect 8202 673480 8208 673492
rect 8260 673480 8266 673532
rect 440878 673480 440884 673532
rect 440936 673520 440942 673532
rect 580166 673520 580172 673532
rect 440936 673492 580172 673520
rect 440936 673480 440942 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 8018 654100 8024 654152
rect 8076 654140 8082 654152
rect 8202 654140 8208 654152
rect 8076 654112 8208 654140
rect 8076 654100 8082 654112
rect 8202 654100 8208 654112
rect 8260 654100 8266 654152
rect 129550 650020 129556 650072
rect 129608 650060 129614 650072
rect 580166 650060 580172 650072
rect 129608 650032 580172 650060
rect 129608 650020 129614 650032
rect 580166 650020 580172 650032
rect 580224 650020 580230 650072
rect 131942 638936 131948 638988
rect 132000 638976 132006 638988
rect 580166 638976 580172 638988
rect 132000 638948 580172 638976
rect 132000 638936 132006 638948
rect 580166 638936 580172 638948
rect 580224 638936 580230 638988
rect 8018 634788 8024 634840
rect 8076 634828 8082 634840
rect 8202 634828 8208 634840
rect 8076 634800 8208 634828
rect 8076 634788 8082 634800
rect 8202 634788 8208 634800
rect 8260 634788 8266 634840
rect 439498 626560 439504 626612
rect 439556 626600 439562 626612
rect 580166 626600 580172 626612
rect 439556 626572 580172 626600
rect 439556 626560 439562 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 3050 623772 3056 623824
rect 3108 623812 3114 623824
rect 434254 623812 434260 623824
rect 3108 623784 434260 623812
rect 3108 623772 3114 623784
rect 434254 623772 434260 623784
rect 434312 623772 434318 623824
rect 8018 615476 8024 615528
rect 8076 615516 8082 615528
rect 8202 615516 8208 615528
rect 8076 615488 8208 615516
rect 8076 615476 8082 615488
rect 8202 615476 8208 615488
rect 8260 615476 8266 615528
rect 130930 603100 130936 603152
rect 130988 603140 130994 603152
rect 580166 603140 580172 603152
rect 130988 603112 580172 603140
rect 130988 603100 130994 603112
rect 580166 603100 580172 603112
rect 580224 603100 580230 603152
rect 8018 596164 8024 596216
rect 8076 596204 8082 596216
rect 8202 596204 8208 596216
rect 8076 596176 8208 596204
rect 8076 596164 8082 596176
rect 8202 596164 8208 596176
rect 8260 596164 8266 596216
rect 133966 592016 133972 592068
rect 134024 592056 134030 592068
rect 580166 592056 580172 592068
rect 134024 592028 580172 592056
rect 134024 592016 134030 592028
rect 580166 592016 580172 592028
rect 580224 592016 580230 592068
rect 126238 583652 126244 583704
rect 126296 583692 126302 583704
rect 302786 583692 302792 583704
rect 126296 583664 302792 583692
rect 126296 583652 126302 583664
rect 302786 583652 302792 583664
rect 302844 583652 302850 583704
rect 270402 583584 270408 583636
rect 270460 583624 270466 583636
rect 307018 583624 307024 583636
rect 270460 583596 307024 583624
rect 270460 583584 270466 583596
rect 307018 583584 307024 583596
rect 307076 583584 307082 583636
rect 282822 583516 282828 583568
rect 282880 583556 282886 583568
rect 313458 583556 313464 583568
rect 282880 583528 313464 583556
rect 282880 583516 282886 583528
rect 313458 583516 313464 583528
rect 313516 583516 313522 583568
rect 199378 583448 199384 583500
rect 199436 583488 199442 583500
rect 317690 583488 317696 583500
rect 199436 583460 317696 583488
rect 199436 583448 199442 583460
rect 317690 583448 317696 583460
rect 317748 583448 317754 583500
rect 128998 583380 129004 583432
rect 129056 583420 129062 583432
rect 347498 583420 347504 583432
rect 129056 583392 347504 583420
rect 129056 583380 129062 583392
rect 347498 583380 347504 583392
rect 347556 583380 347562 583432
rect 124858 583312 124864 583364
rect 124916 583352 124922 583364
rect 324130 583352 324136 583364
rect 124916 583324 324136 583352
rect 124916 583312 124922 583324
rect 324130 583312 324136 583324
rect 324188 583312 324194 583364
rect 131022 583244 131028 583296
rect 131080 583284 131086 583296
rect 349522 583284 349528 583296
rect 131080 583256 349528 583284
rect 131080 583244 131086 583256
rect 349522 583244 349528 583256
rect 349580 583244 349586 583296
rect 289722 583176 289728 583228
rect 289780 583216 289786 583228
rect 328362 583216 328368 583228
rect 289780 583188 328368 583216
rect 289780 583176 289786 583188
rect 328362 583176 328368 583188
rect 328420 583176 328426 583228
rect 275922 583108 275928 583160
rect 275980 583148 275986 583160
rect 319714 583148 319720 583160
rect 275980 583120 319720 583148
rect 275980 583108 275986 583120
rect 319714 583108 319720 583120
rect 319772 583108 319778 583160
rect 281166 583040 281172 583092
rect 281224 583080 281230 583092
rect 326154 583080 326160 583092
rect 281224 583052 326160 583080
rect 281224 583040 281230 583052
rect 326154 583040 326160 583052
rect 326212 583040 326218 583092
rect 293862 582972 293868 583024
rect 293920 583012 293926 583024
rect 338850 583012 338856 583024
rect 293920 582984 338856 583012
rect 293920 582972 293926 582984
rect 338850 582972 338856 582984
rect 338908 582972 338914 583024
rect 300394 582904 300400 582956
rect 300452 582944 300458 582956
rect 353754 582944 353760 582956
rect 300452 582916 353760 582944
rect 300452 582904 300458 582916
rect 353754 582904 353760 582916
rect 353812 582904 353818 582956
rect 300486 582836 300492 582888
rect 300544 582876 300550 582888
rect 355962 582876 355968 582888
rect 300544 582848 355968 582876
rect 300544 582836 300550 582848
rect 355962 582836 355968 582848
rect 356020 582836 356026 582888
rect 291102 582768 291108 582820
rect 291160 582808 291166 582820
rect 351730 582808 351736 582820
rect 291160 582780 351736 582808
rect 291160 582768 291166 582780
rect 351730 582768 351736 582780
rect 351788 582768 351794 582820
rect 274542 582700 274548 582752
rect 274600 582740 274606 582752
rect 368658 582740 368664 582752
rect 274600 582712 368664 582740
rect 274600 582700 274606 582712
rect 368658 582700 368664 582712
rect 368716 582700 368722 582752
rect 298922 582632 298928 582684
rect 298980 582672 298986 582684
rect 341058 582672 341064 582684
rect 298980 582644 341064 582672
rect 298980 582632 298986 582644
rect 341058 582632 341064 582644
rect 341116 582632 341122 582684
rect 357986 582632 357992 582684
rect 358044 582672 358050 582684
rect 379054 582672 379060 582684
rect 358044 582644 379060 582672
rect 358044 582632 358050 582644
rect 379054 582632 379060 582644
rect 379112 582632 379118 582684
rect 300302 582564 300308 582616
rect 300360 582604 300366 582616
rect 362402 582604 362408 582616
rect 300360 582576 362408 582604
rect 300360 582564 300366 582576
rect 362402 582564 362408 582576
rect 362460 582564 362466 582616
rect 366634 582564 366640 582616
rect 366692 582604 366698 582616
rect 377582 582604 377588 582616
rect 366692 582576 377588 582604
rect 366692 582564 366698 582576
rect 377582 582564 377588 582576
rect 377640 582564 377646 582616
rect 299290 582496 299296 582548
rect 299348 582536 299354 582548
rect 332594 582536 332600 582548
rect 299348 582508 332600 582536
rect 299348 582496 299354 582508
rect 332594 582496 332600 582508
rect 332652 582496 332658 582548
rect 370866 582496 370872 582548
rect 370924 582536 370930 582548
rect 377306 582536 377312 582548
rect 370924 582508 377312 582536
rect 370924 582496 370930 582508
rect 377306 582496 377312 582508
rect 377364 582496 377370 582548
rect 298738 582428 298744 582480
rect 298796 582468 298802 582480
rect 321922 582468 321928 582480
rect 298796 582440 321928 582468
rect 298796 582428 298802 582440
rect 321922 582428 321928 582440
rect 321980 582428 321986 582480
rect 372890 582428 372896 582480
rect 372948 582468 372954 582480
rect 377490 582468 377496 582480
rect 372948 582440 377496 582468
rect 372948 582428 372954 582440
rect 377490 582428 377496 582440
rect 377548 582428 377554 582480
rect 298830 582360 298836 582412
rect 298888 582400 298894 582412
rect 309226 582400 309232 582412
rect 298888 582372 309232 582400
rect 298888 582360 298894 582372
rect 309226 582360 309232 582372
rect 309284 582360 309290 582412
rect 299198 579640 299204 579692
rect 299256 579680 299262 579692
rect 304810 579680 304816 579692
rect 299256 579652 304816 579680
rect 299256 579640 299262 579652
rect 304810 579640 304816 579652
rect 304868 579640 304874 579692
rect 438210 579640 438216 579692
rect 438268 579680 438274 579692
rect 580166 579680 580172 579692
rect 438268 579652 580172 579680
rect 438268 579640 438274 579652
rect 580166 579640 580172 579652
rect 580224 579640 580230 579692
rect 7650 579572 7656 579624
rect 7708 579612 7714 579624
rect 7926 579612 7932 579624
rect 7708 579584 7932 579612
rect 7708 579572 7714 579584
rect 7926 579572 7932 579584
rect 7984 579572 7990 579624
rect 305086 579572 305092 579624
rect 305144 579612 305150 579624
rect 315206 579612 315212 579624
rect 305144 579584 315212 579612
rect 305144 579572 305150 579584
rect 315206 579572 315212 579584
rect 315264 579572 315270 579624
rect 330754 579572 330760 579624
rect 330812 579612 330818 579624
rect 334802 579612 334808 579624
rect 330812 579584 334808 579612
rect 330812 579572 330818 579584
rect 334802 579572 334808 579584
rect 334860 579572 334866 579624
rect 330662 579504 330668 579556
rect 330720 579544 330726 579556
rect 335170 579544 335176 579556
rect 330720 579516 335176 579544
rect 330720 579504 330726 579516
rect 335170 579504 335176 579516
rect 335228 579504 335234 579556
rect 300210 579436 300216 579488
rect 300268 579476 300274 579488
rect 310974 579476 310980 579488
rect 300268 579448 310980 579476
rect 300268 579436 300274 579448
rect 310974 579436 310980 579448
rect 311032 579436 311038 579488
rect 330570 579436 330576 579488
rect 330628 579476 330634 579488
rect 338666 579476 338672 579488
rect 330628 579448 338672 579476
rect 330628 579436 330634 579448
rect 338666 579436 338672 579448
rect 338724 579436 338730 579488
rect 336550 579408 336556 579420
rect 306944 579380 309916 579408
rect 299474 579300 299480 579352
rect 299532 579340 299538 579352
rect 300670 579340 300676 579352
rect 299532 579312 300676 579340
rect 299532 579300 299538 579312
rect 300670 579300 300676 579312
rect 300728 579300 300734 579352
rect 305086 579340 305092 579352
rect 305012 579312 305092 579340
rect 299566 579164 299572 579216
rect 299624 579204 299630 579216
rect 305012 579204 305040 579312
rect 305086 579300 305092 579312
rect 305144 579300 305150 579352
rect 305178 579300 305184 579352
rect 305236 579300 305242 579352
rect 305196 579272 305224 579300
rect 299624 579176 305040 579204
rect 305104 579244 305224 579272
rect 299624 579164 299630 579176
rect 157334 579028 157340 579080
rect 157392 579068 157398 579080
rect 162394 579068 162400 579080
rect 157392 579040 162400 579068
rect 157392 579028 157398 579040
rect 162394 579028 162400 579040
rect 162452 579028 162458 579080
rect 176654 579028 176660 579080
rect 176712 579068 176718 579080
rect 181714 579068 181720 579080
rect 176712 579040 181720 579068
rect 176712 579028 176718 579040
rect 181714 579028 181720 579040
rect 181772 579028 181778 579080
rect 195974 579028 195980 579080
rect 196032 579068 196038 579080
rect 201034 579068 201040 579080
rect 196032 579040 201040 579068
rect 196032 579028 196038 579040
rect 201034 579028 201040 579040
rect 201092 579028 201098 579080
rect 215294 579028 215300 579080
rect 215352 579068 215358 579080
rect 220354 579068 220360 579080
rect 215352 579040 220360 579068
rect 215352 579028 215358 579040
rect 220354 579028 220360 579040
rect 220412 579028 220418 579080
rect 234614 579028 234620 579080
rect 234672 579068 234678 579080
rect 239674 579068 239680 579080
rect 234672 579040 239680 579068
rect 234672 579028 234678 579040
rect 239674 579028 239680 579040
rect 239732 579028 239738 579080
rect 253934 579028 253940 579080
rect 253992 579068 253998 579080
rect 258994 579068 259000 579080
rect 253992 579040 259000 579068
rect 253992 579028 253998 579040
rect 258994 579028 259000 579040
rect 259052 579028 259058 579080
rect 300210 579068 300216 579080
rect 297100 579040 300216 579068
rect 130378 578960 130384 579012
rect 130436 579000 130442 579012
rect 152550 579000 152556 579012
rect 130436 578972 152556 579000
rect 130436 578960 130442 578972
rect 152550 578960 152556 578972
rect 152608 578960 152614 579012
rect 171870 579000 171876 579012
rect 162136 578972 171876 579000
rect 125686 578892 125692 578944
rect 125744 578932 125750 578944
rect 137830 578932 137836 578944
rect 125744 578904 137836 578932
rect 125744 578892 125750 578904
rect 137830 578892 137836 578904
rect 137888 578892 137894 578944
rect 147582 578892 147588 578944
rect 147640 578932 147646 578944
rect 152274 578932 152280 578944
rect 147640 578904 152280 578932
rect 147640 578892 147646 578904
rect 152274 578892 152280 578904
rect 152332 578892 152338 578944
rect 152366 578892 152372 578944
rect 152424 578932 152430 578944
rect 157242 578932 157248 578944
rect 152424 578904 157248 578932
rect 152424 578892 152430 578904
rect 157242 578892 157248 578904
rect 157300 578892 157306 578944
rect 138658 578756 138664 578808
rect 138716 578796 138722 578808
rect 152458 578796 152464 578808
rect 138716 578768 152464 578796
rect 138716 578756 138722 578768
rect 152458 578756 152464 578768
rect 152516 578756 152522 578808
rect 152550 578756 152556 578808
rect 152608 578796 152614 578808
rect 152608 578768 157288 578796
rect 152608 578756 152614 578768
rect 122742 578688 122748 578740
rect 122800 578728 122806 578740
rect 147582 578728 147588 578740
rect 122800 578700 128400 578728
rect 122800 578688 122806 578700
rect 128372 578660 128400 578700
rect 138032 578700 147588 578728
rect 138032 578660 138060 578700
rect 147582 578688 147588 578700
rect 147640 578688 147646 578740
rect 157260 578728 157288 578768
rect 162136 578728 162164 578972
rect 171870 578960 171876 578972
rect 171928 578960 171934 579012
rect 191190 579000 191196 579012
rect 181456 578972 191196 579000
rect 171594 578932 171600 578944
rect 157260 578700 162164 578728
rect 162228 578904 171600 578932
rect 128372 578632 138060 578660
rect 138106 578620 138112 578672
rect 138164 578660 138170 578672
rect 139578 578660 139584 578672
rect 138164 578632 139584 578660
rect 138164 578620 138170 578632
rect 139578 578620 139584 578632
rect 139636 578620 139642 578672
rect 152274 578620 152280 578672
rect 152332 578660 152338 578672
rect 162228 578660 162256 578904
rect 171594 578892 171600 578904
rect 171652 578892 171658 578944
rect 171686 578892 171692 578944
rect 171744 578932 171750 578944
rect 176562 578932 176568 578944
rect 171744 578904 176568 578932
rect 171744 578892 171750 578904
rect 176562 578892 176568 578904
rect 176620 578892 176626 578944
rect 162302 578756 162308 578808
rect 162360 578796 162366 578808
rect 171778 578796 171784 578808
rect 162360 578768 171784 578796
rect 162360 578756 162366 578768
rect 171778 578756 171784 578768
rect 171836 578756 171842 578808
rect 171870 578756 171876 578808
rect 171928 578796 171934 578808
rect 171928 578768 176608 578796
rect 171928 578756 171934 578768
rect 176580 578728 176608 578768
rect 181456 578728 181484 578972
rect 191190 578960 191196 578972
rect 191248 578960 191254 579012
rect 210510 579000 210516 579012
rect 200776 578972 210516 579000
rect 190914 578932 190920 578944
rect 176580 578700 181484 578728
rect 181548 578904 190920 578932
rect 152332 578632 162256 578660
rect 152332 578620 152338 578632
rect 171594 578620 171600 578672
rect 171652 578660 171658 578672
rect 181548 578660 181576 578904
rect 190914 578892 190920 578904
rect 190972 578892 190978 578944
rect 191006 578892 191012 578944
rect 191064 578932 191070 578944
rect 195882 578932 195888 578944
rect 191064 578904 195888 578932
rect 191064 578892 191070 578904
rect 195882 578892 195888 578904
rect 195940 578892 195946 578944
rect 181622 578756 181628 578808
rect 181680 578796 181686 578808
rect 191098 578796 191104 578808
rect 181680 578768 191104 578796
rect 181680 578756 181686 578768
rect 191098 578756 191104 578768
rect 191156 578756 191162 578808
rect 191190 578756 191196 578808
rect 191248 578796 191254 578808
rect 191248 578768 195928 578796
rect 191248 578756 191254 578768
rect 195900 578728 195928 578768
rect 200776 578728 200804 578972
rect 210510 578960 210516 578972
rect 210568 578960 210574 579012
rect 229830 579000 229836 579012
rect 220096 578972 229836 579000
rect 210234 578932 210240 578944
rect 195900 578700 200804 578728
rect 200868 578904 210240 578932
rect 171652 578632 181576 578660
rect 171652 578620 171658 578632
rect 190914 578620 190920 578672
rect 190972 578660 190978 578672
rect 200868 578660 200896 578904
rect 210234 578892 210240 578904
rect 210292 578892 210298 578944
rect 210326 578892 210332 578944
rect 210384 578932 210390 578944
rect 215202 578932 215208 578944
rect 210384 578904 215208 578932
rect 210384 578892 210390 578904
rect 215202 578892 215208 578904
rect 215260 578892 215266 578944
rect 200942 578756 200948 578808
rect 201000 578796 201006 578808
rect 210418 578796 210424 578808
rect 201000 578768 210424 578796
rect 201000 578756 201006 578768
rect 210418 578756 210424 578768
rect 210476 578756 210482 578808
rect 210510 578756 210516 578808
rect 210568 578796 210574 578808
rect 210568 578768 215248 578796
rect 210568 578756 210574 578768
rect 215220 578728 215248 578768
rect 220096 578728 220124 578972
rect 229830 578960 229836 578972
rect 229888 578960 229894 579012
rect 249150 579000 249156 579012
rect 239416 578972 249156 579000
rect 229554 578932 229560 578944
rect 215220 578700 220124 578728
rect 220188 578904 229560 578932
rect 190972 578632 200896 578660
rect 190972 578620 190978 578632
rect 210234 578620 210240 578672
rect 210292 578660 210298 578672
rect 220188 578660 220216 578904
rect 229554 578892 229560 578904
rect 229612 578892 229618 578944
rect 229646 578892 229652 578944
rect 229704 578932 229710 578944
rect 234522 578932 234528 578944
rect 229704 578904 234528 578932
rect 229704 578892 229710 578904
rect 234522 578892 234528 578904
rect 234580 578892 234586 578944
rect 220262 578756 220268 578808
rect 220320 578796 220326 578808
rect 229738 578796 229744 578808
rect 220320 578768 229744 578796
rect 220320 578756 220326 578768
rect 229738 578756 229744 578768
rect 229796 578756 229802 578808
rect 229830 578756 229836 578808
rect 229888 578796 229894 578808
rect 229888 578768 234568 578796
rect 229888 578756 229894 578768
rect 234540 578728 234568 578768
rect 239416 578728 239444 578972
rect 249150 578960 249156 578972
rect 249208 578960 249214 579012
rect 268470 579000 268476 579012
rect 258736 578972 268476 579000
rect 248874 578932 248880 578944
rect 234540 578700 239444 578728
rect 239508 578904 248880 578932
rect 210292 578632 220216 578660
rect 210292 578620 210298 578632
rect 229554 578620 229560 578672
rect 229612 578660 229618 578672
rect 239508 578660 239536 578904
rect 248874 578892 248880 578904
rect 248932 578892 248938 578944
rect 248966 578892 248972 578944
rect 249024 578932 249030 578944
rect 253842 578932 253848 578944
rect 249024 578904 253848 578932
rect 249024 578892 249030 578904
rect 253842 578892 253848 578904
rect 253900 578892 253906 578944
rect 239582 578756 239588 578808
rect 239640 578796 239646 578808
rect 249058 578796 249064 578808
rect 239640 578768 249064 578796
rect 239640 578756 239646 578768
rect 249058 578756 249064 578768
rect 249116 578756 249122 578808
rect 249150 578756 249156 578808
rect 249208 578796 249214 578808
rect 249208 578768 253888 578796
rect 249208 578756 249214 578768
rect 253860 578728 253888 578768
rect 258736 578728 258764 578972
rect 268470 578960 268476 578972
rect 268528 578960 268534 579012
rect 282914 578960 282920 579012
rect 282972 579000 282978 579012
rect 297100 579000 297128 579040
rect 300210 579028 300216 579040
rect 300268 579028 300274 579080
rect 282972 578972 297128 579000
rect 282972 578960 282978 578972
rect 297174 578960 297180 579012
rect 297232 579000 297238 579012
rect 299566 579000 299572 579012
rect 297232 578972 299572 579000
rect 297232 578960 297238 578972
rect 299566 578960 299572 578972
rect 299624 578960 299630 579012
rect 268102 578932 268108 578944
rect 253860 578700 258764 578728
rect 258828 578904 268108 578932
rect 229612 578632 239536 578660
rect 229612 578620 229618 578632
rect 248874 578620 248880 578672
rect 248932 578660 248938 578672
rect 258828 578660 258856 578904
rect 268102 578892 268108 578904
rect 268160 578892 268166 578944
rect 268286 578892 268292 578944
rect 268344 578932 268350 578944
rect 273162 578932 273168 578944
rect 268344 578904 273168 578932
rect 268344 578892 268350 578904
rect 273162 578892 273168 578904
rect 273220 578892 273226 578944
rect 277946 578892 277952 578944
rect 278004 578932 278010 578944
rect 294598 578932 294604 578944
rect 278004 578904 294604 578932
rect 278004 578892 278010 578904
rect 294598 578892 294604 578904
rect 294656 578892 294662 578944
rect 300210 578892 300216 578944
rect 300268 578932 300274 578944
rect 305104 578932 305132 579244
rect 300268 578904 305132 578932
rect 300268 578892 300274 578904
rect 278038 578824 278044 578876
rect 278096 578864 278102 578876
rect 278096 578836 287560 578864
rect 278096 578824 278102 578836
rect 258902 578756 258908 578808
rect 258960 578796 258966 578808
rect 268378 578796 268384 578808
rect 258960 578768 268384 578796
rect 258960 578756 258966 578768
rect 268378 578756 268384 578768
rect 268436 578756 268442 578808
rect 268470 578756 268476 578808
rect 268528 578796 268534 578808
rect 282914 578796 282920 578808
rect 268528 578768 273208 578796
rect 268528 578756 268534 578768
rect 273180 578728 273208 578768
rect 273272 578768 282920 578796
rect 273272 578728 273300 578768
rect 282914 578756 282920 578768
rect 282972 578756 282978 578808
rect 273180 578700 273300 578728
rect 248932 578632 258856 578660
rect 248932 578620 248938 578632
rect 268102 578620 268108 578672
rect 268160 578660 268166 578672
rect 278038 578660 278044 578672
rect 268160 578632 278044 578660
rect 268160 578620 268166 578632
rect 278038 578620 278044 578632
rect 278096 578620 278102 578672
rect 287532 578660 287560 578836
rect 287698 578824 287704 578876
rect 287756 578864 287762 578876
rect 289814 578864 289820 578876
rect 287756 578836 289820 578864
rect 287756 578824 287762 578836
rect 289814 578824 289820 578836
rect 289872 578824 289878 578876
rect 298002 578824 298008 578876
rect 298060 578864 298066 578876
rect 298060 578836 304304 578864
rect 298060 578824 298066 578836
rect 299382 578756 299388 578808
rect 299440 578796 299446 578808
rect 300210 578796 300216 578808
rect 299440 578768 300216 578796
rect 299440 578756 299446 578768
rect 300210 578756 300216 578768
rect 300268 578756 300274 578808
rect 304276 578796 304304 578836
rect 306944 578796 306972 579380
rect 309778 579300 309784 579352
rect 309836 579300 309842 579352
rect 304276 578768 306972 578796
rect 297082 578688 297088 578740
rect 297140 578728 297146 578740
rect 300118 578728 300124 578740
rect 297140 578700 300124 578728
rect 297140 578688 297146 578700
rect 300118 578688 300124 578700
rect 300176 578688 300182 578740
rect 309796 578728 309824 579300
rect 309888 579136 309916 579380
rect 330220 579380 336556 579408
rect 309962 579300 309968 579352
rect 310020 579340 310026 579352
rect 310020 579312 310100 579340
rect 310020 579300 310026 579312
rect 309888 579108 310008 579136
rect 309980 579000 310008 579108
rect 310072 579068 310100 579312
rect 315850 579300 315856 579352
rect 315908 579300 315914 579352
rect 330018 579300 330024 579352
rect 330076 579300 330082 579352
rect 315868 579272 315896 579300
rect 330036 579272 330064 579300
rect 315868 579244 330064 579272
rect 330220 579136 330248 579380
rect 336550 579368 336556 579380
rect 336608 579368 336614 579420
rect 342990 579408 342996 579420
rect 338592 579380 342996 579408
rect 330570 579300 330576 579352
rect 330628 579300 330634 579352
rect 330662 579300 330668 579352
rect 330720 579300 330726 579352
rect 330754 579300 330760 579352
rect 330812 579300 330818 579352
rect 334434 579300 334440 579352
rect 334492 579300 334498 579352
rect 334710 579300 334716 579352
rect 334768 579300 334774 579352
rect 334802 579300 334808 579352
rect 334860 579300 334866 579352
rect 334894 579300 334900 579352
rect 334952 579300 334958 579352
rect 335170 579300 335176 579352
rect 335228 579300 335234 579352
rect 329024 579108 330248 579136
rect 329024 579068 329052 579108
rect 310072 579040 329052 579068
rect 309888 578972 310008 579000
rect 309888 578864 309916 578972
rect 322216 578904 327028 578932
rect 322216 578864 322244 578904
rect 309888 578836 317460 578864
rect 317432 578796 317460 578836
rect 321940 578836 322244 578864
rect 327000 578864 327028 578904
rect 330588 578864 330616 579300
rect 327000 578836 330616 578864
rect 321940 578796 321968 578836
rect 330680 578796 330708 579300
rect 317432 578768 321968 578796
rect 322216 578768 330708 578796
rect 304184 578700 309824 578728
rect 297174 578660 297180 578672
rect 287532 578632 297180 578660
rect 297174 578620 297180 578632
rect 297232 578620 297238 578672
rect 115198 578552 115204 578604
rect 115256 578592 115262 578604
rect 115934 578592 115940 578604
rect 115256 578564 115940 578592
rect 115256 578552 115262 578564
rect 115934 578552 115940 578564
rect 115992 578552 115998 578604
rect 129090 578552 129096 578604
rect 129148 578592 129154 578604
rect 287698 578592 287704 578604
rect 129148 578564 287704 578592
rect 129148 578552 129154 578564
rect 287698 578552 287704 578564
rect 287756 578552 287762 578604
rect 294506 578552 294512 578604
rect 294564 578592 294570 578604
rect 304184 578592 304212 578700
rect 322216 578660 322244 578768
rect 330772 578728 330800 579300
rect 294564 578564 304212 578592
rect 309520 578632 322244 578660
rect 322308 578700 330800 578728
rect 294564 578552 294570 578564
rect 119338 578484 119344 578536
rect 119396 578524 119402 578536
rect 125686 578524 125692 578536
rect 119396 578496 125692 578524
rect 119396 578484 119402 578496
rect 125686 578484 125692 578496
rect 125744 578484 125750 578536
rect 137922 578484 137928 578536
rect 137980 578524 137986 578536
rect 138014 578524 138020 578536
rect 137980 578496 138020 578524
rect 137980 578484 137986 578496
rect 138014 578484 138020 578496
rect 138072 578484 138078 578536
rect 157242 578484 157248 578536
rect 157300 578524 157306 578536
rect 157334 578524 157340 578536
rect 157300 578496 157340 578524
rect 157300 578484 157306 578496
rect 157334 578484 157340 578496
rect 157392 578484 157398 578536
rect 176562 578484 176568 578536
rect 176620 578524 176626 578536
rect 176654 578524 176660 578536
rect 176620 578496 176660 578524
rect 176620 578484 176626 578496
rect 176654 578484 176660 578496
rect 176712 578484 176718 578536
rect 195882 578484 195888 578536
rect 195940 578524 195946 578536
rect 195974 578524 195980 578536
rect 195940 578496 195980 578524
rect 195940 578484 195946 578496
rect 195974 578484 195980 578496
rect 196032 578484 196038 578536
rect 215202 578484 215208 578536
rect 215260 578524 215266 578536
rect 215294 578524 215300 578536
rect 215260 578496 215300 578524
rect 215260 578484 215266 578496
rect 215294 578484 215300 578496
rect 215352 578484 215358 578536
rect 234522 578484 234528 578536
rect 234580 578524 234586 578536
rect 234614 578524 234620 578536
rect 234580 578496 234620 578524
rect 234580 578484 234586 578496
rect 234614 578484 234620 578496
rect 234672 578484 234678 578536
rect 253842 578484 253848 578536
rect 253900 578524 253906 578536
rect 253934 578524 253940 578536
rect 253900 578496 253940 578524
rect 253900 578484 253906 578496
rect 253934 578484 253940 578496
rect 253992 578484 253998 578536
rect 273162 578484 273168 578536
rect 273220 578524 273226 578536
rect 273220 578496 282868 578524
rect 273220 578484 273226 578496
rect 138658 578456 138664 578468
rect 128188 578428 138664 578456
rect 125502 578348 125508 578400
rect 125560 578388 125566 578400
rect 128188 578388 128216 578428
rect 138658 578416 138664 578428
rect 138716 578416 138722 578468
rect 139578 578416 139584 578468
rect 139636 578456 139642 578468
rect 152366 578456 152372 578468
rect 139636 578428 152372 578456
rect 139636 578416 139642 578428
rect 152366 578416 152372 578428
rect 152424 578416 152430 578468
rect 152458 578416 152464 578468
rect 152516 578456 152522 578468
rect 162302 578456 162308 578468
rect 152516 578428 162308 578456
rect 152516 578416 152522 578428
rect 162302 578416 162308 578428
rect 162360 578416 162366 578468
rect 162394 578416 162400 578468
rect 162452 578456 162458 578468
rect 171686 578456 171692 578468
rect 162452 578428 171692 578456
rect 162452 578416 162458 578428
rect 171686 578416 171692 578428
rect 171744 578416 171750 578468
rect 171778 578416 171784 578468
rect 171836 578456 171842 578468
rect 181622 578456 181628 578468
rect 171836 578428 181628 578456
rect 171836 578416 171842 578428
rect 181622 578416 181628 578428
rect 181680 578416 181686 578468
rect 181714 578416 181720 578468
rect 181772 578456 181778 578468
rect 191006 578456 191012 578468
rect 181772 578428 191012 578456
rect 181772 578416 181778 578428
rect 191006 578416 191012 578428
rect 191064 578416 191070 578468
rect 191098 578416 191104 578468
rect 191156 578456 191162 578468
rect 200942 578456 200948 578468
rect 191156 578428 200948 578456
rect 191156 578416 191162 578428
rect 200942 578416 200948 578428
rect 201000 578416 201006 578468
rect 201034 578416 201040 578468
rect 201092 578456 201098 578468
rect 210326 578456 210332 578468
rect 201092 578428 210332 578456
rect 201092 578416 201098 578428
rect 210326 578416 210332 578428
rect 210384 578416 210390 578468
rect 210418 578416 210424 578468
rect 210476 578456 210482 578468
rect 220262 578456 220268 578468
rect 210476 578428 220268 578456
rect 210476 578416 210482 578428
rect 220262 578416 220268 578428
rect 220320 578416 220326 578468
rect 220354 578416 220360 578468
rect 220412 578456 220418 578468
rect 229646 578456 229652 578468
rect 220412 578428 229652 578456
rect 220412 578416 220418 578428
rect 229646 578416 229652 578428
rect 229704 578416 229710 578468
rect 229738 578416 229744 578468
rect 229796 578456 229802 578468
rect 239582 578456 239588 578468
rect 229796 578428 239588 578456
rect 229796 578416 229802 578428
rect 239582 578416 239588 578428
rect 239640 578416 239646 578468
rect 239674 578416 239680 578468
rect 239732 578456 239738 578468
rect 248966 578456 248972 578468
rect 239732 578428 248972 578456
rect 239732 578416 239738 578428
rect 248966 578416 248972 578428
rect 249024 578416 249030 578468
rect 249058 578416 249064 578468
rect 249116 578456 249122 578468
rect 258902 578456 258908 578468
rect 249116 578428 258908 578456
rect 249116 578416 249122 578428
rect 258902 578416 258908 578428
rect 258960 578416 258966 578468
rect 258994 578416 259000 578468
rect 259052 578456 259058 578468
rect 268286 578456 268292 578468
rect 259052 578428 268292 578456
rect 259052 578416 259058 578428
rect 268286 578416 268292 578428
rect 268344 578416 268350 578468
rect 268378 578416 268384 578468
rect 268436 578456 268442 578468
rect 277946 578456 277952 578468
rect 268436 578428 277952 578456
rect 268436 578416 268442 578428
rect 277946 578416 277952 578428
rect 278004 578416 278010 578468
rect 282840 578456 282868 578496
rect 300118 578484 300124 578536
rect 300176 578524 300182 578536
rect 309520 578524 309548 578632
rect 300176 578496 309548 578524
rect 300176 578484 300182 578496
rect 294506 578456 294512 578468
rect 282840 578428 294512 578456
rect 294506 578416 294512 578428
rect 294564 578416 294570 578468
rect 294598 578416 294604 578468
rect 294656 578456 294662 578468
rect 297082 578456 297088 578468
rect 294656 578428 297088 578456
rect 294656 578416 294662 578428
rect 297082 578416 297088 578428
rect 297140 578416 297146 578468
rect 313568 578428 314424 578456
rect 125560 578360 128216 578388
rect 125560 578348 125566 578360
rect 129274 578348 129280 578400
rect 129332 578388 129338 578400
rect 313568 578388 313596 578428
rect 129332 578360 313596 578388
rect 129332 578348 129338 578360
rect 85390 578280 85396 578332
rect 85448 578320 85454 578332
rect 125594 578320 125600 578332
rect 85448 578292 125600 578320
rect 85448 578280 85454 578292
rect 125594 578280 125600 578292
rect 125652 578280 125658 578332
rect 125778 578280 125784 578332
rect 125836 578320 125842 578332
rect 125836 578292 313688 578320
rect 125836 578280 125842 578292
rect 85574 578212 85580 578264
rect 85632 578252 85638 578264
rect 85632 578224 313320 578252
rect 85632 578212 85638 578224
rect 313292 577980 313320 578224
rect 313660 578184 313688 578292
rect 314396 578252 314424 578428
rect 322308 578252 322336 578700
rect 334452 578388 334480 579300
rect 314396 578224 322336 578252
rect 325528 578360 334480 578388
rect 325528 578184 325556 578360
rect 334728 578320 334756 579300
rect 313660 578156 325556 578184
rect 325712 578292 334756 578320
rect 325712 578116 325740 578292
rect 334820 578184 334848 579300
rect 334912 578320 334940 579300
rect 335188 578456 335216 579300
rect 338592 578660 338620 579380
rect 342990 579368 342996 579380
rect 343048 579368 343054 579420
rect 343192 579380 345520 579408
rect 338666 579300 338672 579352
rect 338724 579300 338730 579352
rect 338684 579272 338712 579300
rect 338684 579244 339080 579272
rect 339052 579000 339080 579244
rect 343192 579000 343220 579380
rect 345106 579300 345112 579352
rect 345164 579300 345170 579352
rect 339052 578972 343220 579000
rect 335464 578632 338620 578660
rect 338684 578632 338988 578660
rect 335464 578456 335492 578632
rect 335188 578428 335492 578456
rect 334912 578292 335308 578320
rect 335280 578184 335308 578292
rect 338684 578184 338712 578632
rect 338960 578592 338988 578632
rect 338960 578564 339356 578592
rect 339328 578524 339356 578564
rect 345124 578524 345152 579300
rect 345492 578728 345520 579380
rect 360378 579300 360384 579352
rect 360436 579300 360442 579352
rect 364242 579300 364248 579352
rect 364300 579300 364306 579352
rect 375374 579300 375380 579352
rect 375432 579340 375438 579352
rect 378962 579340 378968 579352
rect 375432 579312 378968 579340
rect 375432 579300 375438 579312
rect 378962 579300 378968 579312
rect 379020 579300 379026 579352
rect 360396 578932 360424 579300
rect 360212 578904 360424 578932
rect 360212 578864 360240 578904
rect 360120 578836 360240 578864
rect 360120 578796 360148 578836
rect 350552 578768 360148 578796
rect 350552 578728 350580 578768
rect 345492 578700 350580 578728
rect 339328 578496 345152 578524
rect 364260 578388 364288 579300
rect 339236 578360 364288 578388
rect 339236 578252 339264 578360
rect 334820 578156 334940 578184
rect 335280 578156 338712 578184
rect 338776 578224 339264 578252
rect 316696 578088 325740 578116
rect 316696 577980 316724 578088
rect 334912 578048 334940 578156
rect 338776 578116 338804 578224
rect 335188 578088 338804 578116
rect 335188 578048 335216 578088
rect 334912 578020 335216 578048
rect 313292 577952 316724 577980
rect 110322 575492 110328 575544
rect 110380 575532 110386 575544
rect 296714 575532 296720 575544
rect 110380 575504 296720 575532
rect 110380 575492 110386 575504
rect 296714 575492 296720 575504
rect 296772 575492 296778 575544
rect 281258 572704 281264 572756
rect 281316 572704 281322 572756
rect 281276 572620 281304 572704
rect 281258 572568 281264 572620
rect 281316 572568 281322 572620
rect 7650 569916 7656 569968
rect 7708 569956 7714 569968
rect 7834 569956 7840 569968
rect 7708 569928 7840 569956
rect 7708 569916 7714 569928
rect 7834 569916 7840 569928
rect 7892 569916 7898 569968
rect 271782 569916 271788 569968
rect 271840 569956 271846 569968
rect 296714 569956 296720 569968
rect 271840 569928 296720 569956
rect 271840 569916 271846 569928
rect 296714 569916 296720 569928
rect 296772 569916 296778 569968
rect 281074 569780 281080 569832
rect 281132 569820 281138 569832
rect 281258 569820 281264 569832
rect 281132 569792 281264 569820
rect 281132 569780 281138 569792
rect 281258 569780 281264 569792
rect 281316 569780 281322 569832
rect 7834 563048 7840 563100
rect 7892 563048 7898 563100
rect 129458 563048 129464 563100
rect 129516 563088 129522 563100
rect 296714 563088 296720 563100
rect 129516 563060 296720 563088
rect 129516 563048 129522 563060
rect 296714 563048 296720 563060
rect 296772 563048 296778 563100
rect 7852 562952 7880 563048
rect 7926 562952 7932 562964
rect 7852 562924 7932 562952
rect 7926 562912 7932 562924
rect 7984 562912 7990 562964
rect 200114 562096 200120 562148
rect 200172 562136 200178 562148
rect 209682 562136 209688 562148
rect 200172 562108 209688 562136
rect 200172 562096 200178 562108
rect 209682 562096 209688 562108
rect 209740 562096 209746 562148
rect 195790 562028 195796 562080
rect 195848 562068 195854 562080
rect 214742 562068 214748 562080
rect 195848 562040 214748 562068
rect 195848 562028 195854 562040
rect 214742 562028 214748 562040
rect 214800 562028 214806 562080
rect 195698 561960 195704 562012
rect 195756 562000 195762 562012
rect 205542 562000 205548 562012
rect 195756 561972 205548 562000
rect 195756 561960 195762 561972
rect 205542 561960 205548 561972
rect 205600 561960 205606 562012
rect 197262 561892 197268 561944
rect 197320 561932 197326 561944
rect 208670 561932 208676 561944
rect 197320 561904 208676 561932
rect 197320 561892 197326 561904
rect 208670 561892 208676 561904
rect 208728 561892 208734 561944
rect 195882 561824 195888 561876
rect 195940 561864 195946 561876
rect 211614 561864 211620 561876
rect 195940 561836 211620 561864
rect 195940 561824 195946 561836
rect 211614 561824 211620 561836
rect 211672 561824 211678 561876
rect 197170 561756 197176 561808
rect 197228 561796 197234 561808
rect 200114 561796 200120 561808
rect 197228 561768 200120 561796
rect 197228 561756 197234 561768
rect 200114 561756 200120 561768
rect 200172 561756 200178 561808
rect 209682 561688 209688 561740
rect 209740 561728 209746 561740
rect 217870 561728 217876 561740
rect 209740 561700 217876 561728
rect 209740 561688 209746 561700
rect 217870 561688 217876 561700
rect 217928 561688 217934 561740
rect 281074 560260 281080 560312
rect 281132 560300 281138 560312
rect 281258 560300 281264 560312
rect 281132 560272 281264 560300
rect 281132 560260 281138 560272
rect 281258 560260 281264 560272
rect 281316 560260 281322 560312
rect 197078 560192 197084 560244
rect 197136 560232 197142 560244
rect 202046 560232 202052 560244
rect 197136 560204 202052 560232
rect 197136 560192 197142 560204
rect 202046 560192 202052 560204
rect 202104 560192 202110 560244
rect 418798 556248 418804 556300
rect 418856 556288 418862 556300
rect 511258 556288 511264 556300
rect 418856 556260 511264 556288
rect 418856 556248 418862 556260
rect 511258 556248 511264 556260
rect 511316 556248 511322 556300
rect 273162 556180 273168 556232
rect 273220 556220 273226 556232
rect 297818 556220 297824 556232
rect 273220 556192 297824 556220
rect 273220 556180 273226 556192
rect 297818 556180 297824 556192
rect 297876 556180 297882 556232
rect 378778 556180 378784 556232
rect 378836 556220 378842 556232
rect 484394 556220 484400 556232
rect 378836 556192 484400 556220
rect 378836 556180 378842 556192
rect 484394 556180 484400 556192
rect 484452 556180 484458 556232
rect 109402 554752 109408 554804
rect 109460 554792 109466 554804
rect 110322 554792 110328 554804
rect 109460 554764 110328 554792
rect 109460 554752 109466 554764
rect 110322 554752 110328 554764
rect 110380 554792 110386 554804
rect 115934 554792 115940 554804
rect 110380 554764 115940 554792
rect 110380 554752 110386 554764
rect 115934 554752 115940 554764
rect 115992 554752 115998 554804
rect 92106 553936 92112 553988
rect 92164 553976 92170 553988
rect 115290 553976 115296 553988
rect 92164 553948 115296 553976
rect 92164 553936 92170 553948
rect 115290 553936 115296 553948
rect 115348 553936 115354 553988
rect 89162 553868 89168 553920
rect 89220 553908 89226 553920
rect 156598 553908 156604 553920
rect 89220 553880 156604 553908
rect 89220 553868 89226 553880
rect 156598 553868 156604 553880
rect 156656 553868 156662 553920
rect 115106 553800 115112 553852
rect 115164 553840 115170 553852
rect 128446 553840 128452 553852
rect 115164 553812 128452 553840
rect 115164 553800 115170 553812
rect 128446 553800 128452 553812
rect 128504 553840 128510 553852
rect 128998 553840 129004 553852
rect 128504 553812 129004 553840
rect 128504 553800 128510 553812
rect 128998 553800 129004 553812
rect 129056 553800 129062 553852
rect 95050 553732 95056 553784
rect 95108 553772 95114 553784
rect 120718 553772 120724 553784
rect 95108 553744 120724 553772
rect 95108 553732 95114 553744
rect 120718 553732 120724 553744
rect 120776 553732 120782 553784
rect 100754 553664 100760 553716
rect 100812 553704 100818 553716
rect 129182 553704 129188 553716
rect 100812 553676 129188 553704
rect 100812 553664 100818 553676
rect 129182 553664 129188 553676
rect 129240 553664 129246 553716
rect 106458 553596 106464 553648
rect 106516 553636 106522 553648
rect 137278 553636 137284 553648
rect 106516 553608 137284 553636
rect 106516 553596 106522 553608
rect 137278 553596 137284 553608
rect 137336 553596 137342 553648
rect 103698 553528 103704 553580
rect 103756 553568 103762 553580
rect 141418 553568 141424 553580
rect 103756 553540 141424 553568
rect 103756 553528 103762 553540
rect 141418 553528 141424 553540
rect 141476 553528 141482 553580
rect 97810 553460 97816 553512
rect 97868 553500 97874 553512
rect 151078 553500 151084 553512
rect 97868 553472 151084 553500
rect 97868 553460 97874 553472
rect 151078 553460 151084 553472
rect 151136 553460 151142 553512
rect 112346 553392 112352 553444
rect 112404 553432 112410 553444
rect 116026 553432 116032 553444
rect 112404 553404 116032 553432
rect 112404 553392 112410 553404
rect 116026 553392 116032 553404
rect 116084 553392 116090 553444
rect 281258 553392 281264 553444
rect 281316 553432 281322 553444
rect 281316 553404 281396 553432
rect 281316 553392 281322 553404
rect 281368 553376 281396 553404
rect 128446 553324 128452 553376
rect 128504 553364 128510 553376
rect 128630 553364 128636 553376
rect 128504 553336 128636 553364
rect 128504 553324 128510 553336
rect 128630 553324 128636 553336
rect 128688 553324 128694 553376
rect 281350 553324 281356 553376
rect 281408 553324 281414 553376
rect 89622 552644 89628 552696
rect 89680 552684 89686 552696
rect 128998 552684 129004 552696
rect 89680 552656 129004 552684
rect 89680 552644 89686 552656
rect 128998 552644 129004 552656
rect 129056 552644 129062 552696
rect 271506 550604 271512 550656
rect 271564 550644 271570 550656
rect 271782 550644 271788 550656
rect 271564 550616 271788 550644
rect 271564 550604 271570 550616
rect 271782 550604 271788 550616
rect 271840 550604 271846 550656
rect 281258 550604 281264 550656
rect 281316 550644 281322 550656
rect 281350 550644 281356 550656
rect 281316 550616 281356 550644
rect 281316 550604 281322 550616
rect 281350 550604 281356 550616
rect 281408 550604 281414 550656
rect 8018 550536 8024 550588
rect 8076 550576 8082 550588
rect 8110 550576 8116 550588
rect 8076 550548 8116 550576
rect 8076 550536 8082 550548
rect 8110 550536 8116 550548
rect 8168 550536 8174 550588
rect 281074 550468 281080 550520
rect 281132 550508 281138 550520
rect 281258 550508 281264 550520
rect 281132 550480 281264 550508
rect 281132 550468 281138 550480
rect 281258 550468 281264 550480
rect 281316 550468 281322 550520
rect 85482 549856 85488 549908
rect 85540 549896 85546 549908
rect 86402 549896 86408 549908
rect 85540 549868 86408 549896
rect 85540 549856 85546 549868
rect 86402 549856 86408 549868
rect 86460 549896 86466 549908
rect 199378 549896 199384 549908
rect 86460 549868 199384 549896
rect 86460 549856 86466 549868
rect 199378 549856 199384 549868
rect 199436 549856 199442 549908
rect 271506 545776 271512 545828
rect 271564 545816 271570 545828
rect 271782 545816 271788 545828
rect 271564 545788 271788 545816
rect 271564 545776 271570 545788
rect 271782 545776 271788 545788
rect 271840 545776 271846 545828
rect 128630 543844 128636 543856
rect 128556 543816 128636 543844
rect 128556 543720 128584 543816
rect 128630 543804 128636 543816
rect 128688 543804 128694 543856
rect 128538 543668 128544 543720
rect 128596 543668 128602 543720
rect 118602 542376 118608 542428
rect 118660 542416 118666 542428
rect 155218 542416 155224 542428
rect 118660 542388 155224 542416
rect 118660 542376 118666 542388
rect 155218 542376 155224 542388
rect 155276 542376 155282 542428
rect 8110 540948 8116 541000
rect 8168 540988 8174 541000
rect 8202 540988 8208 541000
rect 8168 540960 8208 540988
rect 8168 540948 8174 540960
rect 8202 540948 8208 540960
rect 8260 540948 8266 541000
rect 271506 540948 271512 541000
rect 271564 540988 271570 541000
rect 271598 540988 271604 541000
rect 271564 540960 271604 540988
rect 271564 540948 271570 540960
rect 271598 540948 271604 540960
rect 271656 540948 271662 541000
rect 281074 540948 281080 541000
rect 281132 540988 281138 541000
rect 281258 540988 281264 541000
rect 281132 540960 281264 540988
rect 281132 540948 281138 540960
rect 281258 540948 281264 540960
rect 281316 540948 281322 541000
rect 3970 538432 3976 538484
rect 4028 538472 4034 538484
rect 4798 538472 4804 538484
rect 4028 538444 4804 538472
rect 4028 538432 4034 538444
rect 4798 538432 4804 538444
rect 4856 538432 4862 538484
rect 286962 538228 286968 538280
rect 287020 538268 287026 538280
rect 297634 538268 297640 538280
rect 287020 538240 297640 538268
rect 287020 538228 287026 538240
rect 297634 538228 297640 538240
rect 297692 538228 297698 538280
rect 117774 536800 117780 536852
rect 117832 536840 117838 536852
rect 140038 536840 140044 536852
rect 117832 536812 140044 536840
rect 117832 536800 117838 536812
rect 140038 536800 140044 536812
rect 140096 536800 140102 536852
rect 128446 534080 128452 534132
rect 128504 534120 128510 534132
rect 128504 534092 128584 534120
rect 128504 534080 128510 534092
rect 128556 534064 128584 534092
rect 281258 534080 281264 534132
rect 281316 534080 281322 534132
rect 128538 534012 128544 534064
rect 128596 534012 128602 534064
rect 281276 534052 281304 534080
rect 281350 534052 281356 534064
rect 281276 534024 281356 534052
rect 281350 534012 281356 534024
rect 281408 534012 281414 534064
rect 117774 532720 117780 532772
rect 117832 532760 117838 532772
rect 153838 532760 153844 532772
rect 117832 532732 153844 532760
rect 117832 532720 117838 532732
rect 153838 532720 153844 532732
rect 153896 532720 153902 532772
rect 294598 532720 294604 532772
rect 294656 532760 294662 532772
rect 297358 532760 297364 532772
rect 294656 532732 297364 532760
rect 294656 532720 294662 532732
rect 297358 532720 297364 532732
rect 297416 532720 297422 532772
rect 128446 531292 128452 531344
rect 128504 531332 128510 531344
rect 128538 531332 128544 531344
rect 128504 531304 128544 531332
rect 128504 531292 128510 531304
rect 128538 531292 128544 531304
rect 128596 531292 128602 531344
rect 271782 531292 271788 531344
rect 271840 531332 271846 531344
rect 271966 531332 271972 531344
rect 271840 531304 271972 531332
rect 271840 531292 271846 531304
rect 271966 531292 271972 531304
rect 272024 531292 272030 531344
rect 281258 531292 281264 531344
rect 281316 531332 281322 531344
rect 281350 531332 281356 531344
rect 281316 531304 281356 531332
rect 281316 531292 281322 531304
rect 281350 531292 281356 531304
rect 281408 531292 281414 531344
rect 117958 529864 117964 529916
rect 118016 529904 118022 529916
rect 119338 529904 119344 529916
rect 118016 529876 119344 529904
rect 118016 529864 118022 529876
rect 119338 529864 119344 529876
rect 119396 529864 119402 529916
rect 118602 525036 118608 525088
rect 118660 525076 118666 525088
rect 128354 525076 128360 525088
rect 118660 525048 128360 525076
rect 118660 525036 118666 525048
rect 128354 525036 128360 525048
rect 128412 525076 128418 525088
rect 129274 525076 129280 525088
rect 128412 525048 129280 525076
rect 128412 525036 128418 525048
rect 129274 525036 129280 525048
rect 129332 525036 129338 525088
rect 271782 524492 271788 524544
rect 271840 524492 271846 524544
rect 281258 524492 281264 524544
rect 281316 524492 281322 524544
rect 70210 524424 70216 524476
rect 70268 524464 70274 524476
rect 82814 524464 82820 524476
rect 70268 524436 82820 524464
rect 70268 524424 70274 524436
rect 82814 524424 82820 524436
rect 82872 524424 82878 524476
rect 128446 524424 128452 524476
rect 128504 524424 128510 524476
rect 128464 524328 128492 524424
rect 271800 524408 271828 524492
rect 281276 524408 281304 524492
rect 271782 524356 271788 524408
rect 271840 524356 271846 524408
rect 281258 524356 281264 524408
rect 281316 524356 281322 524408
rect 128630 524328 128636 524340
rect 128464 524300 128636 524328
rect 128630 524288 128636 524300
rect 128688 524288 128694 524340
rect 8202 521636 8208 521688
rect 8260 521676 8266 521688
rect 8386 521676 8392 521688
rect 8260 521648 8392 521676
rect 8260 521636 8266 521648
rect 8386 521636 8392 521648
rect 8444 521636 8450 521688
rect 280062 521636 280068 521688
rect 280120 521676 280126 521688
rect 297542 521676 297548 521688
rect 280120 521648 297548 521676
rect 280120 521636 280126 521648
rect 297542 521636 297548 521648
rect 297600 521636 297606 521688
rect 128446 521568 128452 521620
rect 128504 521608 128510 521620
rect 129090 521608 129096 521620
rect 128504 521580 129096 521608
rect 128504 521568 128510 521580
rect 129090 521568 129096 521580
rect 129148 521568 129154 521620
rect 293954 521568 293960 521620
rect 294012 521608 294018 521620
rect 294598 521608 294604 521620
rect 294012 521580 294604 521608
rect 294012 521568 294018 521580
rect 294598 521568 294604 521580
rect 294656 521568 294662 521620
rect 85298 521228 85304 521280
rect 85356 521268 85362 521280
rect 293954 521268 293960 521280
rect 85356 521240 293960 521268
rect 85356 521228 85362 521240
rect 293954 521228 293960 521240
rect 294012 521228 294018 521280
rect 199746 521092 199752 521144
rect 199804 521132 199810 521144
rect 222378 521132 222384 521144
rect 199804 521104 222384 521132
rect 199804 521092 199810 521104
rect 222378 521092 222384 521104
rect 222436 521092 222442 521144
rect 199838 521024 199844 521076
rect 199896 521064 199902 521076
rect 222562 521064 222568 521076
rect 199896 521036 222568 521064
rect 199896 521024 199902 521036
rect 222562 521024 222568 521036
rect 222620 521024 222626 521076
rect 196434 520956 196440 521008
rect 196492 520996 196498 521008
rect 222470 520996 222476 521008
rect 196492 520968 222476 520996
rect 196492 520956 196498 520968
rect 222470 520956 222476 520968
rect 222528 520956 222534 521008
rect 117314 520888 117320 520940
rect 117372 520928 117378 520940
rect 128446 520928 128452 520940
rect 117372 520900 128452 520928
rect 117372 520888 117378 520900
rect 128446 520888 128452 520900
rect 128504 520888 128510 520940
rect 195054 520888 195060 520940
rect 195112 520928 195118 520940
rect 222654 520928 222660 520940
rect 195112 520900 222660 520928
rect 195112 520888 195118 520900
rect 222654 520888 222660 520900
rect 222712 520888 222718 520940
rect 128354 518916 128360 518968
rect 128412 518956 128418 518968
rect 128630 518956 128636 518968
rect 128412 518928 128636 518956
rect 128412 518916 128418 518928
rect 128630 518916 128636 518928
rect 128688 518916 128694 518968
rect 278682 518916 278688 518968
rect 278740 518956 278746 518968
rect 297450 518956 297456 518968
rect 278740 518928 297456 518956
rect 278740 518916 278746 518928
rect 297450 518916 297456 518928
rect 297508 518916 297514 518968
rect 89346 518848 89352 518900
rect 89404 518888 89410 518900
rect 122558 518888 122564 518900
rect 89404 518860 122564 518888
rect 89404 518848 89410 518860
rect 122558 518848 122564 518860
rect 122616 518848 122622 518900
rect 122834 518848 122840 518900
rect 122892 518888 122898 518900
rect 129734 518888 129740 518900
rect 122892 518860 129740 518888
rect 122892 518848 122898 518860
rect 129734 518848 129740 518860
rect 129792 518848 129798 518900
rect 109586 518780 109592 518832
rect 109644 518820 109650 518832
rect 113818 518820 113824 518832
rect 109644 518792 113824 518820
rect 109644 518780 109650 518792
rect 113818 518780 113824 518792
rect 113876 518820 113882 518832
rect 115198 518820 115204 518832
rect 113876 518792 115204 518820
rect 113876 518780 113882 518792
rect 115198 518780 115204 518792
rect 115256 518780 115262 518832
rect 127710 518820 127716 518832
rect 122852 518792 127716 518820
rect 99282 518752 99288 518764
rect 91756 518724 99288 518752
rect 86586 518644 86592 518696
rect 86644 518684 86650 518696
rect 86644 518656 89576 518684
rect 86644 518644 86650 518656
rect 89548 518616 89576 518656
rect 91756 518616 91784 518724
rect 99282 518712 99288 518724
rect 99340 518712 99346 518764
rect 99374 518712 99380 518764
rect 99432 518752 99438 518764
rect 122466 518752 122472 518764
rect 99432 518724 104940 518752
rect 122379 518724 122472 518752
rect 99432 518712 99438 518724
rect 104912 518684 104940 518724
rect 122466 518712 122472 518724
rect 122524 518752 122530 518764
rect 122852 518752 122880 518792
rect 127710 518780 127716 518792
rect 127768 518780 127774 518832
rect 122524 518724 122880 518752
rect 122524 518712 122530 518724
rect 109034 518684 109040 518696
rect 104912 518656 109040 518684
rect 109034 518644 109040 518656
rect 109092 518644 109098 518696
rect 109126 518644 109132 518696
rect 109184 518684 109190 518696
rect 109184 518656 115980 518684
rect 109184 518644 109190 518656
rect 89548 518588 91784 518616
rect 115952 518616 115980 518656
rect 122484 518616 122512 518712
rect 115952 518588 122512 518616
rect 129734 518508 129740 518560
rect 129792 518548 129798 518560
rect 130378 518548 130384 518560
rect 129792 518520 130384 518548
rect 129792 518508 129798 518520
rect 130378 518508 130384 518520
rect 130436 518508 130442 518560
rect 97994 518372 98000 518424
rect 98052 518412 98058 518424
rect 127618 518412 127624 518424
rect 98052 518384 127624 518412
rect 98052 518372 98058 518384
rect 127618 518372 127624 518384
rect 127676 518372 127682 518424
rect 106642 518304 106648 518356
rect 106700 518344 106706 518356
rect 144178 518344 144184 518356
rect 106700 518316 144184 518344
rect 106700 518304 106706 518316
rect 144178 518304 144184 518316
rect 144236 518304 144242 518356
rect 100938 518236 100944 518288
rect 100996 518276 101002 518288
rect 152458 518276 152464 518288
rect 100996 518248 152464 518276
rect 100996 518236 101002 518248
rect 152458 518236 152464 518248
rect 152516 518236 152522 518288
rect 196342 518236 196348 518288
rect 196400 518276 196406 518288
rect 218974 518276 218980 518288
rect 196400 518248 218980 518276
rect 196400 518236 196406 518248
rect 218974 518236 218980 518248
rect 219032 518236 219038 518288
rect 92290 518168 92296 518220
rect 92348 518208 92354 518220
rect 127066 518208 127072 518220
rect 92348 518180 127072 518208
rect 92348 518168 92354 518180
rect 127066 518168 127072 518180
rect 127124 518208 127130 518220
rect 297358 518208 297364 518220
rect 127124 518180 297364 518208
rect 127124 518168 127130 518180
rect 297358 518168 297364 518180
rect 297416 518168 297422 518220
rect 205634 517488 205640 517540
rect 205692 517528 205698 517540
rect 206646 517528 206652 517540
rect 205692 517500 206652 517528
rect 205692 517488 205698 517500
rect 206646 517488 206652 517500
rect 206704 517488 206710 517540
rect 505738 517488 505744 517540
rect 505796 517528 505802 517540
rect 506842 517528 506848 517540
rect 505796 517500 506848 517528
rect 505796 517488 505802 517500
rect 506842 517488 506848 517500
rect 506900 517488 506906 517540
rect 282730 516128 282736 516180
rect 282788 516168 282794 516180
rect 297450 516168 297456 516180
rect 282788 516140 297456 516168
rect 282788 516128 282794 516140
rect 297450 516128 297456 516140
rect 297508 516128 297514 516180
rect 271782 514808 271788 514820
rect 271708 514780 271788 514808
rect 271708 514752 271736 514780
rect 271782 514768 271788 514780
rect 271840 514768 271846 514820
rect 281258 514768 281264 514820
rect 281316 514768 281322 514820
rect 271690 514700 271696 514752
rect 271748 514700 271754 514752
rect 281276 514740 281304 514768
rect 281350 514740 281356 514752
rect 281276 514712 281356 514740
rect 281350 514700 281356 514712
rect 281408 514700 281414 514752
rect 271690 511980 271696 512032
rect 271748 512020 271754 512032
rect 271782 512020 271788 512032
rect 271748 511992 271788 512020
rect 271748 511980 271754 511992
rect 271782 511980 271788 511992
rect 271840 511980 271846 512032
rect 281258 511980 281264 512032
rect 281316 512020 281322 512032
rect 281350 512020 281356 512032
rect 281316 511992 281356 512020
rect 281316 511980 281322 511992
rect 281350 511980 281356 511992
rect 281408 511980 281414 512032
rect 281074 511844 281080 511896
rect 281132 511884 281138 511896
rect 281258 511884 281264 511896
rect 281132 511856 281264 511884
rect 281132 511844 281138 511856
rect 281258 511844 281264 511856
rect 281316 511844 281322 511896
rect 293770 509260 293776 509312
rect 293828 509300 293834 509312
rect 296714 509300 296720 509312
rect 293828 509272 296720 509300
rect 293828 509260 293834 509272
rect 296714 509260 296720 509272
rect 296772 509260 296778 509312
rect 128354 509192 128360 509244
rect 128412 509232 128418 509244
rect 128630 509232 128636 509244
rect 128412 509204 128636 509232
rect 128412 509192 128418 509204
rect 128630 509192 128636 509204
rect 128688 509192 128694 509244
rect 271506 507152 271512 507204
rect 271564 507192 271570 507204
rect 271782 507192 271788 507204
rect 271564 507164 271788 507192
rect 271564 507152 271570 507164
rect 271782 507152 271788 507164
rect 271840 507152 271846 507204
rect 380342 506608 380348 506660
rect 380400 506648 380406 506660
rect 380618 506648 380624 506660
rect 380400 506620 380624 506648
rect 380400 506608 380406 506620
rect 380618 506608 380624 506620
rect 380676 506608 380682 506660
rect 191098 506472 191104 506524
rect 191156 506512 191162 506524
rect 296714 506512 296720 506524
rect 191156 506484 296720 506512
rect 191156 506472 191162 506484
rect 296714 506472 296720 506484
rect 296772 506472 296778 506524
rect 297174 505044 297180 505096
rect 297232 505084 297238 505096
rect 298002 505084 298008 505096
rect 297232 505056 298008 505084
rect 297232 505044 297238 505056
rect 298002 505044 298008 505056
rect 298060 505044 298066 505096
rect 8202 502324 8208 502376
rect 8260 502364 8266 502376
rect 8386 502364 8392 502376
rect 8260 502336 8392 502364
rect 8260 502324 8266 502336
rect 8386 502324 8392 502336
rect 8444 502324 8450 502376
rect 271506 502324 271512 502376
rect 271564 502364 271570 502376
rect 271598 502364 271604 502376
rect 271564 502336 271604 502364
rect 271564 502324 271570 502336
rect 271598 502324 271604 502336
rect 271656 502324 271662 502376
rect 281074 502324 281080 502376
rect 281132 502364 281138 502376
rect 281258 502364 281264 502376
rect 281132 502336 281264 502364
rect 281132 502324 281138 502336
rect 281258 502324 281264 502336
rect 281316 502324 281322 502376
rect 96522 500896 96528 500948
rect 96580 500936 96586 500948
rect 380342 500936 380348 500948
rect 96580 500908 380348 500936
rect 96580 500896 96586 500908
rect 380342 500896 380348 500908
rect 380400 500896 380406 500948
rect 103514 500828 103520 500880
rect 103572 500868 103578 500880
rect 104802 500868 104808 500880
rect 103572 500840 104808 500868
rect 103572 500828 103578 500840
rect 104802 500828 104808 500840
rect 104860 500868 104866 500880
rect 377674 500868 377680 500880
rect 104860 500840 377680 500868
rect 104860 500828 104866 500840
rect 377674 500828 377680 500840
rect 377732 500828 377738 500880
rect 129366 500420 129372 500472
rect 129424 500460 129430 500472
rect 377398 500460 377404 500472
rect 129424 500432 377404 500460
rect 129424 500420 129430 500432
rect 377398 500420 377404 500432
rect 377456 500420 377462 500472
rect 130838 500352 130844 500404
rect 130896 500392 130902 500404
rect 380618 500392 380624 500404
rect 130896 500364 380624 500392
rect 130896 500352 130902 500364
rect 380618 500352 380624 500364
rect 380676 500352 380682 500404
rect 130654 500284 130660 500336
rect 130712 500324 130718 500336
rect 580442 500324 580448 500336
rect 130712 500296 580448 500324
rect 130712 500284 130718 500296
rect 580442 500284 580448 500296
rect 580500 500284 580506 500336
rect 70302 500216 70308 500268
rect 70360 500256 70366 500268
rect 95234 500256 95240 500268
rect 70360 500228 95240 500256
rect 70360 500216 70366 500228
rect 95234 500216 95240 500228
rect 95292 500256 95298 500268
rect 96522 500256 96528 500268
rect 95292 500228 96528 500256
rect 95292 500216 95298 500228
rect 96522 500216 96528 500228
rect 96580 500216 96586 500268
rect 130746 500216 130752 500268
rect 130804 500256 130810 500268
rect 580534 500256 580540 500268
rect 130804 500228 580540 500256
rect 130804 500216 130810 500228
rect 580534 500216 580540 500228
rect 580592 500216 580598 500268
rect 128354 499536 128360 499588
rect 128412 499576 128418 499588
rect 128630 499576 128636 499588
rect 128412 499548 128636 499576
rect 128412 499536 128418 499548
rect 128630 499536 128636 499548
rect 128688 499536 128694 499588
rect 298830 499400 298836 499452
rect 298888 499440 298894 499452
rect 302418 499440 302424 499452
rect 298888 499412 302424 499440
rect 298888 499400 298894 499412
rect 302418 499400 302424 499412
rect 302476 499400 302482 499452
rect 324222 499060 324228 499112
rect 324280 499100 324286 499112
rect 379054 499100 379060 499112
rect 324280 499072 379060 499100
rect 324280 499060 324286 499072
rect 379054 499060 379060 499072
rect 379112 499060 379118 499112
rect 298922 498992 298928 499044
rect 298980 499032 298986 499044
rect 310514 499032 310520 499044
rect 298980 499004 310520 499032
rect 298980 498992 298986 499004
rect 310514 498992 310520 499004
rect 310572 498992 310578 499044
rect 321462 498992 321468 499044
rect 321520 499032 321526 499044
rect 378962 499032 378968 499044
rect 321520 499004 378968 499032
rect 321520 498992 321526 499004
rect 378962 498992 378968 499004
rect 379020 498992 379026 499044
rect 300302 498924 300308 498976
rect 300360 498964 300366 498976
rect 311894 498964 311900 498976
rect 300360 498936 311900 498964
rect 300360 498924 300366 498936
rect 311894 498924 311900 498936
rect 311952 498924 311958 498976
rect 317322 498924 317328 498976
rect 317380 498964 317386 498976
rect 377582 498964 377588 498976
rect 317380 498936 377588 498964
rect 317380 498924 317386 498936
rect 377582 498924 377588 498936
rect 377640 498924 377646 498976
rect 309042 498856 309048 498908
rect 309100 498896 309106 498908
rect 377490 498896 377496 498908
rect 309100 498868 377496 498896
rect 309100 498856 309106 498868
rect 377490 498856 377496 498868
rect 377548 498856 377554 498908
rect 118050 498788 118056 498840
rect 118108 498828 118114 498840
rect 302050 498828 302056 498840
rect 118108 498800 302056 498828
rect 118108 498788 118114 498800
rect 302050 498788 302056 498800
rect 302108 498788 302114 498840
rect 375282 498788 375288 498840
rect 375340 498828 375346 498840
rect 478874 498828 478880 498840
rect 375340 498800 478880 498828
rect 375340 498788 375346 498800
rect 478874 498788 478880 498800
rect 478932 498788 478938 498840
rect 131850 498176 131856 498228
rect 131908 498216 131914 498228
rect 579890 498216 579896 498228
rect 131908 498188 579896 498216
rect 131908 498176 131914 498188
rect 579890 498176 579896 498188
rect 579948 498176 579954 498228
rect 116026 498040 116032 498092
rect 116084 498080 116090 498092
rect 347314 498080 347320 498092
rect 116084 498052 347320 498080
rect 116084 498040 116090 498052
rect 347314 498040 347320 498052
rect 347372 498040 347378 498092
rect 120718 497972 120724 498024
rect 120776 498012 120782 498024
rect 121362 498012 121368 498024
rect 120776 497984 121368 498012
rect 120776 497972 120782 497984
rect 121362 497972 121368 497984
rect 121420 498012 121426 498024
rect 338850 498012 338856 498024
rect 121420 497984 338856 498012
rect 121420 497972 121426 497984
rect 338850 497972 338856 497984
rect 338908 497972 338914 498024
rect 128262 497904 128268 497956
rect 128320 497944 128326 497956
rect 334434 497944 334440 497956
rect 128320 497916 334440 497944
rect 128320 497904 128326 497916
rect 334434 497904 334440 497916
rect 334492 497904 334498 497956
rect 335998 497904 336004 497956
rect 336056 497944 336062 497956
rect 349338 497944 349344 497956
rect 336056 497916 349344 497944
rect 336056 497904 336062 497916
rect 349338 497904 349344 497916
rect 349396 497904 349402 497956
rect 111702 497836 111708 497888
rect 111760 497876 111766 497888
rect 115290 497876 115296 497888
rect 111760 497848 115296 497876
rect 111760 497836 111766 497848
rect 115290 497836 115296 497848
rect 115348 497876 115354 497888
rect 313274 497876 313280 497888
rect 115348 497848 313280 497876
rect 115348 497836 115354 497848
rect 313274 497836 313280 497848
rect 313332 497836 313338 497888
rect 318702 497836 318708 497888
rect 318760 497876 318766 497888
rect 355778 497876 355784 497888
rect 318760 497848 355784 497876
rect 318760 497836 318766 497848
rect 355778 497836 355784 497848
rect 355836 497836 355842 497888
rect 155218 497768 155224 497820
rect 155276 497808 155282 497820
rect 319714 497808 319720 497820
rect 155276 497780 319720 497808
rect 155276 497768 155282 497780
rect 319714 497768 319720 497780
rect 319772 497768 319778 497820
rect 320082 497768 320088 497820
rect 320140 497808 320146 497820
rect 357986 497808 357992 497820
rect 320140 497780 357992 497808
rect 320140 497768 320146 497780
rect 357986 497768 357992 497780
rect 358044 497768 358050 497820
rect 284202 497700 284208 497752
rect 284260 497740 284266 497752
rect 368474 497740 368480 497752
rect 284260 497712 368480 497740
rect 284260 497700 284266 497712
rect 368474 497700 368480 497712
rect 368532 497700 368538 497752
rect 291010 497632 291016 497684
rect 291068 497672 291074 497684
rect 377122 497672 377128 497684
rect 291068 497644 377128 497672
rect 291068 497632 291074 497644
rect 377122 497632 377128 497644
rect 377180 497632 377186 497684
rect 108942 497564 108948 497616
rect 109000 497604 109006 497616
rect 116026 497604 116032 497616
rect 109000 497576 116032 497604
rect 109000 497564 109006 497576
rect 116026 497564 116032 497576
rect 116084 497564 116090 497616
rect 127618 497564 127624 497616
rect 127676 497604 127682 497616
rect 128262 497604 128268 497616
rect 127676 497576 128268 497604
rect 127676 497564 127682 497576
rect 128262 497564 128268 497576
rect 128320 497564 128326 497616
rect 281074 497564 281080 497616
rect 281132 497604 281138 497616
rect 281258 497604 281264 497616
rect 281132 497576 281264 497604
rect 281132 497564 281138 497576
rect 281258 497564 281264 497576
rect 281316 497564 281322 497616
rect 284110 497564 284116 497616
rect 284168 497604 284174 497616
rect 374914 497604 374920 497616
rect 284168 497576 374920 497604
rect 284168 497564 284174 497576
rect 374914 497564 374920 497576
rect 374972 497564 374978 497616
rect 83826 497496 83832 497548
rect 83884 497536 83890 497548
rect 127158 497536 127164 497548
rect 83884 497508 127164 497536
rect 83884 497496 83890 497508
rect 127158 497496 127164 497508
rect 127216 497536 127222 497548
rect 360010 497536 360016 497548
rect 127216 497508 360016 497536
rect 127216 497496 127222 497508
rect 360010 497496 360016 497508
rect 360068 497496 360074 497548
rect 111794 497428 111800 497480
rect 111852 497468 111858 497480
rect 125962 497468 125968 497480
rect 111852 497440 125968 497468
rect 111852 497428 111858 497440
rect 125962 497428 125968 497440
rect 126020 497468 126026 497480
rect 372706 497468 372712 497480
rect 126020 497440 372712 497468
rect 126020 497428 126026 497440
rect 372706 497428 372712 497440
rect 372764 497428 372770 497480
rect 289630 497360 289636 497412
rect 289688 497400 289694 497412
rect 366450 497400 366456 497412
rect 289688 497372 366456 497400
rect 289688 497360 289694 497372
rect 366450 497360 366456 497372
rect 366508 497360 366514 497412
rect 285582 497292 285588 497344
rect 285640 497332 285646 497344
rect 345106 497332 345112 497344
rect 285640 497304 345112 497332
rect 285640 497292 285646 497304
rect 345106 497292 345112 497304
rect 345164 497292 345170 497344
rect 292390 497224 292396 497276
rect 292448 497264 292454 497276
rect 351546 497264 351552 497276
rect 292448 497236 351552 497264
rect 292448 497224 292454 497236
rect 351546 497224 351552 497236
rect 351604 497224 351610 497276
rect 275830 497156 275836 497208
rect 275888 497196 275894 497208
rect 306834 497196 306840 497208
rect 275888 497168 306840 497196
rect 275888 497156 275894 497168
rect 306834 497156 306840 497168
rect 306892 497156 306898 497208
rect 307018 497156 307024 497208
rect 307076 497196 307082 497208
rect 362218 497196 362224 497208
rect 307076 497168 362224 497196
rect 307076 497156 307082 497168
rect 362218 497156 362224 497168
rect 362276 497156 362282 497208
rect 277302 497088 277308 497140
rect 277360 497128 277366 497140
rect 317506 497128 317512 497140
rect 277360 497100 317512 497128
rect 277360 497088 277366 497100
rect 317506 497088 317512 497100
rect 317564 497088 317570 497140
rect 334618 497088 334624 497140
rect 334676 497128 334682 497140
rect 343082 497128 343088 497140
rect 334676 497100 343088 497128
rect 334676 497088 334682 497100
rect 343082 497088 343088 497100
rect 343140 497088 343146 497140
rect 288250 497020 288256 497072
rect 288308 497060 288314 497072
rect 321738 497060 321744 497072
rect 288308 497032 321744 497060
rect 288308 497020 288314 497032
rect 321738 497020 321744 497032
rect 321796 497020 321802 497072
rect 307570 496952 307576 497004
rect 307628 496992 307634 497004
rect 315022 496992 315028 497004
rect 307628 496964 315028 496992
rect 307628 496952 307634 496964
rect 315022 496952 315028 496964
rect 315080 496952 315086 497004
rect 315298 496952 315304 497004
rect 315356 496992 315362 497004
rect 323946 496992 323952 497004
rect 315356 496964 323952 496992
rect 315356 496952 315362 496964
rect 323946 496952 323952 496964
rect 324004 496952 324010 497004
rect 155218 496884 155224 496936
rect 155276 496924 155282 496936
rect 155862 496924 155868 496936
rect 155276 496896 155868 496924
rect 155276 496884 155282 496896
rect 155862 496884 155868 496896
rect 155920 496884 155926 496936
rect 304810 496884 304816 496936
rect 304868 496924 304874 496936
rect 309318 496924 309324 496936
rect 304868 496896 309324 496924
rect 304868 496884 304874 496896
rect 309318 496884 309324 496896
rect 309376 496884 309382 496936
rect 324958 496884 324964 496936
rect 325016 496924 325022 496936
rect 328178 496924 328184 496936
rect 325016 496896 328184 496924
rect 325016 496884 325022 496896
rect 328178 496884 328184 496896
rect 328236 496884 328242 496936
rect 331858 496884 331864 496936
rect 331916 496924 331922 496936
rect 336642 496924 336648 496936
rect 331916 496896 336648 496924
rect 331916 496884 331922 496896
rect 336642 496884 336648 496896
rect 336700 496884 336706 496936
rect 129182 496816 129188 496868
rect 129240 496856 129246 496868
rect 364242 496856 364248 496868
rect 129240 496828 364248 496856
rect 129240 496816 129246 496828
rect 364242 496816 364248 496828
rect 364300 496816 364306 496868
rect 297174 495456 297180 495508
rect 297232 495496 297238 495508
rect 298002 495496 298008 495508
rect 297232 495468 298008 495496
rect 297232 495456 297238 495468
rect 298002 495456 298008 495468
rect 298060 495456 298066 495508
rect 308858 492736 308864 492788
rect 308916 492776 308922 492788
rect 309042 492776 309048 492788
rect 308916 492748 309048 492776
rect 308916 492736 308922 492748
rect 309042 492736 309048 492748
rect 309100 492736 309106 492788
rect 302050 492600 302056 492652
rect 302108 492640 302114 492652
rect 302142 492640 302148 492652
rect 302108 492612 302148 492640
rect 302108 492600 302114 492612
rect 302142 492600 302148 492612
rect 302200 492600 302206 492652
rect 301958 491240 301964 491292
rect 302016 491280 302022 491292
rect 302142 491280 302148 491292
rect 302016 491252 302148 491280
rect 302016 491240 302022 491252
rect 302142 491240 302148 491252
rect 302200 491240 302206 491292
rect 299566 490560 299572 490612
rect 299624 490600 299630 490612
rect 300578 490600 300584 490612
rect 299624 490572 300584 490600
rect 299624 490560 299630 490572
rect 300578 490560 300584 490572
rect 300636 490560 300642 490612
rect 128354 489812 128360 489864
rect 128412 489852 128418 489864
rect 128630 489852 128636 489864
rect 128412 489824 128636 489852
rect 128412 489812 128418 489824
rect 128630 489812 128636 489824
rect 128688 489812 128694 489864
rect 271506 487772 271512 487824
rect 271564 487812 271570 487824
rect 271782 487812 271788 487824
rect 271564 487784 271788 487812
rect 271564 487772 271570 487784
rect 271782 487772 271788 487784
rect 271840 487772 271846 487824
rect 281258 485868 281264 485920
rect 281316 485868 281322 485920
rect 8110 485800 8116 485852
rect 8168 485800 8174 485852
rect 8128 485772 8156 485800
rect 281276 485784 281304 485868
rect 438302 485800 438308 485852
rect 438360 485840 438366 485852
rect 580166 485840 580172 485852
rect 438360 485812 580172 485840
rect 438360 485800 438366 485812
rect 580166 485800 580172 485812
rect 580224 485800 580230 485852
rect 8202 485772 8208 485784
rect 8128 485744 8208 485772
rect 8202 485732 8208 485744
rect 8260 485732 8266 485784
rect 281258 485732 281264 485784
rect 281316 485732 281322 485784
rect 271506 483080 271512 483132
rect 271564 483120 271570 483132
rect 271690 483120 271696 483132
rect 271564 483092 271696 483120
rect 271564 483080 271570 483092
rect 271690 483080 271696 483092
rect 271748 483080 271754 483132
rect 7926 482944 7932 482996
rect 7984 482984 7990 482996
rect 8202 482984 8208 482996
rect 7984 482956 8208 482984
rect 7984 482944 7990 482956
rect 8202 482944 8208 482956
rect 8260 482944 8266 482996
rect 271690 482944 271696 482996
rect 271748 482984 271754 482996
rect 271782 482984 271788 482996
rect 271748 482956 271788 482984
rect 271748 482944 271754 482956
rect 271782 482944 271788 482956
rect 271840 482944 271846 482996
rect 301866 481652 301872 481704
rect 301924 481692 301930 481704
rect 301958 481692 301964 481704
rect 301924 481664 301964 481692
rect 301924 481652 301930 481664
rect 301958 481652 301964 481664
rect 302016 481652 302022 481704
rect 308766 481584 308772 481636
rect 308824 481624 308830 481636
rect 308858 481624 308864 481636
rect 308824 481596 308864 481624
rect 308824 481584 308830 481596
rect 308858 481584 308864 481596
rect 308916 481584 308922 481636
rect 3142 481040 3148 481092
rect 3200 481080 3206 481092
rect 4890 481080 4896 481092
rect 3200 481052 4896 481080
rect 3200 481040 3206 481052
rect 4890 481040 4896 481052
rect 4948 481040 4954 481092
rect 128354 480292 128360 480344
rect 128412 480332 128418 480344
rect 128630 480332 128636 480344
rect 128412 480304 128636 480332
rect 128412 480292 128418 480304
rect 128630 480292 128636 480304
rect 128688 480292 128694 480344
rect 271782 476116 271788 476128
rect 271708 476088 271788 476116
rect 271708 476060 271736 476088
rect 271782 476076 271788 476088
rect 271840 476076 271846 476128
rect 281258 476076 281264 476128
rect 281316 476116 281322 476128
rect 281350 476116 281356 476128
rect 281316 476088 281356 476116
rect 281316 476076 281322 476088
rect 281350 476076 281356 476088
rect 281408 476076 281414 476128
rect 271690 476008 271696 476060
rect 271748 476008 271754 476060
rect 281258 473356 281264 473408
rect 281316 473396 281322 473408
rect 281350 473396 281356 473408
rect 281316 473368 281356 473396
rect 281316 473356 281322 473368
rect 281350 473356 281356 473368
rect 281408 473356 281414 473408
rect 308858 473356 308864 473408
rect 308916 473356 308922 473408
rect 308766 473288 308772 473340
rect 308824 473328 308830 473340
rect 308876 473328 308904 473356
rect 308824 473300 308904 473328
rect 308824 473288 308830 473300
rect 302050 469072 302056 469124
rect 302108 469072 302114 469124
rect 302068 468988 302096 469072
rect 302050 468936 302056 468988
rect 302108 468936 302114 468988
rect 271506 468460 271512 468512
rect 271564 468500 271570 468512
rect 271782 468500 271788 468512
rect 271564 468472 271788 468500
rect 271564 468460 271570 468472
rect 271782 468460 271788 468472
rect 271840 468460 271846 468512
rect 281258 466488 281264 466540
rect 281316 466488 281322 466540
rect 8110 466420 8116 466472
rect 8168 466420 8174 466472
rect 8128 466392 8156 466420
rect 281276 466404 281304 466488
rect 8202 466392 8208 466404
rect 8128 466364 8208 466392
rect 8202 466352 8208 466364
rect 8260 466352 8266 466404
rect 281258 466352 281264 466404
rect 281316 466352 281322 466404
rect 271506 463768 271512 463820
rect 271564 463808 271570 463820
rect 271690 463808 271696 463820
rect 271564 463780 271696 463808
rect 271564 463768 271570 463780
rect 271690 463768 271696 463780
rect 271748 463768 271754 463820
rect 271690 463632 271696 463684
rect 271748 463672 271754 463684
rect 271782 463672 271788 463684
rect 271748 463644 271788 463672
rect 271748 463632 271754 463644
rect 271782 463632 271788 463644
rect 271840 463632 271846 463684
rect 306834 463632 306840 463684
rect 306892 463672 306898 463684
rect 307018 463672 307024 463684
rect 306892 463644 307024 463672
rect 306892 463632 306898 463644
rect 307018 463632 307024 463644
rect 307076 463632 307082 463684
rect 130562 462340 130568 462392
rect 130620 462380 130626 462392
rect 580166 462380 580172 462392
rect 130620 462352 580172 462380
rect 130620 462340 130626 462352
rect 580166 462340 580172 462352
rect 580224 462340 580230 462392
rect 281074 458804 281080 458856
rect 281132 458844 281138 458856
rect 281258 458844 281264 458856
rect 281132 458816 281264 458844
rect 281132 458804 281138 458816
rect 281258 458804 281264 458816
rect 281316 458804 281322 458856
rect 271782 456804 271788 456816
rect 271708 456776 271788 456804
rect 271708 456748 271736 456776
rect 271782 456764 271788 456776
rect 271840 456764 271846 456816
rect 271690 456696 271696 456748
rect 271748 456696 271754 456748
rect 7834 453976 7840 454028
rect 7892 454016 7898 454028
rect 8018 454016 8024 454028
rect 7892 453988 8024 454016
rect 7892 453976 7898 453988
rect 8018 453976 8024 453988
rect 8076 453976 8082 454028
rect 3234 451324 3240 451376
rect 3292 451364 3298 451376
rect 261294 451364 261300 451376
rect 3292 451336 261300 451364
rect 3292 451324 3298 451336
rect 261294 451324 261300 451336
rect 261352 451324 261358 451376
rect 134058 451256 134064 451308
rect 134116 451296 134122 451308
rect 579890 451296 579896 451308
rect 134116 451268 579896 451296
rect 134116 451256 134122 451268
rect 579890 451256 579896 451268
rect 579948 451256 579954 451308
rect 271506 449148 271512 449200
rect 271564 449188 271570 449200
rect 271782 449188 271788 449200
rect 271564 449160 271788 449188
rect 271564 449148 271570 449160
rect 271782 449148 271788 449160
rect 271840 449148 271846 449200
rect 302050 448536 302056 448588
rect 302108 448576 302114 448588
rect 302234 448576 302240 448588
rect 302108 448548 302240 448576
rect 302108 448536 302114 448548
rect 302234 448536 302240 448548
rect 302292 448536 302298 448588
rect 281258 447176 281264 447228
rect 281316 447176 281322 447228
rect 281276 447092 281304 447176
rect 261294 447040 261300 447092
rect 261352 447080 261358 447092
rect 265986 447080 265992 447092
rect 261352 447052 265992 447080
rect 261352 447040 261358 447052
rect 265986 447040 265992 447052
rect 266044 447040 266050 447092
rect 281258 447040 281264 447092
rect 281316 447040 281322 447092
rect 271506 444456 271512 444508
rect 271564 444496 271570 444508
rect 271690 444496 271696 444508
rect 271564 444468 271696 444496
rect 271564 444456 271570 444468
rect 271690 444456 271696 444468
rect 271748 444456 271754 444508
rect 7834 444388 7840 444440
rect 7892 444428 7898 444440
rect 7926 444428 7932 444440
rect 7892 444400 7932 444428
rect 7892 444388 7898 444400
rect 7926 444388 7932 444400
rect 7984 444388 7990 444440
rect 265986 444320 265992 444372
rect 266044 444360 266050 444372
rect 266078 444360 266084 444372
rect 266044 444332 266084 444360
rect 266044 444320 266050 444332
rect 266078 444320 266084 444332
rect 266136 444320 266142 444372
rect 271690 444320 271696 444372
rect 271748 444360 271754 444372
rect 271782 444360 271788 444372
rect 271748 444332 271788 444360
rect 271748 444320 271754 444332
rect 271782 444320 271788 444332
rect 271840 444320 271846 444372
rect 306834 444320 306840 444372
rect 306892 444360 306898 444372
rect 307018 444360 307024 444372
rect 306892 444332 307024 444360
rect 306892 444320 306898 444332
rect 307018 444320 307024 444332
rect 307076 444320 307082 444372
rect 308766 442960 308772 443012
rect 308824 443000 308830 443012
rect 308858 443000 308864 443012
rect 308824 442972 308864 443000
rect 308824 442960 308830 442972
rect 308858 442960 308864 442972
rect 308916 442960 308922 443012
rect 281074 439492 281080 439544
rect 281132 439532 281138 439544
rect 281258 439532 281264 439544
rect 281132 439504 281264 439532
rect 281132 439492 281138 439504
rect 281258 439492 281264 439504
rect 281316 439492 281322 439544
rect 301866 438812 301872 438864
rect 301924 438852 301930 438864
rect 302050 438852 302056 438864
rect 301924 438824 302056 438852
rect 301924 438812 301930 438824
rect 302050 438812 302056 438824
rect 302108 438812 302114 438864
rect 266078 437492 266084 437504
rect 266004 437464 266084 437492
rect 266004 437436 266032 437464
rect 266078 437452 266084 437464
rect 266136 437452 266142 437504
rect 271782 437492 271788 437504
rect 271708 437464 271788 437492
rect 271708 437436 271736 437464
rect 271782 437452 271788 437464
rect 271840 437452 271846 437504
rect 265986 437384 265992 437436
rect 266044 437384 266050 437436
rect 271690 437384 271696 437436
rect 271748 437384 271754 437436
rect 306834 434732 306840 434784
rect 306892 434772 306898 434784
rect 307018 434772 307024 434784
rect 306892 434744 307024 434772
rect 306892 434732 306898 434744
rect 307018 434732 307024 434744
rect 307076 434732 307082 434784
rect 128354 431876 128360 431928
rect 128412 431916 128418 431928
rect 128630 431916 128636 431928
rect 128412 431888 128636 431916
rect 128412 431876 128418 431888
rect 128630 431876 128636 431888
rect 128688 431876 128694 431928
rect 265802 429836 265808 429888
rect 265860 429876 265866 429888
rect 266078 429876 266084 429888
rect 265860 429848 266084 429876
rect 265860 429836 265866 429848
rect 266078 429836 266084 429848
rect 266136 429836 266142 429888
rect 271506 429836 271512 429888
rect 271564 429876 271570 429888
rect 271782 429876 271788 429888
rect 271564 429848 271788 429876
rect 271564 429836 271570 429848
rect 271782 429836 271788 429848
rect 271840 429836 271846 429888
rect 301866 429156 301872 429208
rect 301924 429196 301930 429208
rect 302050 429196 302056 429208
rect 301924 429168 302056 429196
rect 301924 429156 301930 429168
rect 302050 429156 302056 429168
rect 302108 429156 302114 429208
rect 281258 427864 281264 427916
rect 281316 427864 281322 427916
rect 8110 427796 8116 427848
rect 8168 427796 8174 427848
rect 8128 427768 8156 427796
rect 281276 427780 281304 427864
rect 302142 427836 302148 427848
rect 302068 427808 302148 427836
rect 302068 427780 302096 427808
rect 302142 427796 302148 427808
rect 302200 427796 302206 427848
rect 8202 427768 8208 427780
rect 8128 427740 8208 427768
rect 8202 427728 8208 427740
rect 8260 427728 8266 427780
rect 281258 427728 281264 427780
rect 281316 427728 281322 427780
rect 302050 427728 302056 427780
rect 302108 427728 302114 427780
rect 265802 425144 265808 425196
rect 265860 425184 265866 425196
rect 265986 425184 265992 425196
rect 265860 425156 265992 425184
rect 265860 425144 265866 425156
rect 265986 425144 265992 425156
rect 266044 425144 266050 425196
rect 271506 425144 271512 425196
rect 271564 425184 271570 425196
rect 271690 425184 271696 425196
rect 271564 425156 271696 425184
rect 271564 425144 271570 425156
rect 271690 425144 271696 425156
rect 271748 425144 271754 425196
rect 7926 425008 7932 425060
rect 7984 425048 7990 425060
rect 8202 425048 8208 425060
rect 7984 425020 8208 425048
rect 7984 425008 7990 425020
rect 8202 425008 8208 425020
rect 8260 425008 8266 425060
rect 265986 425008 265992 425060
rect 266044 425048 266050 425060
rect 266170 425048 266176 425060
rect 266044 425020 266176 425048
rect 266044 425008 266050 425020
rect 266170 425008 266176 425020
rect 266228 425008 266234 425060
rect 271690 425008 271696 425060
rect 271748 425048 271754 425060
rect 271782 425048 271788 425060
rect 271748 425020 271788 425048
rect 271748 425008 271754 425020
rect 271782 425008 271788 425020
rect 271840 425008 271846 425060
rect 308766 423648 308772 423700
rect 308824 423688 308830 423700
rect 308858 423688 308864 423700
rect 308824 423660 308864 423688
rect 308824 423648 308830 423660
rect 308858 423648 308864 423660
rect 308916 423648 308922 423700
rect 281258 423580 281264 423632
rect 281316 423620 281322 423632
rect 281534 423620 281540 423632
rect 281316 423592 281540 423620
rect 281316 423580 281322 423592
rect 281534 423580 281540 423592
rect 281592 423580 281598 423632
rect 128354 422356 128360 422408
rect 128412 422396 128418 422408
rect 128630 422396 128636 422408
rect 128412 422368 128636 422396
rect 128412 422356 128418 422368
rect 128630 422356 128636 422368
rect 128688 422356 128694 422408
rect 302050 418140 302056 418192
rect 302108 418140 302114 418192
rect 302068 418056 302096 418140
rect 302050 418004 302056 418056
rect 302108 418004 302114 418056
rect 7926 415420 7932 415472
rect 7984 415460 7990 415472
rect 8110 415460 8116 415472
rect 7984 415432 8116 415460
rect 7984 415420 7990 415432
rect 8110 415420 8116 415432
rect 8168 415420 8174 415472
rect 132954 415420 132960 415472
rect 133012 415460 133018 415472
rect 579798 415460 579804 415472
rect 133012 415432 579804 415460
rect 133012 415420 133018 415432
rect 579798 415420 579804 415432
rect 579856 415420 579862 415472
rect 281626 413924 281632 413976
rect 281684 413964 281690 413976
rect 281810 413964 281816 413976
rect 281684 413936 281816 413964
rect 281684 413924 281690 413936
rect 281810 413924 281816 413936
rect 281868 413924 281874 413976
rect 265710 411136 265716 411188
rect 265768 411176 265774 411188
rect 265894 411176 265900 411188
rect 265768 411148 265900 411176
rect 265768 411136 265774 411148
rect 265894 411136 265900 411148
rect 265952 411136 265958 411188
rect 254578 411068 254584 411120
rect 254636 411108 254642 411120
rect 269574 411108 269580 411120
rect 254636 411080 269580 411108
rect 254636 411068 254642 411080
rect 269574 411068 269580 411080
rect 269632 411068 269638 411120
rect 254670 411000 254676 411052
rect 254728 411040 254734 411052
rect 266354 411040 266360 411052
rect 254728 411012 266360 411040
rect 254728 411000 254734 411012
rect 266354 411000 266360 411012
rect 266412 411000 266418 411052
rect 258718 410932 258724 410984
rect 258776 410972 258782 410984
rect 266998 410972 267004 410984
rect 258776 410944 267004 410972
rect 258776 410932 258782 410944
rect 266998 410932 267004 410944
rect 267056 410932 267062 410984
rect 226150 410864 226156 410916
rect 226208 410904 226214 410916
rect 270770 410904 270776 410916
rect 226208 410876 270776 410904
rect 226208 410864 226214 410876
rect 270770 410864 270776 410876
rect 270828 410864 270834 410916
rect 223390 410796 223396 410848
rect 223448 410836 223454 410848
rect 266538 410836 266544 410848
rect 223448 410808 266544 410836
rect 223448 410796 223454 410808
rect 266538 410796 266544 410808
rect 266596 410796 266602 410848
rect 246022 410728 246028 410780
rect 246080 410768 246086 410780
rect 270678 410768 270684 410780
rect 246080 410740 270684 410768
rect 246080 410728 246086 410740
rect 270678 410728 270684 410740
rect 270736 410728 270742 410780
rect 211982 410660 211988 410712
rect 212040 410700 212046 410712
rect 258718 410700 258724 410712
rect 212040 410672 258724 410700
rect 212040 410660 212046 410672
rect 258718 410660 258724 410672
rect 258776 410660 258782 410712
rect 258810 410660 258816 410712
rect 258868 410700 258874 410712
rect 266722 410700 266728 410712
rect 258868 410672 266728 410700
rect 258868 410660 258874 410672
rect 266722 410660 266728 410672
rect 266780 410660 266786 410712
rect 206278 410592 206284 410644
rect 206336 410632 206342 410644
rect 270494 410632 270500 410644
rect 206336 410604 270500 410632
rect 206336 410592 206342 410604
rect 270494 410592 270500 410604
rect 270552 410592 270558 410644
rect 203334 410524 203340 410576
rect 203392 410564 203398 410576
rect 254578 410564 254584 410576
rect 203392 410536 254584 410564
rect 203392 410524 203398 410536
rect 254578 410524 254584 410536
rect 254636 410524 254642 410576
rect 257246 410524 257252 410576
rect 257304 410564 257310 410576
rect 269206 410564 269212 410576
rect 257304 410536 269212 410564
rect 257304 410524 257310 410536
rect 269206 410524 269212 410536
rect 269264 410524 269270 410576
rect 240318 410456 240324 410508
rect 240376 410496 240382 410508
rect 266446 410496 266452 410508
rect 240376 410468 266452 410496
rect 240376 410456 240382 410468
rect 266446 410456 266452 410468
rect 266504 410456 266510 410508
rect 237558 410388 237564 410440
rect 237616 410428 237622 410440
rect 258810 410428 258816 410440
rect 237616 410400 258816 410428
rect 237616 410388 237622 410400
rect 258810 410388 258816 410400
rect 258868 410388 258874 410440
rect 260374 410388 260380 410440
rect 260432 410428 260438 410440
rect 267274 410428 267280 410440
rect 260432 410400 267280 410428
rect 260432 410388 260438 410400
rect 267274 410388 267280 410400
rect 267332 410388 267338 410440
rect 234614 410320 234620 410372
rect 234672 410360 234678 410372
rect 257246 410360 257252 410372
rect 234672 410332 257252 410360
rect 234672 410320 234678 410332
rect 257246 410320 257252 410332
rect 257304 410320 257310 410372
rect 257338 410320 257344 410372
rect 257396 410360 257402 410372
rect 269298 410360 269304 410372
rect 257396 410332 269304 410360
rect 257396 410320 257402 410332
rect 269298 410320 269304 410332
rect 269356 410320 269362 410372
rect 231854 410252 231860 410304
rect 231912 410292 231918 410304
rect 270862 410292 270868 410304
rect 231912 410264 270868 410292
rect 231912 410252 231918 410264
rect 270862 410252 270868 410264
rect 270920 410252 270926 410304
rect 228910 410184 228916 410236
rect 228968 410224 228974 410236
rect 270586 410224 270592 410236
rect 228968 410196 270592 410224
rect 228968 410184 228974 410196
rect 270586 410184 270592 410196
rect 270644 410184 270650 410236
rect 200022 410116 200028 410168
rect 200080 410156 200086 410168
rect 217686 410156 217692 410168
rect 200080 410128 217692 410156
rect 200080 410116 200086 410128
rect 217686 410116 217692 410128
rect 217744 410116 217750 410168
rect 251726 410116 251732 410168
rect 251784 410156 251790 410168
rect 257338 410156 257344 410168
rect 251784 410128 257344 410156
rect 251784 410116 251790 410128
rect 257338 410116 257344 410128
rect 257396 410116 257402 410168
rect 257430 410116 257436 410168
rect 257488 410156 257494 410168
rect 269390 410156 269396 410168
rect 257488 410128 269396 410156
rect 257488 410116 257494 410128
rect 269390 410116 269396 410128
rect 269448 410116 269454 410168
rect 195514 410048 195520 410100
rect 195572 410088 195578 410100
rect 220446 410088 220452 410100
rect 195572 410060 220452 410088
rect 195572 410048 195578 410060
rect 220446 410048 220452 410060
rect 220504 410048 220510 410100
rect 269482 410088 269488 410100
rect 258644 410060 269488 410088
rect 195606 409980 195612 410032
rect 195664 410020 195670 410032
rect 214742 410020 214748 410032
rect 195664 409992 214748 410020
rect 195664 409980 195670 409992
rect 214742 409980 214748 409992
rect 214800 409980 214806 410032
rect 248966 409980 248972 410032
rect 249024 410020 249030 410032
rect 258644 410020 258672 410060
rect 269482 410048 269488 410060
rect 269540 410048 269546 410100
rect 266630 410020 266636 410032
rect 249024 409992 258672 410020
rect 258736 409992 266636 410020
rect 249024 409980 249030 409992
rect 199930 409912 199936 409964
rect 199988 409952 199994 409964
rect 209038 409952 209044 409964
rect 199988 409924 209044 409952
rect 199988 409912 199994 409924
rect 209038 409912 209044 409924
rect 209096 409912 209102 409964
rect 243262 409912 243268 409964
rect 243320 409952 243326 409964
rect 258736 409952 258764 409992
rect 266630 409980 266636 409992
rect 266688 409980 266694 410032
rect 243320 409924 258764 409952
rect 243320 409912 243326 409924
rect 263134 409912 263140 409964
rect 263192 409952 263198 409964
rect 267366 409952 267372 409964
rect 263192 409924 267372 409952
rect 263192 409912 263198 409924
rect 267366 409912 267372 409924
rect 267424 409912 267430 409964
rect 196986 409844 196992 409896
rect 197044 409884 197050 409896
rect 200574 409884 200580 409896
rect 197044 409856 200580 409884
rect 197044 409844 197050 409856
rect 200574 409844 200580 409856
rect 200632 409844 200638 409896
rect 265894 409844 265900 409896
rect 265952 409884 265958 409896
rect 268746 409884 268752 409896
rect 265952 409856 268752 409884
rect 265952 409844 265958 409856
rect 268746 409844 268752 409856
rect 268804 409844 268810 409896
rect 196802 409640 196808 409692
rect 196860 409680 196866 409692
rect 202874 409680 202880 409692
rect 196860 409652 202880 409680
rect 196860 409640 196866 409652
rect 202874 409640 202880 409652
rect 202932 409640 202938 409692
rect 196894 409572 196900 409624
rect 196952 409612 196958 409624
rect 205634 409612 205640 409624
rect 196952 409584 205640 409612
rect 196952 409572 196958 409584
rect 205634 409572 205640 409584
rect 205692 409572 205698 409624
rect 195422 409504 195428 409556
rect 195480 409544 195486 409556
rect 209774 409544 209780 409556
rect 195480 409516 209780 409544
rect 195480 409504 195486 409516
rect 209774 409504 209780 409516
rect 209832 409504 209838 409556
rect 195146 409436 195152 409488
rect 195204 409476 195210 409488
rect 212534 409476 212540 409488
rect 195204 409448 212540 409476
rect 195204 409436 195210 409448
rect 212534 409436 212540 409448
rect 212592 409436 212598 409488
rect 196618 409368 196624 409420
rect 196676 409408 196682 409420
rect 215294 409408 215300 409420
rect 196676 409380 215300 409408
rect 196676 409368 196682 409380
rect 215294 409368 215300 409380
rect 215352 409368 215358 409420
rect 196710 409300 196716 409352
rect 196768 409340 196774 409352
rect 219434 409340 219440 409352
rect 196768 409312 219440 409340
rect 196768 409300 196774 409312
rect 219434 409300 219440 409312
rect 219492 409300 219498 409352
rect 195330 409232 195336 409284
rect 195388 409272 195394 409284
rect 219526 409272 219532 409284
rect 195388 409244 219532 409272
rect 195388 409232 195394 409244
rect 219526 409232 219532 409244
rect 219584 409232 219590 409284
rect 196526 409164 196532 409216
rect 196584 409204 196590 409216
rect 222194 409204 222200 409216
rect 196584 409176 222200 409204
rect 196584 409164 196590 409176
rect 222194 409164 222200 409176
rect 222252 409164 222258 409216
rect 195238 409096 195244 409148
rect 195296 409136 195302 409148
rect 222286 409136 222292 409148
rect 195296 409108 222292 409136
rect 195296 409096 195302 409108
rect 222286 409096 222292 409108
rect 222344 409096 222350 409148
rect 8110 408484 8116 408536
rect 8168 408484 8174 408536
rect 271598 408484 271604 408536
rect 271656 408524 271662 408536
rect 271966 408524 271972 408536
rect 271656 408496 271972 408524
rect 271656 408484 271662 408496
rect 271966 408484 271972 408496
rect 272024 408484 272030 408536
rect 8128 408388 8156 408484
rect 8202 408388 8208 408400
rect 8128 408360 8208 408388
rect 8202 408348 8208 408360
rect 8260 408348 8266 408400
rect 265710 408348 265716 408400
rect 265768 408388 265774 408400
rect 266078 408388 266084 408400
rect 265768 408360 266084 408388
rect 265768 408348 265774 408360
rect 266078 408348 266084 408360
rect 266136 408348 266142 408400
rect 188338 407804 188344 407856
rect 188396 407844 188402 407856
rect 380526 407844 380532 407856
rect 188396 407816 380532 407844
rect 188396 407804 188402 407816
rect 380526 407804 380532 407816
rect 380584 407804 380590 407856
rect 70118 407736 70124 407788
rect 70176 407776 70182 407788
rect 104802 407776 104808 407788
rect 70176 407748 104808 407776
rect 70176 407736 70182 407748
rect 104802 407736 104808 407748
rect 104860 407776 104866 407788
rect 416774 407776 416780 407788
rect 104860 407748 416780 407776
rect 104860 407736 104866 407748
rect 416774 407736 416780 407748
rect 416832 407736 416838 407788
rect 155218 407600 155224 407652
rect 155276 407640 155282 407652
rect 155862 407640 155868 407652
rect 155276 407612 155868 407640
rect 155276 407600 155282 407612
rect 155862 407600 155868 407612
rect 155920 407600 155926 407652
rect 155862 407192 155868 407244
rect 155920 407232 155926 407244
rect 416866 407232 416872 407244
rect 155920 407204 416872 407232
rect 155920 407192 155926 407204
rect 416866 407192 416872 407204
rect 416924 407192 416930 407244
rect 127802 407124 127808 407176
rect 127860 407164 127866 407176
rect 411254 407164 411260 407176
rect 127860 407136 411260 407164
rect 127860 407124 127866 407136
rect 411254 407124 411260 407136
rect 411312 407124 411318 407176
rect 197722 406512 197728 406564
rect 197780 406552 197786 406564
rect 293954 406552 293960 406564
rect 197780 406524 293960 406552
rect 197780 406512 197786 406524
rect 293954 406512 293960 406524
rect 294012 406512 294018 406564
rect 199378 406444 199384 406496
rect 199436 406484 199442 406496
rect 402974 406484 402980 406496
rect 199436 406456 402980 406484
rect 199436 406444 199442 406456
rect 402974 406444 402980 406456
rect 403032 406444 403038 406496
rect 293954 406376 293960 406428
rect 294012 406416 294018 406428
rect 294598 406416 294604 406428
rect 294012 406388 294604 406416
rect 294012 406376 294018 406388
rect 294598 406376 294604 406388
rect 294656 406376 294662 406428
rect 308766 404336 308772 404388
rect 308824 404376 308830 404388
rect 308858 404376 308864 404388
rect 308824 404348 308864 404376
rect 308824 404336 308830 404348
rect 308858 404336 308864 404348
rect 308916 404336 308922 404388
rect 301774 401616 301780 401668
rect 301832 401656 301838 401668
rect 302050 401656 302056 401668
rect 301832 401628 302056 401656
rect 301832 401616 301838 401628
rect 302050 401616 302056 401628
rect 302108 401616 302114 401668
rect 8202 400868 8208 400920
rect 8260 400908 8266 400920
rect 8386 400908 8392 400920
rect 8260 400880 8392 400908
rect 8260 400868 8266 400880
rect 8386 400868 8392 400880
rect 8444 400868 8450 400920
rect 120902 398896 120908 398948
rect 120960 398936 120966 398948
rect 121362 398936 121368 398948
rect 120960 398908 121368 398936
rect 120960 398896 120966 398908
rect 121362 398896 121368 398908
rect 121420 398936 121426 398948
rect 125686 398936 125692 398948
rect 121420 398908 125692 398936
rect 121420 398896 121426 398908
rect 125686 398896 125692 398908
rect 125744 398896 125750 398948
rect 71682 398828 71688 398880
rect 71740 398868 71746 398880
rect 85482 398868 85488 398880
rect 71740 398840 85488 398868
rect 71740 398828 71746 398840
rect 85482 398828 85488 398840
rect 85540 398828 85546 398880
rect 110966 398828 110972 398880
rect 111024 398868 111030 398880
rect 111702 398868 111708 398880
rect 111024 398840 111708 398868
rect 111024 398828 111030 398840
rect 111702 398828 111708 398840
rect 111760 398868 111766 398880
rect 126054 398868 126060 398880
rect 111760 398840 126060 398868
rect 111760 398828 111766 398840
rect 126054 398828 126060 398840
rect 126112 398828 126118 398880
rect 113542 398760 113548 398812
rect 113600 398800 113606 398812
rect 113818 398800 113824 398812
rect 113600 398772 113824 398800
rect 113600 398760 113606 398772
rect 113818 398760 113824 398772
rect 113876 398800 113882 398812
rect 126974 398800 126980 398812
rect 113876 398772 126980 398800
rect 113876 398760 113882 398772
rect 126974 398760 126980 398772
rect 127032 398800 127038 398812
rect 127802 398800 127808 398812
rect 127032 398772 127808 398800
rect 127032 398760 127038 398772
rect 127802 398760 127808 398772
rect 127860 398760 127866 398812
rect 271598 398760 271604 398812
rect 271656 398800 271662 398812
rect 271782 398800 271788 398812
rect 271656 398772 271788 398800
rect 271656 398760 271662 398772
rect 271782 398760 271788 398772
rect 271840 398760 271846 398812
rect 85482 398692 85488 398744
rect 85540 398732 85546 398744
rect 90266 398732 90272 398744
rect 85540 398704 90272 398732
rect 85540 398692 85546 398704
rect 90266 398692 90272 398704
rect 90324 398692 90330 398744
rect 125594 398216 125600 398268
rect 125652 398256 125658 398268
rect 128262 398256 128268 398268
rect 125652 398228 128268 398256
rect 125652 398216 125658 398228
rect 128262 398216 128268 398228
rect 128320 398256 128326 398268
rect 138014 398256 138020 398268
rect 128320 398228 138020 398256
rect 128320 398216 128326 398228
rect 138014 398216 138020 398228
rect 138072 398216 138078 398268
rect 100662 398148 100668 398200
rect 100720 398188 100726 398200
rect 113542 398188 113548 398200
rect 100720 398160 113548 398188
rect 100720 398148 100726 398160
rect 113542 398148 113548 398160
rect 113600 398148 113606 398200
rect 75822 398080 75828 398132
rect 75880 398120 75886 398132
rect 115934 398120 115940 398132
rect 75880 398092 115940 398120
rect 75880 398080 75886 398092
rect 115934 398080 115940 398092
rect 115992 398120 115998 398132
rect 127250 398120 127256 398132
rect 115992 398092 127256 398120
rect 115992 398080 115998 398092
rect 127250 398080 127256 398092
rect 127308 398080 127314 398132
rect 128262 398080 128268 398132
rect 128320 398120 128326 398132
rect 155218 398120 155224 398132
rect 128320 398092 155224 398120
rect 128320 398080 128326 398092
rect 155218 398080 155224 398092
rect 155276 398080 155282 398132
rect 80790 397740 80796 397792
rect 80848 397780 80854 397792
rect 124122 397780 124128 397792
rect 80848 397752 124128 397780
rect 80848 397740 80854 397752
rect 124122 397740 124128 397752
rect 124180 397740 124186 397792
rect 105998 397672 106004 397724
rect 106056 397712 106062 397724
rect 130102 397712 130108 397724
rect 106056 397684 130108 397712
rect 106056 397672 106062 397684
rect 130102 397672 130108 397684
rect 130160 397672 130166 397724
rect 95878 397604 95884 397656
rect 95936 397644 95942 397656
rect 126238 397644 126244 397656
rect 95936 397616 126244 397644
rect 95936 397604 95942 397616
rect 126238 397604 126244 397616
rect 126296 397604 126302 397656
rect 85942 397536 85948 397588
rect 86000 397576 86006 397588
rect 128262 397576 128268 397588
rect 86000 397548 128268 397576
rect 86000 397536 86006 397548
rect 128262 397536 128268 397548
rect 128320 397536 128326 397588
rect 115842 397468 115848 397520
rect 115900 397508 115906 397520
rect 127618 397508 127624 397520
rect 115900 397480 127624 397508
rect 115900 397468 115906 397480
rect 127618 397468 127624 397480
rect 127676 397468 127682 397520
rect 124122 397400 124128 397452
rect 124180 397440 124186 397452
rect 124858 397440 124864 397452
rect 124180 397412 124864 397440
rect 124180 397400 124186 397412
rect 124858 397400 124864 397412
rect 124916 397440 124922 397452
rect 125778 397440 125784 397452
rect 124916 397412 125784 397440
rect 124916 397400 124922 397412
rect 125778 397400 125784 397412
rect 125836 397400 125842 397452
rect 71498 396720 71504 396772
rect 71556 396760 71562 396772
rect 117958 396760 117964 396772
rect 71556 396732 117964 396760
rect 71556 396720 71562 396732
rect 117958 396720 117964 396732
rect 118016 396760 118022 396772
rect 126330 396760 126336 396772
rect 118016 396732 126336 396760
rect 118016 396720 118022 396732
rect 126330 396720 126336 396732
rect 126388 396720 126394 396772
rect 8018 396040 8024 396092
rect 8076 396080 8082 396092
rect 8386 396080 8392 396092
rect 8076 396052 8392 396080
rect 8076 396040 8082 396052
rect 8386 396040 8392 396052
rect 8444 396040 8450 396092
rect 83918 395972 83924 396024
rect 83976 396012 83982 396024
rect 84562 396012 84568 396024
rect 83976 395984 84568 396012
rect 83976 395972 83982 395984
rect 84562 395972 84568 395984
rect 84620 395972 84626 396024
rect 96614 395876 96620 395888
rect 83752 395848 96620 395876
rect 71590 395700 71596 395752
rect 71648 395740 71654 395752
rect 83752 395740 83780 395848
rect 96614 395836 96620 395848
rect 96672 395836 96678 395888
rect 84102 395740 84108 395752
rect 71648 395712 83780 395740
rect 83936 395712 84108 395740
rect 71648 395700 71654 395712
rect 83734 395632 83740 395684
rect 83792 395632 83798 395684
rect 72326 395496 72332 395548
rect 72384 395536 72390 395548
rect 83752 395536 83780 395632
rect 72384 395508 83780 395536
rect 83936 395536 83964 395712
rect 84102 395700 84108 395712
rect 84160 395700 84166 395752
rect 84562 395700 84568 395752
rect 84620 395740 84626 395752
rect 84620 395712 99236 395740
rect 84620 395700 84626 395712
rect 84010 395632 84016 395684
rect 84068 395632 84074 395684
rect 99208 395672 99236 395712
rect 99282 395700 99288 395752
rect 99340 395740 99346 395752
rect 108942 395740 108948 395752
rect 99340 395712 108948 395740
rect 99340 395700 99346 395712
rect 108942 395700 108948 395712
rect 109000 395740 109006 395752
rect 125870 395740 125876 395752
rect 109000 395712 125876 395740
rect 109000 395700 109006 395712
rect 125870 395700 125876 395712
rect 125928 395700 125934 395752
rect 126882 395672 126888 395684
rect 99208 395644 126888 395672
rect 126882 395632 126888 395644
rect 126940 395632 126946 395684
rect 84028 395604 84056 395632
rect 168650 395604 168656 395616
rect 84028 395576 168656 395604
rect 168650 395564 168656 395576
rect 168708 395564 168714 395616
rect 179506 395536 179512 395548
rect 83936 395508 179512 395536
rect 72384 395496 72390 395508
rect 179506 395496 179512 395508
rect 179564 395496 179570 395548
rect 8018 394680 8024 394732
rect 8076 394720 8082 394732
rect 8110 394720 8116 394732
rect 8076 394692 8116 394720
rect 8076 394680 8082 394692
rect 8110 394680 8116 394692
rect 8168 394680 8174 394732
rect 308582 394544 308588 394596
rect 308640 394584 308646 394596
rect 308858 394584 308864 394596
rect 308640 394556 308864 394584
rect 308640 394544 308646 394556
rect 308858 394544 308864 394556
rect 308916 394544 308922 394596
rect 128354 393252 128360 393304
rect 128412 393292 128418 393304
rect 128630 393292 128636 393304
rect 128412 393264 128636 393292
rect 128412 393252 128418 393264
rect 128630 393252 128636 393264
rect 128688 393252 128694 393304
rect 402974 393252 402980 393304
rect 403032 393292 403038 393304
rect 403894 393292 403900 393304
rect 403032 393264 403900 393292
rect 403032 393252 403038 393264
rect 403894 393252 403900 393264
rect 403952 393252 403958 393304
rect 266170 392572 266176 392624
rect 266228 392612 266234 392624
rect 436186 392612 436192 392624
rect 266228 392584 436192 392612
rect 266228 392572 266234 392584
rect 436186 392572 436192 392584
rect 436244 392572 436250 392624
rect 301866 391960 301872 392012
rect 301924 392000 301930 392012
rect 302050 392000 302056 392012
rect 301924 391972 302056 392000
rect 301924 391960 301930 391972
rect 302050 391960 302056 391972
rect 302108 391960 302114 392012
rect 126882 391892 126888 391944
rect 126940 391932 126946 391944
rect 199378 391932 199384 391944
rect 126940 391904 199384 391932
rect 126940 391892 126946 391904
rect 199378 391892 199384 391904
rect 199436 391892 199442 391944
rect 458818 389376 458824 389428
rect 458876 389416 458882 389428
rect 475838 389416 475844 389428
rect 458876 389388 475844 389416
rect 458876 389376 458882 389388
rect 475838 389376 475844 389388
rect 475896 389376 475902 389428
rect 416682 389308 416688 389360
rect 416740 389348 416746 389360
rect 464246 389348 464252 389360
rect 416740 389320 464252 389348
rect 416740 389308 416746 389320
rect 464246 389308 464252 389320
rect 464304 389308 464310 389360
rect 418062 389240 418068 389292
rect 418120 389280 418126 389292
rect 487430 389280 487436 389292
rect 418120 389252 487436 389280
rect 418120 389240 418126 389252
rect 487430 389240 487436 389252
rect 487488 389240 487494 389292
rect 8110 389172 8116 389224
rect 8168 389172 8174 389224
rect 416590 389172 416596 389224
rect 416648 389212 416654 389224
rect 499022 389212 499028 389224
rect 416648 389184 499028 389212
rect 416648 389172 416654 389184
rect 499022 389172 499028 389184
rect 499080 389172 499086 389224
rect 8128 389076 8156 389172
rect 271506 389104 271512 389156
rect 271564 389144 271570 389156
rect 271598 389144 271604 389156
rect 271564 389116 271604 389144
rect 271564 389104 271570 389116
rect 271598 389104 271604 389116
rect 271656 389104 271662 389156
rect 297174 389104 297180 389156
rect 297232 389144 297238 389156
rect 298002 389144 298008 389156
rect 297232 389116 298008 389144
rect 297232 389104 297238 389116
rect 298002 389104 298008 389116
rect 298060 389104 298066 389156
rect 8202 389076 8208 389088
rect 8128 389048 8208 389076
rect 8202 389036 8208 389048
rect 8260 389036 8266 389088
rect 126882 386316 126888 386368
rect 126940 386356 126946 386368
rect 130378 386356 130384 386368
rect 126940 386328 130384 386356
rect 126940 386316 126946 386328
rect 130378 386316 130384 386328
rect 130436 386316 130442 386368
rect 281350 386316 281356 386368
rect 281408 386356 281414 386368
rect 281534 386356 281540 386368
rect 281408 386328 281540 386356
rect 281408 386316 281414 386328
rect 281534 386316 281540 386328
rect 281592 386316 281598 386368
rect 306834 386316 306840 386368
rect 306892 386356 306898 386368
rect 307018 386356 307024 386368
rect 306892 386328 307024 386356
rect 306892 386316 306898 386328
rect 307018 386316 307024 386328
rect 307076 386316 307082 386368
rect 344922 385704 344928 385756
rect 344980 385744 344986 385756
rect 408862 385744 408868 385756
rect 344980 385716 408868 385744
rect 344980 385704 344986 385716
rect 408862 385704 408868 385716
rect 408920 385704 408926 385756
rect 294598 385636 294604 385688
rect 294656 385676 294662 385688
rect 388254 385676 388260 385688
rect 294656 385648 388260 385676
rect 294656 385636 294662 385648
rect 388254 385636 388260 385648
rect 388312 385636 388318 385688
rect 365622 385568 365628 385620
rect 365680 385608 365686 385620
rect 392854 385608 392860 385620
rect 365680 385580 392860 385608
rect 365680 385568 365686 385580
rect 392854 385568 392860 385580
rect 392912 385568 392918 385620
rect 349062 385500 349068 385552
rect 349120 385540 349126 385552
rect 385862 385540 385868 385552
rect 349120 385512 385868 385540
rect 349120 385500 349126 385512
rect 385862 385500 385868 385512
rect 385920 385500 385926 385552
rect 355870 385432 355876 385484
rect 355928 385472 355934 385484
rect 399662 385472 399668 385484
rect 355928 385444 399668 385472
rect 355928 385432 355934 385444
rect 399662 385432 399668 385444
rect 399720 385432 399726 385484
rect 353202 385364 353208 385416
rect 353260 385404 353266 385416
rect 402054 385404 402060 385416
rect 353260 385376 402060 385404
rect 353260 385364 353266 385376
rect 402054 385364 402060 385376
rect 402112 385364 402118 385416
rect 357342 385296 357348 385348
rect 357400 385336 357406 385348
rect 406654 385336 406660 385348
rect 357400 385308 406660 385336
rect 357400 385296 357406 385308
rect 406654 385296 406660 385308
rect 406712 385296 406718 385348
rect 347682 385228 347688 385280
rect 347740 385268 347746 385280
rect 397454 385268 397460 385280
rect 347740 385240 397460 385268
rect 347740 385228 347746 385240
rect 397454 385228 397460 385240
rect 397512 385228 397518 385280
rect 343542 385160 343548 385212
rect 343600 385200 343606 385212
rect 395062 385200 395068 385212
rect 343600 385172 395068 385200
rect 343600 385160 343606 385172
rect 395062 385160 395068 385172
rect 395120 385160 395126 385212
rect 355962 385092 355968 385144
rect 356020 385132 356026 385144
rect 413462 385132 413468 385144
rect 356020 385104 413468 385132
rect 356020 385092 356026 385104
rect 413462 385092 413468 385104
rect 413520 385092 413526 385144
rect 367002 385024 367008 385076
rect 367060 385064 367066 385076
rect 390462 385064 390468 385076
rect 367060 385036 390468 385064
rect 367060 385024 367066 385036
rect 390462 385024 390468 385036
rect 390520 385024 390526 385076
rect 126330 384956 126336 385008
rect 126388 384996 126394 385008
rect 130286 384996 130292 385008
rect 126388 384968 130292 384996
rect 126388 384956 126394 384968
rect 130286 384956 130292 384968
rect 130344 384956 130350 385008
rect 271506 384208 271512 384260
rect 271564 384248 271570 384260
rect 271690 384248 271696 384260
rect 271564 384220 271696 384248
rect 271564 384208 271570 384220
rect 271690 384208 271696 384220
rect 271748 384208 271754 384260
rect 128354 383664 128360 383716
rect 128412 383704 128418 383716
rect 128630 383704 128636 383716
rect 128412 383676 128636 383704
rect 128412 383664 128418 383676
rect 128630 383664 128636 383676
rect 128688 383664 128694 383716
rect 301498 381488 301504 381540
rect 301556 381528 301562 381540
rect 301958 381528 301964 381540
rect 301556 381500 301964 381528
rect 301556 381488 301562 381500
rect 301958 381488 301964 381500
rect 302016 381528 302022 381540
rect 380894 381528 380900 381540
rect 302016 381500 380900 381528
rect 302016 381488 302022 381500
rect 380894 381488 380900 381500
rect 380952 381488 380958 381540
rect 8202 379556 8208 379568
rect 8036 379528 8208 379556
rect 8036 379500 8064 379528
rect 8202 379516 8208 379528
rect 8260 379516 8266 379568
rect 297174 379516 297180 379568
rect 297232 379556 297238 379568
rect 298002 379556 298008 379568
rect 297232 379528 298008 379556
rect 297232 379516 297238 379528
rect 298002 379516 298008 379528
rect 298060 379516 298066 379568
rect 8018 379448 8024 379500
rect 8076 379448 8082 379500
rect 271690 379448 271696 379500
rect 271748 379488 271754 379500
rect 271782 379488 271788 379500
rect 271748 379460 271788 379488
rect 271748 379448 271754 379460
rect 271782 379448 271788 379460
rect 271840 379448 271846 379500
rect 281166 376796 281172 376848
rect 281224 376836 281230 376848
rect 281534 376836 281540 376848
rect 281224 376808 281540 376836
rect 281224 376796 281230 376808
rect 281534 376796 281540 376808
rect 281592 376796 281598 376848
rect 306834 376728 306840 376780
rect 306892 376768 306898 376780
rect 307018 376768 307024 376780
rect 306892 376740 307024 376768
rect 306892 376728 306898 376740
rect 307018 376728 307024 376740
rect 307076 376728 307082 376780
rect 308582 376728 308588 376780
rect 308640 376768 308646 376780
rect 308674 376768 308680 376780
rect 308640 376740 308680 376768
rect 308640 376728 308646 376740
rect 308674 376728 308680 376740
rect 308732 376728 308738 376780
rect 351822 376728 351828 376780
rect 351880 376768 351886 376780
rect 380894 376768 380900 376780
rect 351880 376740 380900 376768
rect 351880 376728 351886 376740
rect 380894 376728 380900 376740
rect 380952 376728 380958 376780
rect 281074 376660 281080 376712
rect 281132 376700 281138 376712
rect 281166 376700 281172 376712
rect 281132 376672 281172 376700
rect 281132 376660 281138 376672
rect 281166 376660 281172 376672
rect 281224 376660 281230 376712
rect 7834 375300 7840 375352
rect 7892 375340 7898 375352
rect 8018 375340 8024 375352
rect 7892 375312 8024 375340
rect 7892 375300 7898 375312
rect 8018 375300 8024 375312
rect 8076 375300 8082 375352
rect 129090 374116 129096 374128
rect 128832 374088 129096 374116
rect 128832 374060 128860 374088
rect 129090 374076 129096 374088
rect 129148 374076 129154 374128
rect 128814 374008 128820 374060
rect 128872 374008 128878 374060
rect 364242 374008 364248 374060
rect 364300 374048 364306 374060
rect 380894 374048 380900 374060
rect 364300 374020 380900 374048
rect 364300 374008 364306 374020
rect 380894 374008 380900 374020
rect 380952 374008 380958 374060
rect 414658 374008 414664 374060
rect 414716 374048 414722 374060
rect 456794 374048 456800 374060
rect 414716 374020 456800 374048
rect 414716 374008 414722 374020
rect 456794 374008 456800 374020
rect 456852 374008 456858 374060
rect 128354 373940 128360 373992
rect 128412 373980 128418 373992
rect 128538 373980 128544 373992
rect 128412 373952 128544 373980
rect 128412 373940 128418 373952
rect 128538 373940 128544 373952
rect 128596 373940 128602 373992
rect 347590 369860 347596 369912
rect 347648 369900 347654 369912
rect 380894 369900 380900 369912
rect 347648 369872 380900 369900
rect 347648 369860 347654 369872
rect 380894 369860 380900 369872
rect 380952 369860 380958 369912
rect 128538 369792 128544 369844
rect 128596 369792 128602 369844
rect 128556 369764 128584 369792
rect 128630 369764 128636 369776
rect 128556 369736 128636 369764
rect 128630 369724 128636 369736
rect 128688 369724 128694 369776
rect 281074 367140 281080 367192
rect 281132 367180 281138 367192
rect 281350 367180 281356 367192
rect 281132 367152 281356 367180
rect 281132 367140 281138 367152
rect 281350 367140 281356 367152
rect 281408 367140 281414 367192
rect 281074 367004 281080 367056
rect 281132 367044 281138 367056
rect 281350 367044 281356 367056
rect 281132 367016 281356 367044
rect 281132 367004 281138 367016
rect 281350 367004 281356 367016
rect 281408 367004 281414 367056
rect 306834 367004 306840 367056
rect 306892 367044 306898 367056
rect 307018 367044 307024 367056
rect 306892 367016 307024 367044
rect 306892 367004 306898 367016
rect 307018 367004 307024 367016
rect 307076 367004 307082 367056
rect 2958 366120 2964 366172
rect 3016 366160 3022 366172
rect 4982 366160 4988 366172
rect 3016 366132 4988 366160
rect 3016 366120 3022 366132
rect 4982 366120 4988 366132
rect 5040 366120 5046 366172
rect 308674 365780 308680 365832
rect 308732 365820 308738 365832
rect 308858 365820 308864 365832
rect 308732 365792 308864 365820
rect 308732 365780 308738 365792
rect 308858 365780 308864 365792
rect 308916 365780 308922 365832
rect 7834 365712 7840 365764
rect 7892 365752 7898 365764
rect 8110 365752 8116 365764
rect 7892 365724 8116 365752
rect 7892 365712 7898 365724
rect 8110 365712 8116 365724
rect 8168 365712 8174 365764
rect 128906 365644 128912 365696
rect 128964 365684 128970 365696
rect 197722 365684 197728 365696
rect 128964 365656 197728 365684
rect 128964 365644 128970 365656
rect 197722 365644 197728 365656
rect 197780 365644 197786 365696
rect 308674 365644 308680 365696
rect 308732 365684 308738 365696
rect 308858 365684 308864 365696
rect 308732 365656 308864 365684
rect 308732 365644 308738 365656
rect 308858 365644 308864 365656
rect 308916 365644 308922 365696
rect 333882 362924 333888 362976
rect 333940 362964 333946 362976
rect 380894 362964 380900 362976
rect 333940 362936 380900 362964
rect 333940 362924 333946 362936
rect 380894 362924 380900 362936
rect 380952 362924 380958 362976
rect 8110 360204 8116 360256
rect 8168 360204 8174 360256
rect 128814 360204 128820 360256
rect 128872 360244 128878 360256
rect 129090 360244 129096 360256
rect 128872 360216 129096 360244
rect 128872 360204 128878 360216
rect 129090 360204 129096 360216
rect 129148 360204 129154 360256
rect 271690 360204 271696 360256
rect 271748 360244 271754 360256
rect 271782 360244 271788 360256
rect 271748 360216 271788 360244
rect 271748 360204 271754 360216
rect 271782 360204 271788 360216
rect 271840 360204 271846 360256
rect 8128 360176 8156 360204
rect 8202 360176 8208 360188
rect 8128 360148 8208 360176
rect 8202 360136 8208 360148
rect 8260 360136 8266 360188
rect 281074 357484 281080 357536
rect 281132 357524 281138 357536
rect 281166 357524 281172 357536
rect 281132 357496 281172 357524
rect 281132 357484 281138 357496
rect 281166 357484 281172 357496
rect 281224 357484 281230 357536
rect 306834 357416 306840 357468
rect 306892 357456 306898 357468
rect 307018 357456 307024 357468
rect 306892 357428 307024 357456
rect 306892 357416 306898 357428
rect 307018 357416 307024 357428
rect 307076 357416 307082 357468
rect 308674 357416 308680 357468
rect 308732 357456 308738 357468
rect 308732 357428 308904 357456
rect 308732 357416 308738 357428
rect 308876 357400 308904 357428
rect 281074 357348 281080 357400
rect 281132 357388 281138 357400
rect 281166 357388 281172 357400
rect 281132 357360 281172 357388
rect 281132 357348 281138 357360
rect 281166 357348 281172 357360
rect 281224 357348 281230 357400
rect 308858 357348 308864 357400
rect 308916 357348 308922 357400
rect 185578 355988 185584 356040
rect 185636 356028 185642 356040
rect 188338 356028 188344 356040
rect 185636 356000 188344 356028
rect 185636 355988 185642 356000
rect 188338 355988 188344 356000
rect 188396 355988 188402 356040
rect 8202 354628 8208 354680
rect 8260 354668 8266 354680
rect 8386 354668 8392 354680
rect 8260 354640 8392 354668
rect 8260 354628 8266 354640
rect 8386 354628 8392 354640
rect 8444 354628 8450 354680
rect 354582 353268 354588 353320
rect 354640 353308 354646 353320
rect 380894 353308 380900 353320
rect 354640 353280 380900 353308
rect 354640 353268 354646 353280
rect 380894 353268 380900 353280
rect 380952 353268 380958 353320
rect 129734 350548 129740 350600
rect 129792 350588 129798 350600
rect 130470 350588 130476 350600
rect 129792 350560 130476 350588
rect 129792 350548 129798 350560
rect 130470 350548 130476 350560
rect 130528 350548 130534 350600
rect 128722 347936 128728 347948
rect 128648 347908 128728 347936
rect 128648 347812 128676 347908
rect 128722 347896 128728 347908
rect 128780 347896 128786 347948
rect 281074 347828 281080 347880
rect 281132 347868 281138 347880
rect 281350 347868 281356 347880
rect 281132 347840 281356 347868
rect 281132 347828 281138 347840
rect 281350 347828 281356 347840
rect 281408 347828 281414 347880
rect 128630 347760 128636 347812
rect 128688 347760 128694 347812
rect 128722 347760 128728 347812
rect 128780 347800 128786 347812
rect 129090 347800 129096 347812
rect 128780 347772 129096 347800
rect 128780 347760 128786 347772
rect 129090 347760 129096 347772
rect 129148 347760 129154 347812
rect 281074 347692 281080 347744
rect 281132 347732 281138 347744
rect 281350 347732 281356 347744
rect 281132 347704 281356 347732
rect 281132 347692 281138 347704
rect 281350 347692 281356 347704
rect 281408 347692 281414 347744
rect 306834 347692 306840 347744
rect 306892 347732 306898 347744
rect 306926 347732 306932 347744
rect 306892 347704 306932 347732
rect 306892 347692 306898 347704
rect 306926 347692 306932 347704
rect 306984 347692 306990 347744
rect 365530 347692 365536 347744
rect 365588 347732 365594 347744
rect 386782 347732 386788 347744
rect 365588 347704 386788 347732
rect 365588 347692 365594 347704
rect 386782 347692 386788 347704
rect 386840 347692 386846 347744
rect 360102 347624 360108 347676
rect 360160 347664 360166 347676
rect 391382 347664 391388 347676
rect 360160 347636 391388 347664
rect 360160 347624 360166 347636
rect 391382 347624 391388 347636
rect 391440 347624 391446 347676
rect 358722 347556 358728 347608
rect 358780 347596 358786 347608
rect 393590 347596 393596 347608
rect 358780 347568 393596 347596
rect 358780 347556 358786 347568
rect 393590 347556 393596 347568
rect 393648 347556 393654 347608
rect 362862 347488 362868 347540
rect 362920 347528 362926 347540
rect 398190 347528 398196 347540
rect 362920 347500 398196 347528
rect 362920 347488 362926 347500
rect 398190 347488 398196 347500
rect 398248 347488 398254 347540
rect 362770 347420 362776 347472
rect 362828 347460 362834 347472
rect 402790 347460 402796 347472
rect 362828 347432 402796 347460
rect 362828 347420 362834 347432
rect 402790 347420 402796 347432
rect 402848 347420 402854 347472
rect 350534 347352 350540 347404
rect 350592 347392 350598 347404
rect 395982 347392 395988 347404
rect 350592 347364 395988 347392
rect 350592 347352 350598 347364
rect 395982 347352 395988 347364
rect 396040 347352 396046 347404
rect 342162 347284 342168 347336
rect 342220 347324 342226 347336
rect 388990 347324 388996 347336
rect 342220 347296 388996 347324
rect 342220 347284 342226 347296
rect 388990 347284 388996 347296
rect 389048 347284 389054 347336
rect 361482 347216 361488 347268
rect 361540 347256 361546 347268
rect 407390 347256 407396 347268
rect 361540 347228 407396 347256
rect 361540 347216 361546 347228
rect 407390 347216 407396 347228
rect 407448 347216 407454 347268
rect 354490 347148 354496 347200
rect 354548 347188 354554 347200
rect 400582 347188 400588 347200
rect 354548 347160 400588 347188
rect 354548 347148 354554 347160
rect 400582 347148 400588 347160
rect 400640 347148 400646 347200
rect 361390 347080 361396 347132
rect 361448 347120 361454 347132
rect 414382 347120 414388 347132
rect 361448 347092 414388 347120
rect 361448 347080 361454 347092
rect 414382 347080 414388 347092
rect 414440 347080 414446 347132
rect 274450 347012 274456 347064
rect 274508 347052 274514 347064
rect 310606 347052 310612 347064
rect 274508 347024 310612 347052
rect 274508 347012 274514 347024
rect 310606 347012 310612 347024
rect 310664 347012 310670 347064
rect 333790 347012 333796 347064
rect 333848 347052 333854 347064
rect 411990 347052 411996 347064
rect 333848 347024 411996 347052
rect 333848 347012 333854 347024
rect 411990 347012 411996 347024
rect 412048 347012 412054 347064
rect 130286 346468 130292 346520
rect 130344 346508 130350 346520
rect 132770 346508 132776 346520
rect 130344 346480 132776 346508
rect 130344 346468 130350 346480
rect 132770 346468 132776 346480
rect 132828 346468 132834 346520
rect 308674 346400 308680 346452
rect 308732 346440 308738 346452
rect 308766 346440 308772 346452
rect 308732 346412 308772 346440
rect 308732 346400 308738 346412
rect 308766 346400 308772 346412
rect 308824 346400 308830 346452
rect 128722 345516 128728 345568
rect 128780 345556 128786 345568
rect 129090 345556 129096 345568
rect 128780 345528 129096 345556
rect 128780 345516 128786 345528
rect 129090 345516 129096 345528
rect 129148 345516 129154 345568
rect 8202 345040 8208 345092
rect 8260 345080 8266 345092
rect 8386 345080 8392 345092
rect 8260 345052 8392 345080
rect 8260 345040 8266 345052
rect 8386 345040 8392 345052
rect 8444 345040 8450 345092
rect 504818 345040 504824 345092
rect 504876 345080 504882 345092
rect 579982 345080 579988 345092
rect 504876 345052 579988 345080
rect 504876 345040 504882 345052
rect 579982 345040 579988 345052
rect 580040 345040 580046 345092
rect 135254 342864 135260 342916
rect 135312 342904 135318 342916
rect 191098 342904 191104 342916
rect 135312 342876 191104 342904
rect 135312 342864 135318 342876
rect 191098 342864 191104 342876
rect 191156 342864 191162 342916
rect 199654 342728 199660 342780
rect 199712 342768 199718 342780
rect 200206 342768 200212 342780
rect 199712 342740 200212 342768
rect 199712 342728 199718 342740
rect 200206 342728 200212 342740
rect 200264 342728 200270 342780
rect 128814 342456 128820 342508
rect 128872 342496 128878 342508
rect 135254 342496 135260 342508
rect 128872 342468 135260 342496
rect 128872 342456 128878 342468
rect 135254 342456 135260 342468
rect 135312 342456 135318 342508
rect 503806 341980 503812 342032
rect 503864 342020 503870 342032
rect 504174 342020 504180 342032
rect 503864 341992 504180 342020
rect 503864 341980 503870 341992
rect 504174 341980 504180 341992
rect 504232 341980 504238 342032
rect 126054 340824 126060 340876
rect 126112 340864 126118 340876
rect 408494 340864 408500 340876
rect 126112 340836 408500 340864
rect 126112 340824 126118 340836
rect 408494 340824 408500 340836
rect 408552 340824 408558 340876
rect 504726 340864 504732 340876
rect 504100 340836 504732 340864
rect 127250 340756 127256 340808
rect 127308 340796 127314 340808
rect 404354 340796 404360 340808
rect 127308 340768 404360 340796
rect 127308 340756 127314 340768
rect 404354 340756 404360 340768
rect 404412 340756 404418 340808
rect 503898 340756 503904 340808
rect 503956 340796 503962 340808
rect 504100 340796 504128 340836
rect 504726 340824 504732 340836
rect 504784 340824 504790 340876
rect 503956 340768 504128 340796
rect 503956 340756 503962 340768
rect 127710 340688 127716 340740
rect 127768 340728 127774 340740
rect 381630 340728 381636 340740
rect 127768 340700 381636 340728
rect 127768 340688 127774 340700
rect 381630 340688 381636 340700
rect 381688 340688 381694 340740
rect 130470 340620 130476 340672
rect 130528 340660 130534 340672
rect 381538 340660 381544 340672
rect 130528 340632 381544 340660
rect 130528 340620 130534 340632
rect 381538 340620 381544 340632
rect 381596 340620 381602 340672
rect 132770 340552 132776 340604
rect 132828 340592 132834 340604
rect 383654 340592 383660 340604
rect 132828 340564 383660 340592
rect 132828 340552 132834 340564
rect 383654 340552 383660 340564
rect 383712 340552 383718 340604
rect 173894 340524 173900 340536
rect 166920 340496 173900 340524
rect 130194 340416 130200 340468
rect 130252 340456 130258 340468
rect 138014 340456 138020 340468
rect 130252 340428 138020 340456
rect 130252 340416 130258 340428
rect 138014 340416 138020 340428
rect 138072 340456 138078 340468
rect 154574 340456 154580 340468
rect 138072 340428 154580 340456
rect 138072 340416 138078 340428
rect 154574 340416 154580 340428
rect 154632 340416 154638 340468
rect 166920 340456 166948 340496
rect 173894 340484 173900 340496
rect 173952 340484 173958 340536
rect 202800 340496 205680 340524
rect 202800 340468 202828 340496
rect 164160 340428 166948 340456
rect 157334 340348 157340 340400
rect 157392 340388 157398 340400
rect 164160 340388 164188 340428
rect 183462 340416 183468 340468
rect 183520 340456 183526 340468
rect 183520 340428 186268 340456
rect 183520 340416 183526 340428
rect 157392 340360 164188 340388
rect 186240 340388 186268 340428
rect 202782 340416 202788 340468
rect 202840 340416 202846 340468
rect 205652 340456 205680 340496
rect 240134 340484 240140 340536
rect 240192 340484 240198 340536
rect 259380 340496 259500 340524
rect 215202 340456 215208 340468
rect 205652 340428 215208 340456
rect 215202 340416 215208 340428
rect 215260 340416 215266 340468
rect 240042 340416 240048 340468
rect 240100 340456 240106 340468
rect 240152 340456 240180 340484
rect 240100 340428 240180 340456
rect 240100 340416 240106 340428
rect 249702 340416 249708 340468
rect 249760 340456 249766 340468
rect 259380 340456 259408 340496
rect 259472 340468 259500 340496
rect 269022 340484 269028 340536
rect 269080 340484 269086 340536
rect 280154 340524 280160 340536
rect 278700 340496 280160 340524
rect 249760 340428 259408 340456
rect 249760 340416 249766 340428
rect 259454 340416 259460 340468
rect 259512 340416 259518 340468
rect 269040 340456 269068 340484
rect 269114 340456 269120 340468
rect 269040 340428 269120 340456
rect 269114 340416 269120 340428
rect 269172 340416 269178 340468
rect 273254 340416 273260 340468
rect 273312 340456 273318 340468
rect 278700 340456 278728 340496
rect 280154 340484 280160 340496
rect 280212 340484 280218 340536
rect 340800 340496 350396 340524
rect 273312 340428 278728 340456
rect 273312 340416 273318 340428
rect 333238 340416 333244 340468
rect 333296 340456 333302 340468
rect 340800 340456 340828 340496
rect 333296 340428 340828 340456
rect 333296 340416 333302 340428
rect 193214 340388 193220 340400
rect 186240 340360 193220 340388
rect 157392 340348 157398 340360
rect 193214 340348 193220 340360
rect 193272 340348 193278 340400
rect 224954 340348 224960 340400
rect 225012 340388 225018 340400
rect 230474 340388 230480 340400
rect 225012 340360 230480 340388
rect 225012 340348 225018 340360
rect 230474 340348 230480 340360
rect 230532 340348 230538 340400
rect 292482 340388 292488 340400
rect 284956 340360 292488 340388
rect 173986 340280 173992 340332
rect 174044 340320 174050 340332
rect 183462 340320 183468 340332
rect 174044 340292 183468 340320
rect 174044 340280 174050 340292
rect 183462 340280 183468 340292
rect 183520 340280 183526 340332
rect 215386 340280 215392 340332
rect 215444 340320 215450 340332
rect 224862 340320 224868 340332
rect 215444 340292 224868 340320
rect 215444 340280 215450 340292
rect 224862 340280 224868 340292
rect 224920 340280 224926 340332
rect 280154 340280 280160 340332
rect 280212 340320 280218 340332
rect 284956 340320 284984 340360
rect 292482 340348 292488 340360
rect 292540 340348 292546 340400
rect 304276 340360 318840 340388
rect 280212 340292 284984 340320
rect 280212 340280 280218 340292
rect 292666 340280 292672 340332
rect 292724 340320 292730 340332
rect 304276 340320 304304 340360
rect 318812 340332 318840 340360
rect 318886 340348 318892 340400
rect 318944 340388 318950 340400
rect 331122 340388 331128 340400
rect 318944 340360 331128 340388
rect 318944 340348 318950 340360
rect 331122 340348 331128 340360
rect 331180 340348 331186 340400
rect 292724 340292 304304 340320
rect 292724 340280 292730 340292
rect 318794 340280 318800 340332
rect 318852 340280 318858 340332
rect 350368 340320 350396 340496
rect 367020 340428 369716 340456
rect 357434 340388 357440 340400
rect 357360 340360 357440 340388
rect 357360 340320 357388 340360
rect 357434 340348 357440 340360
rect 357492 340348 357498 340400
rect 362218 340348 362224 340400
rect 362276 340388 362282 340400
rect 367020 340388 367048 340428
rect 362276 340360 367048 340388
rect 369688 340388 369716 340428
rect 381722 340388 381728 340400
rect 369688 340360 381728 340388
rect 362276 340348 362282 340360
rect 381722 340348 381728 340360
rect 381780 340348 381786 340400
rect 350368 340292 357388 340320
rect 114462 340212 114468 340264
rect 114520 340252 114526 340264
rect 126054 340252 126060 340264
rect 114520 340224 126060 340252
rect 114520 340212 114526 340224
rect 126054 340212 126060 340224
rect 126112 340212 126118 340264
rect 331122 340212 331128 340264
rect 331180 340252 331186 340264
rect 333238 340252 333244 340264
rect 331180 340224 333244 340252
rect 331180 340212 331186 340224
rect 333238 340212 333244 340224
rect 333296 340212 333302 340264
rect 357434 340212 357440 340264
rect 357492 340252 357498 340264
rect 362218 340252 362224 340264
rect 357492 340224 362224 340252
rect 357492 340212 357498 340224
rect 362218 340212 362224 340224
rect 362276 340212 362282 340264
rect 110322 340144 110328 340196
rect 110380 340184 110386 340196
rect 127250 340184 127256 340196
rect 110380 340156 127256 340184
rect 110380 340144 110386 340156
rect 127250 340144 127256 340156
rect 127308 340144 127314 340196
rect 196342 338988 196348 339040
rect 196400 339028 196406 339040
rect 209774 339028 209780 339040
rect 196400 339000 209780 339028
rect 196400 338988 196406 339000
rect 209774 338988 209780 339000
rect 209832 338988 209838 339040
rect 199746 338920 199752 338972
rect 199804 338960 199810 338972
rect 213914 338960 213920 338972
rect 199804 338932 213920 338960
rect 199804 338920 199810 338932
rect 213914 338920 213920 338932
rect 213972 338920 213978 338972
rect 199838 338852 199844 338904
rect 199896 338892 199902 338904
rect 215294 338892 215300 338904
rect 199896 338864 215300 338892
rect 199896 338852 199902 338864
rect 215294 338852 215300 338864
rect 215352 338852 215358 338904
rect 196434 338784 196440 338836
rect 196492 338824 196498 338836
rect 222194 338824 222200 338836
rect 196492 338796 222200 338824
rect 196492 338784 196498 338796
rect 222194 338784 222200 338796
rect 222252 338784 222258 338836
rect 257982 338784 257988 338836
rect 258040 338824 258046 338836
rect 267274 338824 267280 338836
rect 258040 338796 267280 338824
rect 258040 338784 258046 338796
rect 267274 338784 267280 338796
rect 267332 338784 267338 338836
rect 195054 338716 195060 338768
rect 195112 338756 195118 338768
rect 220814 338756 220820 338768
rect 195112 338728 220820 338756
rect 195112 338716 195118 338728
rect 220814 338716 220820 338728
rect 220872 338716 220878 338768
rect 237282 338716 237288 338768
rect 237340 338756 237346 338768
rect 267366 338756 267372 338768
rect 237340 338728 267372 338756
rect 237340 338716 237346 338728
rect 267366 338716 267372 338728
rect 267424 338716 267430 338768
rect 262122 338580 262128 338632
rect 262180 338620 262186 338632
rect 268746 338620 268752 338632
rect 262180 338592 268752 338620
rect 262180 338580 262186 338592
rect 268746 338580 268752 338592
rect 268804 338580 268810 338632
rect 281074 338104 281080 338156
rect 281132 338144 281138 338156
rect 281258 338144 281264 338156
rect 281132 338116 281264 338144
rect 281132 338104 281138 338116
rect 281258 338104 281264 338116
rect 281316 338104 281322 338156
rect 306834 338104 306840 338156
rect 306892 338144 306898 338156
rect 307018 338144 307024 338156
rect 306892 338116 307024 338144
rect 306892 338104 306898 338116
rect 307018 338104 307024 338116
rect 307076 338104 307082 338156
rect 308766 338104 308772 338156
rect 308824 338104 308830 338156
rect 350258 338104 350264 338156
rect 350316 338144 350322 338156
rect 350534 338144 350540 338156
rect 350316 338116 350540 338144
rect 350316 338104 350322 338116
rect 350534 338104 350540 338116
rect 350592 338104 350598 338156
rect 107562 338036 107568 338088
rect 107620 338076 107626 338088
rect 301498 338076 301504 338088
rect 107620 338048 281212 338076
rect 107620 338036 107626 338048
rect 97902 337968 97908 338020
rect 97960 338008 97966 338020
rect 127066 338008 127072 338020
rect 97960 337980 127072 338008
rect 97960 337968 97966 337980
rect 127066 337968 127072 337980
rect 127124 337968 127130 338020
rect 231854 337968 231860 338020
rect 231912 338008 231918 338020
rect 244826 338008 244832 338020
rect 231912 337980 244832 338008
rect 231912 337968 231918 337980
rect 244826 337968 244832 337980
rect 244884 337968 244890 338020
rect 250990 337968 250996 338020
rect 251048 338008 251054 338020
rect 260190 338008 260196 338020
rect 251048 337980 260196 338008
rect 251048 337968 251054 337980
rect 260190 337968 260196 337980
rect 260248 337968 260254 338020
rect 281184 338008 281212 338048
rect 281368 338048 301504 338076
rect 281368 338008 281396 338048
rect 301498 338036 301504 338048
rect 301556 338036 301562 338088
rect 281184 337980 281396 338008
rect 308784 338008 308812 338104
rect 308858 338008 308864 338020
rect 308784 337980 308864 338008
rect 308858 337968 308864 337980
rect 308916 337968 308922 338020
rect 112806 337900 112812 337952
rect 112864 337940 112870 337952
rect 113082 337940 113088 337952
rect 112864 337912 113088 337940
rect 112864 337900 112870 337912
rect 113082 337900 113088 337912
rect 113140 337940 113146 337952
rect 127158 337940 127164 337952
rect 113140 337912 127164 337940
rect 113140 337900 113146 337912
rect 127158 337900 127164 337912
rect 127216 337900 127222 337952
rect 226150 337900 226156 337952
rect 226208 337940 226214 337952
rect 248506 337940 248512 337952
rect 226208 337912 248512 337940
rect 226208 337900 226214 337912
rect 248506 337900 248512 337912
rect 248564 337900 248570 337952
rect 253750 337900 253756 337952
rect 253808 337940 253814 337952
rect 263134 337940 263140 337952
rect 253808 337912 263140 337940
rect 253808 337900 253814 337912
rect 263134 337900 263140 337912
rect 263192 337900 263198 337952
rect 122650 337832 122656 337884
rect 122708 337872 122714 337884
rect 127710 337872 127716 337884
rect 122708 337844 127716 337872
rect 122708 337832 122714 337844
rect 127710 337832 127716 337844
rect 127768 337832 127774 337884
rect 220446 337832 220452 337884
rect 220504 337872 220510 337884
rect 239398 337872 239404 337884
rect 220504 337844 239404 337872
rect 220504 337832 220510 337844
rect 239398 337832 239404 337844
rect 239456 337832 239462 337884
rect 211798 337764 211804 337816
rect 211856 337804 211862 337816
rect 240778 337804 240784 337816
rect 211856 337776 240784 337804
rect 211856 337764 211862 337776
rect 240778 337764 240784 337776
rect 240836 337764 240842 337816
rect 242158 337764 242164 337816
rect 242216 337804 242222 337816
rect 246022 337804 246028 337816
rect 242216 337776 246028 337804
rect 242216 337764 242222 337776
rect 246022 337764 246028 337776
rect 246080 337764 246086 337816
rect 249058 337764 249064 337816
rect 249116 337804 249122 337816
rect 257430 337804 257436 337816
rect 249116 337776 257436 337804
rect 249116 337764 249122 337776
rect 257430 337764 257436 337776
rect 257488 337764 257494 337816
rect 92750 337696 92756 337748
rect 92808 337736 92814 337748
rect 93762 337736 93768 337748
rect 92808 337708 93768 337736
rect 92808 337696 92814 337708
rect 93762 337696 93768 337708
rect 93820 337696 93826 337748
rect 102870 337696 102876 337748
rect 102928 337736 102934 337748
rect 103422 337736 103428 337748
rect 102928 337708 103428 337736
rect 102928 337696 102934 337708
rect 103422 337696 103428 337708
rect 103480 337696 103486 337748
rect 203334 337696 203340 337748
rect 203392 337736 203398 337748
rect 207658 337736 207664 337748
rect 203392 337708 207664 337736
rect 203392 337696 203398 337708
rect 207658 337696 207664 337708
rect 207716 337696 207722 337748
rect 214742 337696 214748 337748
rect 214800 337736 214806 337748
rect 258718 337736 258724 337748
rect 214800 337708 258724 337736
rect 214800 337696 214806 337708
rect 258718 337696 258724 337708
rect 258776 337696 258782 337748
rect 206094 337628 206100 337680
rect 206152 337668 206158 337680
rect 255590 337668 255596 337680
rect 206152 337640 255596 337668
rect 206152 337628 206158 337640
rect 255590 337628 255596 337640
rect 255648 337628 255654 337680
rect 117958 337560 117964 337612
rect 118016 337600 118022 337612
rect 128170 337600 128176 337612
rect 118016 337572 128176 337600
rect 118016 337560 118022 337572
rect 128170 337560 128176 337572
rect 128228 337600 128234 337612
rect 297266 337600 297272 337612
rect 128228 337572 297272 337600
rect 128228 337560 128234 337572
rect 297266 337560 297272 337572
rect 297324 337560 297330 337612
rect 401502 337560 401508 337612
rect 401560 337600 401566 337612
rect 460566 337600 460572 337612
rect 401560 337572 460572 337600
rect 401560 337560 401566 337572
rect 460566 337560 460572 337572
rect 460624 337560 460630 337612
rect 72878 337492 72884 337544
rect 72936 337532 72942 337544
rect 130286 337532 130292 337544
rect 72936 337504 130292 337532
rect 72936 337492 72942 337504
rect 130286 337492 130292 337504
rect 130344 337532 130350 337544
rect 299566 337532 299572 337544
rect 130344 337504 299572 337532
rect 130344 337492 130350 337504
rect 299566 337492 299572 337504
rect 299624 337492 299630 337544
rect 411162 337492 411168 337544
rect 411220 337532 411226 337544
rect 472158 337532 472164 337544
rect 411220 337504 472164 337532
rect 411220 337492 411226 337504
rect 472158 337492 472164 337504
rect 472216 337492 472222 337544
rect 77846 337424 77852 337476
rect 77904 337464 77910 337476
rect 99282 337464 99288 337476
rect 77904 337436 99288 337464
rect 77904 337424 77910 337436
rect 99282 337424 99288 337436
rect 99340 337464 99346 337476
rect 329834 337464 329840 337476
rect 99340 337436 329840 337464
rect 99340 337424 99346 337436
rect 329834 337424 329840 337436
rect 329892 337424 329898 337476
rect 408402 337424 408408 337476
rect 408460 337464 408466 337476
rect 483750 337464 483756 337476
rect 408460 337436 483756 337464
rect 408460 337424 408466 337436
rect 483750 337424 483756 337436
rect 483808 337424 483814 337476
rect 87782 337356 87788 337408
rect 87840 337396 87846 337408
rect 117222 337396 117228 337408
rect 87840 337368 117228 337396
rect 87840 337356 87846 337368
rect 117222 337356 117228 337368
rect 117280 337396 117286 337408
rect 380434 337396 380440 337408
rect 117280 337368 380440 337396
rect 117280 337356 117286 337368
rect 380434 337356 380440 337368
rect 380492 337356 380498 337408
rect 413922 337356 413928 337408
rect 413980 337396 413986 337408
rect 495342 337396 495348 337408
rect 413980 337368 495348 337396
rect 413980 337356 413986 337368
rect 495342 337356 495348 337368
rect 495400 337356 495406 337408
rect 223206 337288 223212 337340
rect 223264 337328 223270 337340
rect 237650 337328 237656 337340
rect 223264 337300 237656 337328
rect 223264 337288 223270 337300
rect 237650 337288 237656 337300
rect 237708 337288 237714 337340
rect 239398 337288 239404 337340
rect 239456 337328 239462 337340
rect 246298 337328 246304 337340
rect 239456 337300 246304 337328
rect 239456 337288 239462 337300
rect 246298 337288 246304 337300
rect 246356 337288 246362 337340
rect 228910 337220 228916 337272
rect 228968 337260 228974 337272
rect 235994 337260 236000 337272
rect 228968 337232 236000 337260
rect 228968 337220 228974 337232
rect 235994 337220 236000 337232
rect 236052 337220 236058 337272
rect 242802 337220 242808 337272
rect 242860 337260 242866 337272
rect 249058 337260 249064 337272
rect 242860 337232 249064 337260
rect 242860 337220 242866 337232
rect 249058 337220 249064 337232
rect 249116 337220 249122 337272
rect 251726 337220 251732 337272
rect 251784 337260 251790 337272
rect 260098 337260 260104 337272
rect 251784 337232 260104 337260
rect 251784 337220 251790 337232
rect 260098 337220 260104 337232
rect 260156 337220 260162 337272
rect 271782 336880 271788 336932
rect 271840 336880 271846 336932
rect 200574 336812 200580 336864
rect 200632 336852 200638 336864
rect 201402 336852 201408 336864
rect 200632 336824 201408 336852
rect 200632 336812 200638 336824
rect 201402 336812 201408 336824
rect 201460 336812 201466 336864
rect 234614 336812 234620 336864
rect 234672 336852 234678 336864
rect 237466 336852 237472 336864
rect 234672 336824 237472 336852
rect 234672 336812 234678 336824
rect 237466 336812 237472 336824
rect 237524 336812 237530 336864
rect 237558 336812 237564 336864
rect 237616 336852 237622 336864
rect 239398 336852 239404 336864
rect 237616 336824 239404 336852
rect 237616 336812 237622 336824
rect 239398 336812 239404 336824
rect 239456 336812 239462 336864
rect 240042 336812 240048 336864
rect 240100 336852 240106 336864
rect 243078 336852 243084 336864
rect 240100 336824 243084 336852
rect 240100 336812 240106 336824
rect 243078 336812 243084 336824
rect 243136 336812 243142 336864
rect 247678 336812 247684 336864
rect 247736 336852 247742 336864
rect 248782 336852 248788 336864
rect 247736 336824 248788 336852
rect 247736 336812 247742 336824
rect 248782 336812 248788 336824
rect 248840 336812 248846 336864
rect 254486 336812 254492 336864
rect 254544 336852 254550 336864
rect 258442 336852 258448 336864
rect 254544 336824 258448 336852
rect 254544 336812 254550 336824
rect 258442 336812 258448 336824
rect 258500 336812 258506 336864
rect 265894 336812 265900 336864
rect 265952 336852 265958 336864
rect 269666 336852 269672 336864
rect 265952 336824 269672 336852
rect 265952 336812 265958 336824
rect 269666 336812 269672 336824
rect 269724 336812 269730 336864
rect 271690 336812 271696 336864
rect 271748 336852 271754 336864
rect 271800 336852 271828 336880
rect 271748 336824 271828 336852
rect 271748 336812 271754 336824
rect 2958 336744 2964 336796
rect 3016 336784 3022 336796
rect 434714 336784 434720 336796
rect 3016 336756 434720 336784
rect 3016 336744 3022 336756
rect 434714 336744 434720 336756
rect 434772 336744 434778 336796
rect 82722 336676 82728 336728
rect 82780 336716 82786 336728
rect 125962 336716 125968 336728
rect 82780 336688 125968 336716
rect 82780 336676 82786 336688
rect 125962 336676 125968 336688
rect 126020 336676 126026 336728
rect 258166 336676 258172 336728
rect 258224 336716 258230 336728
rect 258442 336716 258448 336728
rect 258224 336688 258448 336716
rect 258224 336676 258230 336688
rect 258442 336676 258448 336688
rect 258500 336676 258506 336728
rect 128722 335996 128728 336048
rect 128780 336036 128786 336048
rect 129090 336036 129096 336048
rect 128780 336008 129096 336036
rect 128780 335996 128786 336008
rect 129090 335996 129096 336008
rect 129148 335996 129154 336048
rect 503622 331168 503628 331220
rect 503680 331208 503686 331220
rect 503990 331208 503996 331220
rect 503680 331180 503996 331208
rect 503680 331168 503686 331180
rect 503990 331168 503996 331180
rect 504048 331168 504054 331220
rect 271414 330488 271420 330540
rect 271472 330528 271478 330540
rect 271598 330528 271604 330540
rect 271472 330500 271604 330528
rect 271472 330488 271478 330500
rect 271598 330488 271604 330500
rect 271656 330488 271662 330540
rect 244826 328448 244832 328500
rect 244884 328488 244890 328500
rect 248690 328488 248696 328500
rect 244884 328460 248696 328488
rect 244884 328448 244890 328460
rect 248690 328448 248696 328460
rect 248748 328448 248754 328500
rect 281166 328448 281172 328500
rect 281224 328488 281230 328500
rect 281258 328488 281264 328500
rect 281224 328460 281264 328488
rect 281224 328448 281230 328460
rect 281258 328448 281264 328460
rect 281316 328448 281322 328500
rect 307018 328380 307024 328432
rect 307076 328380 307082 328432
rect 503530 328380 503536 328432
rect 503588 328420 503594 328432
rect 503714 328420 503720 328432
rect 503588 328392 503720 328420
rect 503588 328380 503594 328392
rect 503714 328380 503720 328392
rect 503772 328380 503778 328432
rect 307036 328296 307064 328380
rect 307018 328244 307024 328296
rect 307076 328244 307082 328296
rect 308766 327156 308772 327208
rect 308824 327196 308830 327208
rect 308824 327168 308904 327196
rect 308824 327156 308830 327168
rect 308876 327140 308904 327168
rect 258166 327088 258172 327140
rect 258224 327128 258230 327140
rect 258350 327128 258356 327140
rect 258224 327100 258356 327128
rect 258224 327088 258230 327100
rect 258350 327088 258356 327100
rect 258408 327088 258414 327140
rect 308858 327088 308864 327140
rect 308916 327088 308922 327140
rect 128722 327020 128728 327072
rect 128780 327060 128786 327072
rect 129090 327060 129096 327072
rect 128780 327032 129096 327060
rect 128780 327020 128786 327032
rect 129090 327020 129096 327032
rect 129148 327020 129154 327072
rect 8018 325660 8024 325712
rect 8076 325700 8082 325712
rect 8202 325700 8208 325712
rect 8076 325672 8208 325700
rect 8076 325660 8082 325672
rect 8202 325660 8208 325672
rect 8260 325660 8266 325712
rect 128354 325660 128360 325712
rect 128412 325700 128418 325712
rect 128446 325700 128452 325712
rect 128412 325672 128452 325700
rect 128412 325660 128418 325672
rect 128446 325660 128452 325672
rect 128504 325660 128510 325712
rect 271414 325660 271420 325712
rect 271472 325700 271478 325712
rect 271506 325700 271512 325712
rect 271472 325672 271512 325700
rect 271472 325660 271478 325672
rect 271506 325660 271512 325672
rect 271564 325660 271570 325712
rect 503990 323552 503996 323604
rect 504048 323592 504054 323604
rect 504174 323592 504180 323604
rect 504048 323564 504180 323592
rect 504048 323552 504054 323564
rect 504174 323552 504180 323564
rect 504232 323552 504238 323604
rect 2958 322940 2964 322992
rect 3016 322980 3022 322992
rect 5074 322980 5080 322992
rect 3016 322952 5080 322980
rect 3016 322940 3022 322952
rect 5074 322940 5080 322952
rect 5132 322940 5138 322992
rect 271506 322872 271512 322924
rect 271564 322912 271570 322924
rect 271690 322912 271696 322924
rect 271564 322884 271696 322912
rect 271564 322872 271570 322884
rect 271690 322872 271696 322884
rect 271748 322872 271754 322924
rect 130010 321580 130016 321632
rect 130068 321620 130074 321632
rect 580166 321620 580172 321632
rect 130068 321592 580172 321620
rect 130068 321580 130074 321592
rect 580166 321580 580172 321592
rect 580224 321580 580230 321632
rect 122558 321512 122564 321564
rect 122616 321552 122622 321564
rect 122742 321552 122748 321564
rect 122616 321524 122748 321552
rect 122616 321512 122622 321524
rect 122742 321512 122748 321524
rect 122800 321512 122806 321564
rect 132678 321512 132684 321564
rect 132736 321552 132742 321564
rect 132862 321552 132868 321564
rect 132736 321524 132868 321552
rect 132736 321512 132742 321524
rect 132862 321512 132868 321524
rect 132920 321512 132926 321564
rect 281258 321512 281264 321564
rect 281316 321552 281322 321564
rect 281350 321552 281356 321564
rect 281316 321524 281356 321552
rect 281316 321512 281322 321524
rect 281350 321512 281356 321524
rect 281408 321512 281414 321564
rect 255774 318792 255780 318844
rect 255832 318832 255838 318844
rect 255866 318832 255872 318844
rect 255832 318804 255872 318832
rect 255832 318792 255838 318804
rect 255866 318792 255872 318804
rect 255924 318792 255930 318844
rect 503530 318792 503536 318844
rect 503588 318832 503594 318844
rect 503714 318832 503720 318844
rect 503588 318804 503720 318832
rect 503588 318792 503594 318804
rect 503714 318792 503720 318804
rect 503772 318792 503778 318844
rect 503990 318792 503996 318844
rect 504048 318832 504054 318844
rect 504174 318832 504180 318844
rect 504048 318804 504180 318832
rect 504048 318792 504054 318804
rect 504174 318792 504180 318804
rect 504232 318792 504238 318844
rect 122466 318724 122472 318776
rect 122524 318764 122530 318776
rect 122742 318764 122748 318776
rect 122524 318736 122748 318764
rect 122524 318724 122530 318736
rect 122742 318724 122748 318736
rect 122800 318724 122806 318776
rect 132402 318724 132408 318776
rect 132460 318764 132466 318776
rect 132862 318764 132868 318776
rect 132460 318736 132868 318764
rect 132460 318724 132466 318736
rect 132862 318724 132868 318736
rect 132920 318724 132926 318776
rect 257706 318724 257712 318776
rect 257764 318764 257770 318776
rect 257982 318764 257988 318776
rect 257764 318736 257988 318764
rect 257764 318724 257770 318736
rect 257982 318724 257988 318736
rect 258040 318724 258046 318776
rect 281074 318724 281080 318776
rect 281132 318764 281138 318776
rect 281350 318764 281356 318776
rect 281132 318736 281356 318764
rect 281132 318724 281138 318736
rect 281350 318724 281356 318736
rect 281408 318724 281414 318776
rect 504358 318724 504364 318776
rect 504416 318764 504422 318776
rect 504450 318764 504456 318776
rect 504416 318736 504456 318764
rect 504416 318724 504422 318736
rect 504450 318724 504456 318736
rect 504508 318724 504514 318776
rect 258166 317432 258172 317484
rect 258224 317472 258230 317484
rect 258626 317472 258632 317484
rect 258224 317444 258632 317472
rect 258224 317432 258230 317444
rect 258626 317432 258632 317444
rect 258684 317432 258690 317484
rect 503438 313896 503444 313948
rect 503496 313936 503502 313948
rect 503714 313936 503720 313948
rect 503496 313908 503720 313936
rect 503496 313896 503502 313908
rect 503714 313896 503720 313908
rect 503772 313896 503778 313948
rect 503622 311856 503628 311908
rect 503680 311896 503686 311908
rect 503990 311896 503996 311908
rect 503680 311868 503996 311896
rect 503680 311856 503686 311868
rect 503990 311856 503996 311868
rect 504048 311856 504054 311908
rect 503622 311720 503628 311772
rect 503680 311760 503686 311772
rect 503990 311760 503996 311772
rect 503680 311732 503996 311760
rect 503680 311720 503686 311732
rect 503990 311720 503996 311732
rect 504048 311720 504054 311772
rect 128722 311584 128728 311636
rect 128780 311624 128786 311636
rect 129090 311624 129096 311636
rect 128780 311596 129096 311624
rect 128780 311584 128786 311596
rect 129090 311584 129096 311596
rect 129148 311584 129154 311636
rect 131758 310496 131764 310548
rect 131816 310536 131822 310548
rect 580166 310536 580172 310548
rect 131816 310508 580172 310536
rect 131816 310496 131822 310508
rect 580166 310496 580172 310508
rect 580224 310496 580230 310548
rect 504358 309204 504364 309256
rect 504416 309244 504422 309256
rect 504450 309244 504456 309256
rect 504416 309216 504456 309244
rect 504416 309204 504422 309216
rect 504450 309204 504456 309216
rect 504508 309204 504514 309256
rect 122466 309136 122472 309188
rect 122524 309176 122530 309188
rect 122650 309176 122656 309188
rect 122524 309148 122656 309176
rect 122524 309136 122530 309148
rect 122650 309136 122656 309148
rect 122708 309136 122714 309188
rect 132402 309136 132408 309188
rect 132460 309176 132466 309188
rect 132770 309176 132776 309188
rect 132460 309148 132776 309176
rect 132460 309136 132466 309148
rect 132770 309136 132776 309148
rect 132828 309136 132834 309188
rect 257706 309136 257712 309188
rect 257764 309176 257770 309188
rect 257798 309176 257804 309188
rect 257764 309148 257804 309176
rect 257764 309136 257770 309148
rect 257798 309136 257804 309148
rect 257856 309136 257862 309188
rect 281074 309136 281080 309188
rect 281132 309176 281138 309188
rect 281258 309176 281264 309188
rect 281132 309148 281264 309176
rect 281132 309136 281138 309148
rect 281258 309136 281264 309148
rect 281316 309136 281322 309188
rect 307018 309136 307024 309188
rect 307076 309176 307082 309188
rect 307076 309148 307156 309176
rect 307076 309136 307082 309148
rect 307128 309120 307156 309148
rect 503438 309136 503444 309188
rect 503496 309176 503502 309188
rect 503806 309176 503812 309188
rect 503496 309148 503812 309176
rect 503496 309136 503502 309148
rect 503806 309136 503812 309148
rect 503864 309136 503870 309188
rect 307110 309068 307116 309120
rect 307168 309068 307174 309120
rect 504174 309068 504180 309120
rect 504232 309108 504238 309120
rect 504358 309108 504364 309120
rect 504232 309080 504364 309108
rect 504232 309068 504238 309080
rect 504358 309068 504364 309080
rect 504416 309068 504422 309120
rect 2958 307776 2964 307828
rect 3016 307816 3022 307828
rect 5166 307816 5172 307828
rect 3016 307788 5172 307816
rect 3016 307776 3022 307788
rect 5166 307776 5172 307788
rect 5224 307776 5230 307828
rect 307110 307776 307116 307828
rect 307168 307816 307174 307828
rect 307202 307816 307208 307828
rect 307168 307788 307208 307816
rect 307168 307776 307174 307788
rect 307202 307776 307208 307788
rect 307260 307776 307266 307828
rect 128722 307028 128728 307080
rect 128780 307068 128786 307080
rect 129090 307068 129096 307080
rect 128780 307040 129096 307068
rect 128780 307028 128786 307040
rect 129090 307028 129096 307040
rect 129148 307028 129154 307080
rect 8018 306348 8024 306400
rect 8076 306388 8082 306400
rect 8202 306388 8208 306400
rect 8076 306360 8208 306388
rect 8076 306348 8082 306360
rect 8202 306348 8208 306360
rect 8260 306348 8266 306400
rect 271782 303560 271788 303612
rect 271840 303600 271846 303612
rect 271966 303600 271972 303612
rect 271840 303572 271972 303600
rect 271840 303560 271846 303572
rect 271966 303560 271972 303572
rect 272024 303560 272030 303612
rect 281258 302200 281264 302252
rect 281316 302200 281322 302252
rect 281276 302172 281304 302200
rect 281350 302172 281356 302184
rect 281276 302144 281356 302172
rect 281350 302132 281356 302144
rect 281408 302132 281414 302184
rect 128630 299480 128636 299532
rect 128688 299520 128694 299532
rect 128814 299520 128820 299532
rect 128688 299492 128820 299520
rect 128688 299480 128694 299492
rect 128814 299480 128820 299492
rect 128872 299480 128878 299532
rect 307018 299480 307024 299532
rect 307076 299520 307082 299532
rect 307202 299520 307208 299532
rect 307076 299492 307208 299520
rect 307076 299480 307082 299492
rect 307202 299480 307208 299492
rect 307260 299480 307266 299532
rect 308674 299480 308680 299532
rect 308732 299520 308738 299532
rect 308766 299520 308772 299532
rect 308732 299492 308772 299520
rect 308732 299480 308738 299492
rect 308766 299480 308772 299492
rect 308824 299480 308830 299532
rect 504174 299480 504180 299532
rect 504232 299520 504238 299532
rect 504450 299520 504456 299532
rect 504232 299492 504456 299520
rect 504232 299480 504238 299492
rect 504450 299480 504456 299492
rect 504508 299480 504514 299532
rect 255498 299412 255504 299464
rect 255556 299452 255562 299464
rect 255590 299452 255596 299464
rect 255556 299424 255596 299452
rect 255556 299412 255562 299424
rect 255590 299412 255596 299424
rect 255648 299412 255654 299464
rect 257706 299412 257712 299464
rect 257764 299452 257770 299464
rect 257890 299452 257896 299464
rect 257764 299424 257896 299452
rect 257764 299412 257770 299424
rect 257890 299412 257896 299424
rect 257948 299412 257954 299464
rect 258258 299412 258264 299464
rect 258316 299452 258322 299464
rect 258350 299452 258356 299464
rect 258316 299424 258356 299452
rect 258316 299412 258322 299424
rect 258350 299412 258356 299424
rect 258408 299412 258414 299464
rect 281074 299412 281080 299464
rect 281132 299452 281138 299464
rect 281350 299452 281356 299464
rect 281132 299424 281356 299452
rect 281132 299412 281138 299424
rect 281350 299412 281356 299424
rect 281408 299412 281414 299464
rect 504450 298052 504456 298104
rect 504508 298092 504514 298104
rect 504726 298092 504732 298104
rect 504508 298064 504732 298092
rect 504508 298052 504514 298064
rect 504726 298052 504732 298064
rect 504784 298052 504790 298104
rect 128722 297372 128728 297424
rect 128780 297412 128786 297424
rect 129090 297412 129096 297424
rect 128780 297384 129096 297412
rect 128780 297372 128786 297384
rect 129090 297372 129096 297384
rect 129148 297372 129154 297424
rect 2958 293972 2964 294024
rect 3016 294012 3022 294024
rect 434806 294012 434812 294024
rect 3016 293984 434812 294012
rect 3016 293972 3022 293984
rect 434806 293972 434812 293984
rect 434864 293972 434870 294024
rect 308674 292544 308680 292596
rect 308732 292584 308738 292596
rect 308858 292584 308864 292596
rect 308732 292556 308864 292584
rect 308732 292544 308738 292556
rect 308858 292544 308864 292556
rect 308916 292544 308922 292596
rect 322842 291932 322848 291984
rect 322900 291972 322906 291984
rect 378686 291972 378692 291984
rect 322900 291944 378692 291972
rect 322900 291932 322906 291944
rect 378686 291932 378692 291944
rect 378744 291932 378750 291984
rect 300762 291864 300768 291916
rect 300820 291904 300826 291916
rect 378594 291904 378600 291916
rect 300820 291876 378600 291904
rect 300820 291864 300826 291876
rect 378594 291864 378600 291876
rect 378652 291864 378658 291916
rect 198918 291796 198924 291848
rect 198976 291836 198982 291848
rect 231854 291836 231860 291848
rect 198976 291808 231860 291836
rect 198976 291796 198982 291808
rect 231854 291796 231860 291808
rect 231912 291796 231918 291848
rect 300670 291796 300676 291848
rect 300728 291836 300734 291848
rect 378870 291836 378876 291848
rect 300728 291808 378876 291836
rect 300728 291796 300734 291808
rect 378870 291796 378876 291808
rect 378928 291796 378934 291848
rect 128446 290436 128452 290488
rect 128504 290476 128510 290488
rect 128630 290476 128636 290488
rect 128504 290448 128636 290476
rect 128504 290436 128510 290448
rect 128630 290436 128636 290448
rect 128688 290436 128694 290488
rect 255498 289892 255504 289944
rect 255556 289932 255562 289944
rect 255556 289904 255636 289932
rect 255556 289892 255562 289904
rect 255608 289876 255636 289904
rect 258258 289892 258264 289944
rect 258316 289932 258322 289944
rect 258316 289904 258396 289932
rect 258316 289892 258322 289904
rect 258368 289876 258396 289904
rect 255590 289824 255596 289876
rect 255648 289824 255654 289876
rect 257706 289824 257712 289876
rect 257764 289864 257770 289876
rect 257798 289864 257804 289876
rect 257764 289836 257804 289864
rect 257764 289824 257770 289836
rect 257798 289824 257804 289836
rect 257856 289824 257862 289876
rect 258350 289824 258356 289876
rect 258408 289824 258414 289876
rect 281074 289824 281080 289876
rect 281132 289864 281138 289876
rect 281258 289864 281264 289876
rect 281132 289836 281264 289864
rect 281132 289824 281138 289836
rect 281258 289824 281264 289836
rect 281316 289824 281322 289876
rect 504542 288396 504548 288448
rect 504600 288436 504606 288448
rect 504726 288436 504732 288448
rect 504600 288408 504732 288436
rect 504600 288396 504606 288408
rect 504726 288396 504732 288408
rect 504784 288396 504790 288448
rect 128722 287716 128728 287768
rect 128780 287756 128786 287768
rect 129090 287756 129096 287768
rect 128780 287728 129096 287756
rect 128780 287716 128786 287728
rect 129090 287716 129096 287728
rect 129148 287716 129154 287768
rect 8018 287036 8024 287088
rect 8076 287076 8082 287088
rect 8202 287076 8208 287088
rect 8076 287048 8208 287076
rect 8076 287036 8082 287048
rect 8202 287036 8208 287048
rect 8260 287036 8266 287088
rect 271782 284248 271788 284300
rect 271840 284288 271846 284300
rect 271966 284288 271972 284300
rect 271840 284260 271972 284288
rect 271840 284248 271846 284260
rect 271966 284248 271972 284260
rect 272024 284248 272030 284300
rect 308582 283568 308588 283620
rect 308640 283608 308646 283620
rect 308858 283608 308864 283620
rect 308640 283580 308864 283608
rect 308640 283568 308646 283580
rect 308858 283568 308864 283580
rect 308916 283568 308922 283620
rect 503714 283024 503720 283076
rect 503772 283064 503778 283076
rect 503772 283036 503852 283064
rect 503772 283024 503778 283036
rect 503824 283008 503852 283036
rect 503806 282956 503812 283008
rect 503864 282956 503870 283008
rect 132678 282888 132684 282940
rect 132736 282928 132742 282940
rect 132862 282928 132868 282940
rect 132736 282900 132868 282928
rect 132736 282888 132742 282900
rect 132862 282888 132868 282900
rect 132920 282888 132926 282940
rect 257798 282888 257804 282940
rect 257856 282928 257862 282940
rect 257982 282928 257988 282940
rect 257856 282900 257988 282928
rect 257856 282888 257862 282900
rect 257982 282888 257988 282900
rect 258040 282888 258046 282940
rect 281258 282888 281264 282940
rect 281316 282888 281322 282940
rect 281276 282860 281304 282888
rect 281350 282860 281356 282872
rect 281276 282832 281356 282860
rect 281350 282820 281356 282832
rect 281408 282820 281414 282872
rect 128446 280100 128452 280152
rect 128504 280140 128510 280152
rect 128630 280140 128636 280152
rect 128504 280112 128636 280140
rect 128504 280100 128510 280112
rect 128630 280100 128636 280112
rect 128688 280100 128694 280152
rect 281350 280100 281356 280152
rect 281408 280140 281414 280152
rect 281626 280140 281632 280152
rect 281408 280112 281632 280140
rect 281408 280100 281414 280112
rect 281626 280100 281632 280112
rect 281684 280100 281690 280152
rect 308582 278740 308588 278792
rect 308640 278780 308646 278792
rect 308674 278780 308680 278792
rect 308640 278752 308680 278780
rect 308640 278740 308646 278752
rect 308674 278740 308680 278752
rect 308732 278740 308738 278792
rect 504450 278672 504456 278724
rect 504508 278712 504514 278724
rect 504542 278712 504548 278724
rect 504508 278684 504548 278712
rect 504508 278672 504514 278684
rect 504542 278672 504548 278684
rect 504600 278672 504606 278724
rect 258258 275952 258264 276004
rect 258316 275992 258322 276004
rect 258350 275992 258356 276004
rect 258316 275964 258356 275992
rect 258316 275952 258322 275964
rect 258350 275952 258356 275964
rect 258408 275952 258414 276004
rect 131574 274660 131580 274712
rect 131632 274700 131638 274712
rect 579982 274700 579988 274712
rect 131632 274672 579988 274700
rect 131632 274660 131638 274672
rect 579982 274660 579988 274672
rect 580040 274660 580046 274712
rect 128722 274252 128728 274304
rect 128780 274292 128786 274304
rect 129090 274292 129096 274304
rect 128780 274264 129096 274292
rect 128780 274252 128786 274264
rect 129090 274252 129096 274264
rect 129148 274252 129154 274304
rect 503622 273300 503628 273352
rect 503680 273340 503686 273352
rect 503990 273340 503996 273352
rect 503680 273312 503996 273340
rect 503680 273300 503686 273312
rect 503990 273300 503996 273312
rect 504048 273300 504054 273352
rect 503622 273164 503628 273216
rect 503680 273204 503686 273216
rect 503990 273204 503996 273216
rect 503680 273176 503996 273204
rect 503680 273164 503686 273176
rect 503990 273164 503996 273176
rect 504048 273164 504054 273216
rect 281350 270580 281356 270632
rect 281408 270620 281414 270632
rect 281626 270620 281632 270632
rect 281408 270592 281632 270620
rect 281408 270580 281414 270592
rect 281626 270580 281632 270592
rect 281684 270580 281690 270632
rect 128446 270512 128452 270564
rect 128504 270552 128510 270564
rect 128630 270552 128636 270564
rect 128504 270524 128636 270552
rect 128504 270512 128510 270524
rect 128630 270512 128636 270524
rect 128688 270512 128694 270564
rect 307018 270552 307024 270564
rect 306944 270524 307024 270552
rect 306944 270496 306972 270524
rect 307018 270512 307024 270524
rect 307076 270512 307082 270564
rect 281074 270444 281080 270496
rect 281132 270484 281138 270496
rect 281350 270484 281356 270496
rect 281132 270456 281356 270484
rect 281132 270444 281138 270456
rect 281350 270444 281356 270456
rect 281408 270444 281414 270496
rect 306926 270444 306932 270496
rect 306984 270444 306990 270496
rect 308674 269084 308680 269136
rect 308732 269124 308738 269136
rect 308858 269124 308864 269136
rect 308732 269096 308864 269124
rect 308732 269084 308738 269096
rect 308858 269084 308864 269096
rect 308916 269084 308922 269136
rect 306742 269016 306748 269068
rect 306800 269056 306806 269068
rect 306926 269056 306932 269068
rect 306800 269028 306932 269056
rect 306800 269016 306806 269028
rect 306926 269016 306932 269028
rect 306984 269016 306990 269068
rect 128722 268404 128728 268456
rect 128780 268444 128786 268456
rect 129090 268444 129096 268456
rect 128780 268416 129096 268444
rect 128780 268404 128786 268416
rect 129090 268404 129096 268416
rect 129148 268404 129154 268456
rect 8018 267724 8024 267776
rect 8076 267764 8082 267776
rect 8202 267764 8208 267776
rect 8076 267736 8208 267764
rect 8076 267724 8082 267736
rect 8202 267724 8208 267736
rect 8260 267724 8266 267776
rect 2866 264936 2872 264988
rect 2924 264976 2930 264988
rect 5258 264976 5264 264988
rect 2924 264948 5264 264976
rect 2924 264936 2930 264948
rect 5258 264936 5264 264948
rect 5316 264936 5322 264988
rect 271598 264868 271604 264920
rect 271656 264908 271662 264920
rect 271782 264908 271788 264920
rect 271656 264880 271788 264908
rect 271656 264868 271662 264880
rect 271782 264868 271788 264880
rect 271840 264868 271846 264920
rect 503714 263644 503720 263696
rect 503772 263684 503778 263696
rect 503990 263684 503996 263696
rect 503772 263656 503996 263684
rect 503772 263644 503778 263656
rect 503990 263644 503996 263656
rect 504048 263644 504054 263696
rect 131666 263576 131672 263628
rect 131724 263616 131730 263628
rect 580166 263616 580172 263628
rect 131724 263588 580172 263616
rect 131724 263576 131730 263588
rect 580166 263576 580172 263588
rect 580224 263576 580230 263628
rect 503714 263508 503720 263560
rect 503772 263548 503778 263560
rect 503990 263548 503996 263560
rect 503772 263520 503996 263548
rect 503772 263508 503778 263520
rect 503990 263508 503996 263520
rect 504048 263508 504054 263560
rect 255682 260856 255688 260908
rect 255740 260856 255746 260908
rect 281074 260856 281080 260908
rect 281132 260896 281138 260908
rect 281258 260896 281264 260908
rect 281132 260868 281264 260896
rect 281132 260856 281138 260868
rect 281258 260856 281264 260868
rect 281316 260856 281322 260908
rect 128078 260788 128084 260840
rect 128136 260828 128142 260840
rect 128538 260828 128544 260840
rect 128136 260800 128544 260828
rect 128136 260788 128142 260800
rect 128538 260788 128544 260800
rect 128596 260788 128602 260840
rect 255700 260772 255728 260856
rect 504266 260788 504272 260840
rect 504324 260828 504330 260840
rect 504542 260828 504548 260840
rect 504324 260800 504548 260828
rect 504324 260788 504330 260800
rect 504542 260788 504548 260800
rect 504600 260788 504606 260840
rect 255682 260720 255688 260772
rect 255740 260720 255746 260772
rect 306742 259428 306748 259480
rect 306800 259468 306806 259480
rect 307018 259468 307024 259480
rect 306800 259440 307024 259468
rect 306800 259428 306806 259440
rect 307018 259428 307024 259440
rect 307076 259428 307082 259480
rect 128722 258748 128728 258800
rect 128780 258788 128786 258800
rect 129090 258788 129096 258800
rect 128780 258760 129096 258788
rect 128780 258748 128786 258760
rect 129090 258748 129096 258760
rect 129148 258748 129154 258800
rect 271414 255212 271420 255264
rect 271472 255252 271478 255264
rect 271782 255252 271788 255264
rect 271472 255224 271788 255252
rect 271472 255212 271478 255224
rect 271782 255212 271788 255224
rect 271840 255212 271846 255264
rect 503622 253988 503628 254040
rect 503680 254028 503686 254040
rect 503990 254028 503996 254040
rect 503680 254000 503996 254028
rect 503680 253988 503686 254000
rect 503990 253988 503996 254000
rect 504048 253988 504054 254040
rect 503622 253852 503628 253904
rect 503680 253892 503686 253904
rect 503990 253892 503996 253904
rect 503680 253864 503996 253892
rect 503680 253852 503686 253864
rect 503990 253852 503996 253864
rect 504048 253852 504054 253904
rect 504266 253784 504272 253836
rect 504324 253824 504330 253836
rect 504542 253824 504548 253836
rect 504324 253796 504548 253824
rect 504324 253784 504330 253796
rect 504542 253784 504548 253796
rect 504600 253784 504606 253836
rect 307018 251472 307024 251524
rect 307076 251472 307082 251524
rect 307036 251388 307064 251472
rect 307018 251336 307024 251388
rect 307076 251336 307082 251388
rect 2866 251200 2872 251252
rect 2924 251240 2930 251252
rect 434898 251240 434904 251252
rect 2924 251212 434904 251240
rect 2924 251200 2930 251212
rect 434898 251200 434904 251212
rect 434956 251200 434962 251252
rect 7742 251132 7748 251184
rect 7800 251172 7806 251184
rect 7926 251172 7932 251184
rect 7800 251144 7932 251172
rect 7800 251132 7806 251144
rect 7926 251132 7932 251144
rect 7984 251132 7990 251184
rect 504082 251132 504088 251184
rect 504140 251172 504146 251184
rect 504266 251172 504272 251184
rect 504140 251144 504272 251172
rect 504140 251132 504146 251144
rect 504266 251132 504272 251144
rect 504324 251132 504330 251184
rect 128722 249092 128728 249144
rect 128780 249132 128786 249144
rect 129090 249132 129096 249144
rect 128780 249104 129096 249132
rect 128780 249092 128786 249104
rect 129090 249092 129096 249104
rect 129148 249092 129154 249144
rect 258442 249092 258448 249144
rect 258500 249092 258506 249144
rect 258460 249008 258488 249092
rect 258442 248956 258448 249008
rect 258500 248956 258506 249008
rect 271414 245624 271420 245676
rect 271472 245664 271478 245676
rect 271506 245664 271512 245676
rect 271472 245636 271512 245664
rect 271472 245624 271478 245636
rect 271506 245624 271512 245636
rect 271564 245624 271570 245676
rect 308582 245352 308588 245404
rect 308640 245392 308646 245404
rect 308858 245392 308864 245404
rect 308640 245364 308864 245392
rect 308640 245352 308646 245364
rect 308858 245352 308864 245364
rect 308916 245352 308922 245404
rect 503714 244400 503720 244452
rect 503772 244440 503778 244452
rect 503772 244412 503852 244440
rect 503772 244400 503778 244412
rect 503824 244384 503852 244412
rect 503806 244332 503812 244384
rect 503864 244332 503870 244384
rect 271506 242156 271512 242208
rect 271564 242196 271570 242208
rect 271782 242196 271788 242208
rect 271564 242168 271788 242196
rect 271564 242156 271570 242168
rect 271782 242156 271788 242168
rect 271840 242156 271846 242208
rect 307018 241544 307024 241596
rect 307076 241584 307082 241596
rect 307202 241584 307208 241596
rect 307076 241556 307208 241584
rect 307076 241544 307082 241556
rect 307202 241544 307208 241556
rect 307260 241544 307266 241596
rect 7742 241476 7748 241528
rect 7800 241516 7806 241528
rect 8018 241516 8024 241528
rect 7800 241488 8024 241516
rect 7800 241476 7806 241488
rect 8018 241476 8024 241488
rect 8076 241476 8082 241528
rect 281074 241476 281080 241528
rect 281132 241516 281138 241528
rect 281258 241516 281264 241528
rect 281132 241488 281264 241516
rect 281132 241476 281138 241488
rect 281258 241476 281264 241488
rect 281316 241476 281322 241528
rect 504082 241476 504088 241528
rect 504140 241516 504146 241528
rect 504450 241516 504456 241528
rect 504140 241488 504456 241516
rect 504140 241476 504146 241488
rect 504450 241476 504456 241488
rect 504508 241476 504514 241528
rect 281074 241340 281080 241392
rect 281132 241380 281138 241392
rect 281258 241380 281264 241392
rect 281132 241352 281264 241380
rect 281132 241340 281138 241352
rect 281258 241340 281264 241352
rect 281316 241340 281322 241392
rect 258258 240116 258264 240168
rect 258316 240156 258322 240168
rect 258442 240156 258448 240168
rect 258316 240128 258448 240156
rect 258316 240116 258322 240128
rect 258442 240116 258448 240128
rect 258500 240116 258506 240168
rect 128722 239436 128728 239488
rect 128780 239476 128786 239488
rect 129090 239476 129096 239488
rect 128780 239448 129096 239476
rect 128780 239436 128786 239448
rect 129090 239436 129096 239448
rect 129148 239436 129154 239488
rect 258258 238688 258264 238740
rect 258316 238728 258322 238740
rect 258442 238728 258448 238740
rect 258316 238700 258448 238728
rect 258316 238688 258322 238700
rect 258442 238688 258448 238700
rect 258500 238688 258506 238740
rect 255406 236648 255412 236700
rect 255464 236688 255470 236700
rect 255590 236688 255596 236700
rect 255464 236660 255596 236688
rect 255464 236648 255470 236660
rect 255590 236648 255596 236660
rect 255648 236648 255654 236700
rect 308582 235288 308588 235340
rect 308640 235328 308646 235340
rect 308766 235328 308772 235340
rect 308640 235300 308772 235328
rect 308640 235288 308646 235300
rect 308766 235288 308772 235300
rect 308824 235288 308830 235340
rect 8018 234716 8024 234728
rect 7944 234688 8024 234716
rect 7944 234592 7972 234688
rect 8018 234676 8024 234688
rect 8076 234676 8082 234728
rect 503622 234676 503628 234728
rect 503680 234716 503686 234728
rect 503990 234716 503996 234728
rect 503680 234688 503996 234716
rect 503680 234676 503686 234688
rect 503990 234676 503996 234688
rect 504048 234676 504054 234728
rect 504450 234716 504456 234728
rect 504376 234688 504456 234716
rect 504376 234592 504404 234688
rect 504450 234676 504456 234688
rect 504508 234676 504514 234728
rect 7926 234540 7932 234592
rect 7984 234540 7990 234592
rect 503622 234540 503628 234592
rect 503680 234580 503686 234592
rect 503990 234580 503996 234592
rect 503680 234552 503996 234580
rect 503680 234540 503686 234552
rect 503990 234540 503996 234552
rect 504048 234540 504054 234592
rect 504358 234540 504364 234592
rect 504416 234540 504422 234592
rect 128630 231820 128636 231872
rect 128688 231860 128694 231872
rect 128814 231860 128820 231872
rect 128688 231832 128820 231860
rect 128688 231820 128694 231832
rect 128814 231820 128820 231832
rect 128872 231820 128878 231872
rect 257982 231820 257988 231872
rect 258040 231860 258046 231872
rect 258166 231860 258172 231872
rect 258040 231832 258172 231860
rect 258040 231820 258046 231832
rect 258166 231820 258172 231832
rect 258224 231820 258230 231872
rect 281074 231820 281080 231872
rect 281132 231860 281138 231872
rect 281258 231860 281264 231872
rect 281132 231832 281264 231860
rect 281132 231820 281138 231832
rect 281258 231820 281264 231832
rect 281316 231820 281322 231872
rect 306926 231820 306932 231872
rect 306984 231820 306990 231872
rect 7742 231752 7748 231804
rect 7800 231792 7806 231804
rect 7926 231792 7932 231804
rect 7800 231764 7932 231792
rect 7800 231752 7806 231764
rect 7926 231752 7932 231764
rect 7984 231752 7990 231804
rect 306944 231792 306972 231820
rect 307018 231792 307024 231804
rect 306944 231764 307024 231792
rect 307018 231752 307024 231764
rect 307076 231752 307082 231804
rect 504174 231752 504180 231804
rect 504232 231792 504238 231804
rect 504358 231792 504364 231804
rect 504232 231764 504364 231792
rect 504232 231752 504238 231764
rect 504358 231752 504364 231764
rect 504416 231752 504422 231804
rect 306926 230460 306932 230512
rect 306984 230500 306990 230512
rect 307018 230500 307024 230512
rect 306984 230472 307024 230500
rect 306984 230460 306990 230472
rect 307018 230460 307024 230472
rect 307076 230460 307082 230512
rect 128722 229712 128728 229764
rect 128780 229752 128786 229764
rect 129090 229752 129096 229764
rect 128780 229724 129096 229752
rect 128780 229712 128786 229724
rect 129090 229712 129096 229724
rect 129148 229712 129154 229764
rect 132678 227740 132684 227792
rect 132736 227780 132742 227792
rect 580074 227780 580080 227792
rect 132736 227752 580080 227780
rect 132736 227740 132742 227752
rect 580074 227740 580080 227752
rect 580132 227740 580138 227792
rect 271690 227672 271696 227724
rect 271748 227712 271754 227724
rect 271874 227712 271880 227724
rect 271748 227684 271880 227712
rect 271748 227672 271754 227684
rect 271874 227672 271880 227684
rect 271932 227672 271938 227724
rect 503714 225088 503720 225140
rect 503772 225128 503778 225140
rect 503772 225100 503852 225128
rect 503772 225088 503778 225100
rect 503824 225072 503852 225100
rect 503806 225020 503812 225072
rect 503864 225020 503870 225072
rect 122558 224884 122564 224936
rect 122616 224924 122622 224936
rect 122742 224924 122748 224936
rect 122616 224896 122748 224924
rect 122616 224884 122622 224896
rect 122742 224884 122748 224896
rect 122800 224884 122806 224936
rect 2774 222504 2780 222556
rect 2832 222544 2838 222556
rect 6178 222544 6184 222556
rect 2832 222516 6184 222544
rect 2832 222504 2838 222516
rect 6178 222504 6184 222516
rect 6236 222504 6242 222556
rect 7742 222164 7748 222216
rect 7800 222204 7806 222216
rect 8018 222204 8024 222216
rect 7800 222176 8024 222204
rect 7800 222164 7806 222176
rect 8018 222164 8024 222176
rect 8076 222164 8082 222216
rect 255590 222164 255596 222216
rect 255648 222204 255654 222216
rect 255682 222204 255688 222216
rect 255648 222176 255688 222204
rect 255648 222164 255654 222176
rect 255682 222164 255688 222176
rect 255740 222164 255746 222216
rect 281074 222164 281080 222216
rect 281132 222204 281138 222216
rect 281166 222204 281172 222216
rect 281132 222176 281172 222204
rect 281132 222164 281138 222176
rect 281166 222164 281172 222176
rect 281224 222164 281230 222216
rect 308674 222164 308680 222216
rect 308732 222204 308738 222216
rect 308732 222176 308812 222204
rect 308732 222164 308738 222176
rect 308784 222148 308812 222176
rect 504174 222164 504180 222216
rect 504232 222204 504238 222216
rect 504450 222204 504456 222216
rect 504232 222176 504456 222204
rect 504232 222164 504238 222176
rect 504450 222164 504456 222176
rect 504508 222164 504514 222216
rect 213914 222096 213920 222148
rect 213972 222136 213978 222148
rect 214190 222136 214196 222148
rect 213972 222108 214196 222136
rect 213972 222096 213978 222108
rect 214190 222096 214196 222108
rect 214248 222096 214254 222148
rect 307018 222096 307024 222148
rect 307076 222136 307082 222148
rect 307110 222136 307116 222148
rect 307076 222108 307116 222136
rect 307076 222096 307082 222108
rect 307110 222096 307116 222108
rect 307168 222096 307174 222148
rect 308766 222096 308772 222148
rect 308824 222096 308830 222148
rect 308674 220804 308680 220856
rect 308732 220844 308738 220856
rect 308766 220844 308772 220856
rect 308732 220816 308772 220844
rect 308732 220804 308738 220816
rect 308766 220804 308772 220816
rect 308824 220804 308830 220856
rect 128722 220056 128728 220108
rect 128780 220096 128786 220108
rect 129090 220096 129096 220108
rect 128780 220068 129096 220096
rect 128780 220056 128786 220068
rect 129090 220056 129096 220068
rect 129148 220056 129154 220108
rect 271690 218016 271696 218068
rect 271748 218056 271754 218068
rect 271966 218056 271972 218068
rect 271748 218028 271972 218056
rect 271748 218016 271754 218028
rect 271966 218016 271972 218028
rect 272024 218016 272030 218068
rect 132770 216656 132776 216708
rect 132828 216696 132834 216708
rect 579798 216696 579804 216708
rect 132828 216668 579804 216696
rect 132828 216656 132834 216668
rect 579798 216656 579804 216668
rect 579856 216656 579862 216708
rect 308306 215976 308312 216028
rect 308364 216016 308370 216028
rect 308674 216016 308680 216028
rect 308364 215988 308680 216016
rect 308364 215976 308370 215988
rect 308674 215976 308680 215988
rect 308732 215976 308738 216028
rect 8018 215404 8024 215416
rect 7944 215376 8024 215404
rect 7944 215280 7972 215376
rect 8018 215364 8024 215376
rect 8076 215364 8082 215416
rect 122742 215404 122748 215416
rect 122668 215376 122748 215404
rect 122668 215280 122696 215376
rect 122742 215364 122748 215376
rect 122800 215364 122806 215416
rect 128446 215364 128452 215416
rect 128504 215364 128510 215416
rect 258534 215404 258540 215416
rect 258460 215376 258540 215404
rect 128464 215280 128492 215364
rect 258460 215280 258488 215376
rect 258534 215364 258540 215376
rect 258592 215364 258598 215416
rect 503622 215364 503628 215416
rect 503680 215404 503686 215416
rect 503990 215404 503996 215416
rect 503680 215376 503996 215404
rect 503680 215364 503686 215376
rect 503990 215364 503996 215376
rect 504048 215364 504054 215416
rect 504450 215404 504456 215416
rect 504284 215376 504456 215404
rect 281166 215296 281172 215348
rect 281224 215296 281230 215348
rect 7926 215228 7932 215280
rect 7984 215228 7990 215280
rect 122650 215228 122656 215280
rect 122708 215228 122714 215280
rect 128446 215228 128452 215280
rect 128504 215228 128510 215280
rect 258442 215228 258448 215280
rect 258500 215228 258506 215280
rect 281184 215200 281212 215296
rect 504284 215280 504312 215376
rect 504450 215364 504456 215376
rect 504508 215364 504514 215416
rect 297266 215228 297272 215280
rect 297324 215268 297330 215280
rect 298002 215268 298008 215280
rect 297324 215240 298008 215268
rect 297324 215228 297330 215240
rect 298002 215228 298008 215240
rect 298060 215228 298066 215280
rect 503622 215228 503628 215280
rect 503680 215268 503686 215280
rect 503990 215268 503996 215280
rect 503680 215240 503996 215268
rect 503680 215228 503686 215240
rect 503990 215228 503996 215240
rect 504048 215228 504054 215280
rect 504266 215228 504272 215280
rect 504324 215228 504330 215280
rect 281258 215200 281264 215212
rect 281184 215172 281264 215200
rect 281258 215160 281264 215172
rect 281316 215160 281322 215212
rect 214190 212508 214196 212560
rect 214248 212548 214254 212560
rect 214374 212548 214380 212560
rect 214248 212520 214380 212548
rect 214248 212508 214254 212520
rect 214374 212508 214380 212520
rect 214432 212508 214438 212560
rect 255590 212508 255596 212560
rect 255648 212548 255654 212560
rect 255682 212548 255688 212560
rect 255648 212520 255688 212548
rect 255648 212508 255654 212520
rect 255682 212508 255688 212520
rect 255740 212508 255746 212560
rect 257798 212508 257804 212560
rect 257856 212548 257862 212560
rect 257982 212548 257988 212560
rect 257856 212520 257988 212548
rect 257856 212508 257862 212520
rect 257982 212508 257988 212520
rect 258040 212508 258046 212560
rect 271506 212508 271512 212560
rect 271564 212548 271570 212560
rect 271966 212548 271972 212560
rect 271564 212520 271972 212548
rect 271564 212508 271570 212520
rect 271966 212508 271972 212520
rect 272024 212508 272030 212560
rect 275646 212508 275652 212560
rect 275704 212548 275710 212560
rect 275922 212548 275928 212560
rect 275704 212520 275928 212548
rect 275704 212508 275710 212520
rect 275922 212508 275928 212520
rect 275980 212508 275986 212560
rect 307018 212508 307024 212560
rect 307076 212548 307082 212560
rect 307202 212548 307208 212560
rect 307076 212520 307208 212548
rect 307076 212508 307082 212520
rect 307202 212508 307208 212520
rect 307260 212508 307266 212560
rect 255590 211488 255596 211540
rect 255648 211528 255654 211540
rect 256142 211528 256148 211540
rect 255648 211500 256148 211528
rect 255648 211488 255654 211500
rect 256142 211488 256148 211500
rect 256200 211488 256206 211540
rect 297818 211080 297824 211132
rect 297876 211120 297882 211132
rect 303890 211120 303896 211132
rect 297876 211092 303896 211120
rect 297876 211080 297882 211092
rect 303890 211080 303896 211092
rect 303948 211080 303954 211132
rect 2774 210400 2780 210452
rect 2832 210440 2838 210452
rect 3050 210440 3056 210452
rect 2832 210412 3056 210440
rect 2832 210400 2838 210412
rect 3050 210400 3056 210412
rect 3108 210400 3114 210452
rect 128722 210400 128728 210452
rect 128780 210440 128786 210452
rect 129090 210440 129096 210452
rect 128780 210412 129096 210440
rect 128780 210400 128786 210412
rect 129090 210400 129096 210412
rect 129148 210400 129154 210452
rect 132862 210400 132868 210452
rect 132920 210440 132926 210452
rect 133506 210440 133512 210452
rect 132920 210412 133512 210440
rect 132920 210400 132926 210412
rect 133506 210400 133512 210412
rect 133564 210400 133570 210452
rect 268470 210400 268476 210452
rect 268528 210440 268534 210452
rect 268838 210440 268844 210452
rect 268528 210412 268844 210440
rect 268528 210400 268534 210412
rect 268838 210400 268844 210412
rect 268896 210400 268902 210452
rect 290918 210400 290924 210452
rect 290976 210440 290982 210452
rect 291102 210440 291108 210452
rect 290976 210412 291108 210440
rect 290976 210400 290982 210412
rect 291102 210400 291108 210412
rect 291160 210400 291166 210452
rect 297726 210400 297732 210452
rect 297784 210440 297790 210452
rect 311986 210440 311992 210452
rect 297784 210412 311992 210440
rect 297784 210400 297790 210412
rect 311986 210400 311992 210412
rect 312044 210400 312050 210452
rect 3050 207000 3056 207052
rect 3108 207040 3114 207052
rect 434990 207040 434996 207052
rect 3108 207012 434996 207040
rect 3108 207000 3114 207012
rect 434990 207000 434996 207012
rect 435048 207000 435054 207052
rect 503714 205776 503720 205828
rect 503772 205816 503778 205828
rect 503772 205788 503852 205816
rect 503772 205776 503778 205788
rect 503824 205760 503852 205788
rect 503806 205708 503812 205760
rect 503864 205708 503870 205760
rect 297266 205640 297272 205692
rect 297324 205680 297330 205692
rect 297818 205680 297824 205692
rect 297324 205652 297824 205680
rect 297324 205640 297330 205652
rect 297818 205640 297824 205652
rect 297876 205640 297882 205692
rect 503714 205640 503720 205692
rect 503772 205680 503778 205692
rect 503990 205680 503996 205692
rect 503772 205652 503996 205680
rect 503772 205640 503778 205652
rect 503990 205640 503996 205652
rect 504048 205640 504054 205692
rect 504174 205640 504180 205692
rect 504232 205680 504238 205692
rect 504232 205652 504312 205680
rect 504232 205640 504238 205652
rect 504284 205624 504312 205652
rect 8018 205572 8024 205624
rect 8076 205612 8082 205624
rect 8076 205584 8156 205612
rect 8076 205572 8082 205584
rect 8128 205556 8156 205584
rect 308398 205572 308404 205624
rect 308456 205612 308462 205624
rect 308582 205612 308588 205624
rect 308456 205584 308588 205612
rect 308456 205572 308462 205584
rect 308582 205572 308588 205584
rect 308640 205572 308646 205624
rect 504266 205572 504272 205624
rect 504324 205572 504330 205624
rect 8110 205504 8116 205556
rect 8168 205504 8174 205556
rect 196618 205096 196624 205148
rect 196676 205136 196682 205148
rect 230566 205136 230572 205148
rect 196676 205108 230572 205136
rect 196676 205096 196682 205108
rect 230566 205096 230572 205108
rect 230624 205096 230630 205148
rect 195146 205028 195152 205080
rect 195204 205068 195210 205080
rect 229554 205068 229560 205080
rect 195204 205040 229560 205068
rect 195204 205028 195210 205040
rect 229554 205028 229560 205040
rect 229612 205028 229618 205080
rect 195238 204960 195244 205012
rect 195296 205000 195302 205012
rect 231210 205000 231216 205012
rect 195296 204972 231216 205000
rect 195296 204960 195302 204972
rect 231210 204960 231216 204972
rect 231268 204960 231274 205012
rect 294874 204960 294880 205012
rect 294932 205000 294938 205012
rect 378318 205000 378324 205012
rect 294932 204972 378324 205000
rect 294932 204960 294938 204972
rect 378318 204960 378324 204972
rect 378376 204960 378382 205012
rect 196526 204892 196532 204944
rect 196584 204932 196590 204944
rect 233234 204932 233240 204944
rect 196584 204904 233240 204932
rect 196584 204892 196590 204904
rect 233234 204892 233240 204904
rect 233292 204892 233298 204944
rect 237466 204892 237472 204944
rect 237524 204932 237530 204944
rect 237742 204932 237748 204944
rect 237524 204904 237748 204932
rect 237524 204892 237530 204904
rect 237742 204892 237748 204904
rect 237800 204892 237806 204944
rect 286226 204892 286232 204944
rect 286284 204932 286290 204944
rect 378226 204932 378232 204944
rect 286284 204904 378232 204932
rect 286284 204892 286290 204904
rect 378226 204892 378232 204904
rect 378284 204892 378290 204944
rect 199470 204212 199476 204264
rect 199528 204252 199534 204264
rect 244734 204252 244740 204264
rect 199528 204224 244740 204252
rect 199528 204212 199534 204224
rect 244734 204212 244740 204224
rect 244792 204212 244798 204264
rect 255774 204212 255780 204264
rect 255832 204252 255838 204264
rect 266906 204252 266912 204264
rect 255832 204224 266912 204252
rect 255832 204212 255838 204224
rect 266906 204212 266912 204224
rect 266964 204212 266970 204264
rect 319162 204212 319168 204264
rect 319220 204252 319226 204264
rect 380066 204252 380072 204264
rect 319220 204224 380072 204252
rect 319220 204212 319226 204224
rect 380066 204212 380072 204224
rect 380124 204212 380130 204264
rect 197630 204144 197636 204196
rect 197688 204184 197694 204196
rect 245654 204184 245660 204196
rect 197688 204156 245660 204184
rect 197688 204144 197694 204156
rect 245654 204144 245660 204156
rect 245712 204144 245718 204196
rect 250530 204144 250536 204196
rect 250588 204184 250594 204196
rect 267826 204184 267832 204196
rect 250588 204156 267832 204184
rect 250588 204144 250594 204156
rect 267826 204144 267832 204156
rect 267884 204144 267890 204196
rect 313550 204144 313556 204196
rect 313608 204184 313614 204196
rect 378134 204184 378140 204196
rect 313608 204156 378140 204184
rect 313608 204144 313614 204156
rect 378134 204144 378140 204156
rect 378192 204144 378198 204196
rect 197446 204076 197452 204128
rect 197504 204116 197510 204128
rect 251910 204116 251916 204128
rect 197504 204088 251916 204116
rect 197504 204076 197510 204088
rect 251910 204076 251916 204088
rect 251968 204076 251974 204128
rect 253566 204076 253572 204128
rect 253624 204116 253630 204128
rect 268654 204116 268660 204128
rect 253624 204088 268660 204116
rect 253624 204076 253630 204088
rect 268654 204076 268660 204088
rect 268712 204076 268718 204128
rect 314930 204076 314936 204128
rect 314988 204116 314994 204128
rect 380158 204116 380164 204128
rect 314988 204088 380164 204116
rect 314988 204076 314994 204088
rect 380158 204076 380164 204088
rect 380216 204076 380222 204128
rect 199378 204008 199384 204060
rect 199436 204048 199442 204060
rect 254026 204048 254032 204060
rect 199436 204020 254032 204048
rect 199436 204008 199442 204020
rect 254026 204008 254032 204020
rect 254084 204008 254090 204060
rect 255958 204008 255964 204060
rect 256016 204048 256022 204060
rect 268378 204048 268384 204060
rect 256016 204020 268384 204048
rect 256016 204008 256022 204020
rect 268378 204008 268384 204020
rect 268436 204008 268442 204060
rect 308398 204008 308404 204060
rect 308456 204048 308462 204060
rect 377214 204048 377220 204060
rect 308456 204020 377220 204048
rect 308456 204008 308462 204020
rect 377214 204008 377220 204020
rect 377272 204008 377278 204060
rect 199194 203940 199200 203992
rect 199252 203980 199258 203992
rect 258442 203980 258448 203992
rect 199252 203952 258448 203980
rect 199252 203940 199258 203952
rect 258442 203940 258448 203952
rect 258500 203940 258506 203992
rect 306650 203940 306656 203992
rect 306708 203980 306714 203992
rect 380710 203980 380716 203992
rect 306708 203952 380716 203980
rect 306708 203940 306714 203952
rect 380710 203940 380716 203952
rect 380768 203940 380774 203992
rect 197722 203872 197728 203924
rect 197780 203912 197786 203924
rect 257154 203912 257160 203924
rect 197780 203884 257160 203912
rect 197780 203872 197786 203884
rect 257154 203872 257160 203884
rect 257212 203872 257218 203924
rect 259822 203872 259828 203924
rect 259880 203912 259886 203924
rect 267182 203912 267188 203924
rect 259880 203884 267188 203912
rect 259880 203872 259886 203884
rect 267182 203872 267188 203884
rect 267240 203872 267246 203924
rect 301406 203872 301412 203924
rect 301464 203912 301470 203924
rect 379514 203912 379520 203924
rect 301464 203884 379520 203912
rect 301464 203872 301470 203884
rect 379514 203872 379520 203884
rect 379572 203872 379578 203924
rect 197906 203804 197912 203856
rect 197964 203844 197970 203856
rect 260374 203844 260380 203856
rect 197964 203816 260380 203844
rect 197964 203804 197970 203816
rect 260374 203804 260380 203816
rect 260432 203804 260438 203856
rect 299382 203804 299388 203856
rect 299440 203844 299446 203856
rect 380250 203844 380256 203856
rect 299440 203816 380256 203844
rect 299440 203804 299446 203816
rect 380250 203804 380256 203816
rect 380308 203804 380314 203856
rect 198182 203736 198188 203788
rect 198240 203776 198246 203788
rect 262766 203776 262772 203788
rect 198240 203748 262772 203776
rect 198240 203736 198246 203748
rect 262766 203736 262772 203748
rect 262824 203736 262830 203788
rect 292482 203736 292488 203788
rect 292540 203776 292546 203788
rect 379790 203776 379796 203788
rect 292540 203748 379796 203776
rect 292540 203736 292546 203748
rect 379790 203736 379796 203748
rect 379848 203736 379854 203788
rect 197538 203668 197544 203720
rect 197596 203708 197602 203720
rect 262950 203708 262956 203720
rect 197596 203680 262956 203708
rect 197596 203668 197602 203680
rect 262950 203668 262956 203680
rect 263008 203668 263014 203720
rect 287514 203668 287520 203720
rect 287572 203708 287578 203720
rect 379606 203708 379612 203720
rect 287572 203680 379612 203708
rect 287572 203668 287578 203680
rect 379606 203668 379612 203680
rect 379664 203668 379670 203720
rect 197814 203600 197820 203652
rect 197872 203640 197878 203652
rect 265434 203640 265440 203652
rect 197872 203612 265440 203640
rect 197872 203600 197878 203612
rect 265434 203600 265440 203612
rect 265492 203600 265498 203652
rect 271782 203600 271788 203652
rect 271840 203640 271846 203652
rect 369854 203640 369860 203652
rect 271840 203612 369860 203640
rect 271840 203600 271846 203612
rect 369854 203600 369860 203612
rect 369912 203600 369918 203652
rect 197998 203532 198004 203584
rect 198056 203572 198062 203584
rect 267182 203572 267188 203584
rect 198056 203544 267188 203572
rect 198056 203532 198062 203544
rect 267182 203532 267188 203544
rect 267240 203532 267246 203584
rect 280522 203532 280528 203584
rect 280580 203572 280586 203584
rect 379882 203572 379888 203584
rect 280580 203544 379888 203572
rect 280580 203532 280586 203544
rect 379882 203532 379888 203544
rect 379940 203532 379946 203584
rect 198090 203464 198096 203516
rect 198148 203504 198154 203516
rect 238754 203504 238760 203516
rect 198148 203476 238760 203504
rect 198148 203464 198154 203476
rect 238754 203464 238760 203476
rect 238812 203464 238818 203516
rect 240962 203464 240968 203516
rect 241020 203504 241026 203516
rect 268562 203504 268568 203516
rect 241020 203476 268568 203504
rect 241020 203464 241026 203476
rect 268562 203464 268568 203476
rect 268620 203464 268626 203516
rect 296162 203464 296168 203516
rect 296220 203504 296226 203516
rect 353294 203504 353300 203516
rect 296220 203476 353300 203504
rect 296220 203464 296226 203476
rect 353294 203464 353300 203476
rect 353352 203464 353358 203516
rect 209682 203396 209688 203448
rect 209740 203436 209746 203448
rect 243170 203436 243176 203448
rect 209740 203408 243176 203436
rect 209740 203396 209746 203408
rect 243170 203396 243176 203408
rect 243228 203396 243234 203448
rect 294414 203396 294420 203448
rect 294472 203436 294478 203448
rect 340874 203436 340880 203448
rect 294472 203408 340880 203436
rect 294472 203396 294478 203408
rect 340874 203396 340880 203408
rect 340932 203396 340938 203448
rect 198366 203328 198372 203380
rect 198424 203368 198430 203380
rect 225138 203368 225144 203380
rect 198424 203340 225144 203368
rect 198424 203328 198430 203340
rect 225138 203328 225144 203340
rect 225196 203328 225202 203380
rect 302878 203328 302884 203380
rect 302936 203368 302942 203380
rect 331214 203368 331220 203380
rect 302936 203340 331220 203368
rect 302936 203328 302942 203340
rect 331214 203328 331220 203340
rect 331272 203328 331278 203380
rect 297910 203260 297916 203312
rect 297968 203300 297974 203312
rect 325142 203300 325148 203312
rect 297968 203272 325148 203300
rect 297968 203260 297974 203272
rect 325142 203260 325148 203272
rect 325200 203260 325206 203312
rect 315206 203192 315212 203244
rect 315264 203232 315270 203244
rect 335998 203232 336004 203244
rect 315264 203204 336004 203232
rect 315264 203192 315270 203204
rect 335998 203192 336004 203204
rect 336056 203192 336062 203244
rect 308950 203124 308956 203176
rect 309008 203164 309014 203176
rect 321738 203164 321744 203176
rect 309008 203136 321744 203164
rect 309008 203124 309014 203136
rect 321738 203124 321744 203136
rect 321796 203124 321802 203176
rect 128446 202852 128452 202904
rect 128504 202892 128510 202904
rect 128630 202892 128636 202904
rect 128504 202864 128636 202892
rect 128504 202852 128510 202864
rect 128630 202852 128636 202864
rect 128688 202852 128694 202904
rect 258810 202892 258816 202904
rect 258552 202864 258816 202892
rect 196710 202784 196716 202836
rect 196768 202824 196774 202836
rect 196768 202796 220768 202824
rect 196768 202784 196774 202796
rect 195330 202716 195336 202768
rect 195388 202756 195394 202768
rect 220630 202756 220636 202768
rect 195388 202728 220636 202756
rect 195388 202716 195394 202728
rect 220630 202716 220636 202728
rect 220688 202716 220694 202768
rect 220740 202756 220768 202796
rect 220814 202784 220820 202836
rect 220872 202824 220878 202836
rect 221274 202824 221280 202836
rect 220872 202796 221280 202824
rect 220872 202784 220878 202796
rect 221274 202784 221280 202796
rect 221332 202784 221338 202836
rect 239674 202784 239680 202836
rect 239732 202824 239738 202836
rect 240134 202824 240140 202836
rect 239732 202796 240140 202824
rect 239732 202784 239738 202796
rect 240134 202784 240140 202796
rect 240192 202784 240198 202836
rect 240502 202784 240508 202836
rect 240560 202824 240566 202836
rect 242158 202824 242164 202836
rect 240560 202796 242164 202824
rect 240560 202784 240566 202796
rect 242158 202784 242164 202796
rect 242216 202784 242222 202836
rect 242250 202784 242256 202836
rect 242308 202824 242314 202836
rect 242802 202824 242808 202836
rect 242308 202796 242808 202824
rect 242308 202784 242314 202796
rect 242802 202784 242808 202796
rect 242860 202784 242866 202836
rect 251450 202784 251456 202836
rect 251508 202824 251514 202836
rect 258552 202824 258580 202864
rect 258810 202852 258816 202864
rect 258868 202852 258874 202904
rect 504174 202852 504180 202904
rect 504232 202892 504238 202904
rect 504266 202892 504272 202904
rect 504232 202864 504272 202892
rect 504232 202852 504238 202864
rect 504266 202852 504272 202864
rect 504324 202852 504330 202904
rect 258994 202824 259000 202836
rect 251508 202796 258580 202824
rect 258644 202796 259000 202824
rect 251508 202784 251514 202796
rect 226886 202756 226892 202768
rect 220740 202728 226892 202756
rect 226886 202716 226892 202728
rect 226944 202716 226950 202768
rect 236362 202716 236368 202768
rect 236420 202756 236426 202768
rect 258644 202756 258672 202796
rect 258994 202784 259000 202796
rect 259052 202784 259058 202836
rect 260098 202784 260104 202836
rect 260156 202824 260162 202836
rect 263594 202824 263600 202836
rect 260156 202796 263600 202824
rect 260156 202784 260162 202796
rect 263594 202784 263600 202796
rect 263652 202784 263658 202836
rect 266262 202784 266268 202836
rect 266320 202824 266326 202836
rect 269390 202824 269396 202836
rect 266320 202796 269396 202824
rect 266320 202784 266326 202796
rect 269390 202784 269396 202796
rect 269448 202784 269454 202836
rect 289262 202784 289268 202836
rect 289320 202824 289326 202836
rect 289722 202824 289728 202836
rect 289320 202796 289728 202824
rect 289320 202784 289326 202796
rect 289722 202784 289728 202796
rect 289780 202784 289786 202836
rect 290550 202784 290556 202836
rect 290608 202824 290614 202836
rect 291010 202824 291016 202836
rect 290608 202796 291016 202824
rect 290608 202784 290614 202796
rect 291010 202784 291016 202796
rect 291068 202784 291074 202836
rect 291378 202784 291384 202836
rect 291436 202824 291442 202836
rect 292390 202824 292396 202836
rect 291436 202796 292396 202824
rect 291436 202784 291442 202796
rect 292390 202784 292396 202796
rect 292448 202784 292454 202836
rect 293126 202784 293132 202836
rect 293184 202824 293190 202836
rect 293862 202824 293868 202836
rect 293184 202796 293868 202824
rect 293184 202784 293190 202796
rect 293862 202784 293868 202796
rect 293920 202784 293926 202836
rect 295794 202784 295800 202836
rect 295852 202824 295858 202836
rect 296438 202824 296444 202836
rect 295852 202796 296444 202824
rect 295852 202784 295858 202796
rect 296438 202784 296444 202796
rect 296496 202784 296502 202836
rect 300118 202784 300124 202836
rect 300176 202824 300182 202836
rect 300670 202824 300676 202836
rect 300176 202796 300676 202824
rect 300176 202784 300182 202796
rect 300670 202784 300676 202796
rect 300728 202784 300734 202836
rect 307110 202824 307116 202836
rect 300964 202796 307116 202824
rect 236420 202728 258672 202756
rect 236420 202716 236426 202728
rect 258718 202716 258724 202768
rect 258776 202756 258782 202768
rect 263870 202756 263876 202768
rect 258776 202728 263876 202756
rect 258776 202716 258782 202728
rect 263870 202716 263876 202728
rect 263928 202716 263934 202768
rect 264882 202716 264888 202768
rect 264940 202756 264946 202768
rect 269482 202756 269488 202768
rect 264940 202728 269488 202756
rect 264940 202716 264946 202728
rect 269482 202716 269488 202728
rect 269540 202716 269546 202768
rect 299474 202716 299480 202768
rect 299532 202756 299538 202768
rect 300964 202756 300992 202796
rect 307110 202784 307116 202796
rect 307168 202784 307174 202836
rect 311894 202784 311900 202836
rect 311952 202824 311958 202836
rect 312538 202824 312544 202836
rect 311952 202796 312544 202824
rect 311952 202784 311958 202796
rect 312538 202784 312544 202796
rect 312596 202784 312602 202836
rect 312630 202784 312636 202836
rect 312688 202824 312694 202836
rect 319162 202824 319168 202836
rect 312688 202796 319168 202824
rect 312688 202784 312694 202796
rect 319162 202784 319168 202796
rect 319220 202784 319226 202836
rect 319254 202784 319260 202836
rect 319312 202824 319318 202836
rect 320082 202824 320088 202836
rect 319312 202796 320088 202824
rect 319312 202784 319318 202796
rect 320082 202784 320088 202796
rect 320140 202784 320146 202836
rect 350994 202784 351000 202836
rect 351052 202824 351058 202836
rect 351822 202824 351828 202836
rect 351052 202796 351828 202824
rect 351052 202784 351058 202796
rect 351822 202784 351828 202796
rect 351880 202784 351886 202836
rect 352742 202784 352748 202836
rect 352800 202824 352806 202836
rect 353202 202824 353208 202836
rect 352800 202796 353208 202824
rect 352800 202784 352806 202796
rect 353202 202784 353208 202796
rect 353260 202784 353266 202836
rect 353294 202784 353300 202836
rect 353352 202824 353358 202836
rect 413002 202824 413008 202836
rect 353352 202796 413008 202824
rect 353352 202784 353358 202796
rect 413002 202784 413008 202796
rect 413060 202784 413066 202836
rect 413094 202784 413100 202836
rect 413152 202824 413158 202836
rect 414658 202824 414664 202836
rect 413152 202796 414664 202824
rect 413152 202784 413158 202796
rect 414658 202784 414664 202796
rect 414716 202784 414722 202836
rect 415026 202784 415032 202836
rect 415084 202824 415090 202836
rect 417418 202824 417424 202836
rect 415084 202796 417424 202824
rect 415084 202784 415090 202796
rect 417418 202784 417424 202796
rect 417476 202784 417482 202836
rect 417510 202784 417516 202836
rect 417568 202824 417574 202836
rect 418062 202824 418068 202836
rect 417568 202796 418068 202824
rect 417568 202784 417574 202796
rect 418062 202784 418068 202796
rect 418120 202784 418126 202836
rect 299532 202728 300992 202756
rect 299532 202716 299538 202728
rect 301038 202716 301044 202768
rect 301096 202756 301102 202768
rect 307202 202756 307208 202768
rect 301096 202728 307208 202756
rect 301096 202716 301102 202728
rect 307202 202716 307208 202728
rect 307260 202716 307266 202768
rect 310422 202716 310428 202768
rect 310480 202756 310486 202768
rect 375650 202756 375656 202768
rect 310480 202728 375656 202756
rect 310480 202716 310486 202728
rect 375650 202716 375656 202728
rect 375708 202716 375714 202768
rect 375742 202716 375748 202768
rect 375800 202756 375806 202768
rect 378778 202756 378784 202768
rect 375800 202728 378784 202756
rect 375800 202716 375806 202728
rect 378778 202716 378784 202728
rect 378836 202716 378842 202768
rect 400582 202716 400588 202768
rect 400640 202756 400646 202768
rect 401502 202756 401508 202768
rect 400640 202728 401508 202756
rect 400640 202716 400646 202728
rect 401502 202716 401508 202728
rect 401560 202716 401566 202768
rect 401594 202716 401600 202768
rect 401652 202756 401658 202768
rect 458818 202756 458824 202768
rect 401652 202728 458824 202756
rect 401652 202716 401658 202728
rect 458818 202716 458824 202728
rect 458876 202716 458882 202768
rect 200022 202648 200028 202700
rect 200080 202688 200086 202700
rect 238202 202688 238208 202700
rect 200080 202660 238208 202688
rect 200080 202648 200086 202660
rect 238202 202648 238208 202660
rect 238260 202648 238266 202700
rect 240778 202648 240784 202700
rect 240836 202688 240842 202700
rect 242342 202688 242348 202700
rect 240836 202660 242348 202688
rect 240836 202648 240842 202660
rect 242342 202648 242348 202660
rect 242400 202648 242406 202700
rect 250898 202648 250904 202700
rect 250956 202688 250962 202700
rect 269206 202688 269212 202700
rect 250956 202660 269212 202688
rect 250956 202648 250962 202660
rect 269206 202648 269212 202660
rect 269264 202648 269270 202700
rect 299106 202648 299112 202700
rect 299164 202688 299170 202700
rect 304994 202688 305000 202700
rect 299164 202660 305000 202688
rect 299164 202648 299170 202660
rect 304994 202648 305000 202660
rect 305052 202648 305058 202700
rect 306926 202648 306932 202700
rect 306984 202688 306990 202700
rect 320634 202688 320640 202700
rect 306984 202660 320640 202688
rect 306984 202648 306990 202660
rect 320634 202648 320640 202660
rect 320692 202648 320698 202700
rect 344002 202648 344008 202700
rect 344060 202688 344066 202700
rect 344060 202660 347820 202688
rect 344060 202648 344066 202660
rect 156598 202580 156604 202632
rect 156656 202620 156662 202632
rect 169110 202620 169116 202632
rect 156656 202592 169116 202620
rect 156656 202580 156662 202592
rect 169110 202580 169116 202592
rect 169168 202580 169174 202632
rect 198274 202580 198280 202632
rect 198332 202620 198338 202632
rect 202874 202620 202880 202632
rect 198332 202592 202880 202620
rect 198332 202580 198338 202592
rect 202874 202580 202880 202592
rect 202932 202580 202938 202632
rect 207658 202580 207664 202632
rect 207716 202620 207722 202632
rect 239306 202620 239312 202632
rect 207716 202592 239312 202620
rect 207716 202580 207722 202592
rect 239306 202580 239312 202592
rect 239364 202580 239370 202632
rect 239398 202580 239404 202632
rect 239456 202620 239462 202632
rect 243814 202620 243820 202632
rect 239456 202592 243820 202620
rect 239456 202580 239462 202592
rect 243814 202580 243820 202592
rect 243872 202580 243878 202632
rect 248966 202580 248972 202632
rect 249024 202620 249030 202632
rect 268102 202620 268108 202632
rect 249024 202592 268108 202620
rect 249024 202580 249030 202592
rect 268102 202580 268108 202592
rect 268160 202580 268166 202632
rect 283926 202580 283932 202632
rect 283984 202620 283990 202632
rect 284202 202620 284208 202632
rect 283984 202592 284208 202620
rect 283984 202580 283990 202592
rect 284202 202580 284208 202592
rect 284260 202580 284266 202632
rect 299014 202580 299020 202632
rect 299072 202620 299078 202632
rect 305638 202620 305644 202632
rect 299072 202592 305644 202620
rect 299072 202580 299078 202592
rect 305638 202580 305644 202592
rect 305696 202580 305702 202632
rect 307202 202580 307208 202632
rect 307260 202620 307266 202632
rect 309502 202620 309508 202632
rect 307260 202592 309508 202620
rect 307260 202580 307266 202592
rect 309502 202580 309508 202592
rect 309560 202580 309566 202632
rect 311158 202580 311164 202632
rect 311216 202620 311222 202632
rect 331858 202620 331864 202632
rect 311216 202592 331864 202620
rect 311216 202580 311222 202592
rect 331858 202580 331864 202592
rect 331916 202580 331922 202632
rect 342070 202580 342076 202632
rect 342128 202620 342134 202632
rect 342128 202592 347728 202620
rect 342128 202580 342134 202592
rect 153838 202512 153844 202564
rect 153896 202552 153902 202564
rect 178034 202552 178040 202564
rect 153896 202524 178040 202552
rect 153896 202512 153902 202524
rect 178034 202512 178040 202524
rect 178092 202512 178098 202564
rect 196986 202512 196992 202564
rect 197044 202552 197050 202564
rect 241514 202552 241520 202564
rect 197044 202524 241520 202552
rect 197044 202512 197050 202524
rect 241514 202512 241520 202524
rect 241572 202512 241578 202564
rect 247494 202512 247500 202564
rect 247552 202552 247558 202564
rect 247552 202524 253796 202552
rect 247552 202512 247558 202524
rect 130102 202444 130108 202496
rect 130160 202484 130166 202496
rect 134426 202484 134432 202496
rect 130160 202456 134432 202484
rect 130160 202444 130166 202456
rect 134426 202444 134432 202456
rect 134484 202444 134490 202496
rect 152458 202444 152464 202496
rect 152516 202484 152522 202496
rect 176930 202484 176936 202496
rect 152516 202456 176936 202484
rect 152516 202444 152522 202456
rect 176930 202444 176936 202456
rect 176988 202444 176994 202496
rect 195514 202444 195520 202496
rect 195572 202484 195578 202496
rect 241054 202484 241060 202496
rect 195572 202456 241060 202484
rect 195572 202444 195578 202456
rect 241054 202444 241060 202456
rect 241112 202444 241118 202496
rect 243722 202444 243728 202496
rect 243780 202484 243786 202496
rect 252646 202484 252652 202496
rect 243780 202456 252652 202484
rect 243780 202444 243786 202456
rect 252646 202444 252652 202456
rect 252704 202444 252710 202496
rect 253768 202484 253796 202524
rect 253842 202512 253848 202564
rect 253900 202552 253906 202564
rect 267918 202552 267924 202564
rect 253900 202524 267924 202552
rect 253900 202512 253906 202524
rect 267918 202512 267924 202524
rect 267976 202512 267982 202564
rect 299290 202512 299296 202564
rect 299348 202552 299354 202564
rect 302234 202552 302240 202564
rect 299348 202524 302240 202552
rect 299348 202512 299354 202524
rect 302234 202512 302240 202524
rect 302292 202512 302298 202564
rect 302326 202512 302332 202564
rect 302384 202552 302390 202564
rect 302970 202552 302976 202564
rect 302384 202524 302976 202552
rect 302384 202512 302390 202524
rect 302970 202512 302976 202524
rect 303028 202512 303034 202564
rect 307294 202512 307300 202564
rect 307352 202552 307358 202564
rect 325694 202552 325700 202564
rect 307352 202524 325700 202552
rect 307352 202512 307358 202524
rect 325694 202512 325700 202524
rect 325752 202512 325758 202564
rect 253768 202456 253888 202484
rect 151078 202376 151084 202428
rect 151136 202416 151142 202428
rect 182174 202416 182180 202428
rect 151136 202388 182180 202416
rect 151136 202376 151142 202388
rect 182174 202376 182180 202388
rect 182232 202376 182238 202428
rect 199930 202376 199936 202428
rect 199988 202416 199994 202428
rect 246482 202416 246488 202428
rect 199988 202388 246488 202416
rect 199988 202376 199994 202388
rect 246482 202376 246488 202388
rect 246540 202376 246546 202428
rect 137278 202308 137284 202360
rect 137336 202348 137342 202360
rect 168374 202348 168380 202360
rect 137336 202320 168380 202348
rect 137336 202308 137342 202320
rect 168374 202308 168380 202320
rect 168432 202308 168438 202360
rect 195606 202308 195612 202360
rect 195664 202348 195670 202360
rect 245194 202348 245200 202360
rect 195664 202320 245200 202348
rect 195664 202308 195670 202320
rect 245194 202308 245200 202320
rect 245252 202308 245258 202360
rect 247586 202308 247592 202360
rect 247644 202348 247650 202360
rect 253474 202348 253480 202360
rect 247644 202320 253480 202348
rect 247644 202308 247650 202320
rect 253474 202308 253480 202320
rect 253532 202308 253538 202360
rect 253860 202348 253888 202456
rect 254118 202444 254124 202496
rect 254176 202484 254182 202496
rect 266262 202484 266268 202496
rect 254176 202456 266268 202484
rect 254176 202444 254182 202456
rect 266262 202444 266268 202456
rect 266320 202444 266326 202496
rect 267642 202444 267648 202496
rect 267700 202484 267706 202496
rect 269298 202484 269304 202496
rect 267700 202456 269304 202484
rect 267700 202444 267706 202456
rect 269298 202444 269304 202456
rect 269356 202444 269362 202496
rect 273990 202444 273996 202496
rect 274048 202484 274054 202496
rect 274542 202484 274548 202496
rect 274048 202456 274548 202484
rect 274048 202444 274054 202456
rect 274542 202444 274548 202456
rect 274600 202444 274606 202496
rect 280982 202444 280988 202496
rect 281040 202484 281046 202496
rect 281258 202484 281264 202496
rect 281040 202456 281264 202484
rect 281040 202444 281046 202456
rect 281258 202444 281264 202456
rect 281316 202444 281322 202496
rect 282270 202444 282276 202496
rect 282328 202484 282334 202496
rect 282730 202484 282736 202496
rect 282328 202456 282736 202484
rect 282328 202444 282334 202456
rect 282730 202444 282736 202456
rect 282788 202444 282794 202496
rect 288802 202444 288808 202496
rect 288860 202484 288866 202496
rect 315298 202484 315304 202496
rect 288860 202456 315304 202484
rect 288860 202444 288866 202456
rect 315298 202444 315304 202456
rect 315356 202444 315362 202496
rect 333146 202444 333152 202496
rect 333204 202484 333210 202496
rect 333882 202484 333888 202496
rect 333204 202456 333888 202484
rect 333204 202444 333210 202456
rect 333882 202444 333888 202456
rect 333940 202444 333946 202496
rect 341426 202444 341432 202496
rect 341484 202484 341490 202496
rect 342162 202484 342168 202496
rect 341484 202456 342168 202484
rect 341484 202444 341490 202456
rect 342162 202444 342168 202456
rect 342220 202444 342226 202496
rect 343174 202444 343180 202496
rect 343232 202484 343238 202496
rect 343542 202484 343548 202496
rect 343232 202456 343548 202484
rect 343232 202444 343238 202456
rect 343542 202444 343548 202456
rect 343600 202444 343606 202496
rect 346670 202444 346676 202496
rect 346728 202484 346734 202496
rect 347590 202484 347596 202496
rect 346728 202456 347596 202484
rect 346728 202444 346734 202456
rect 347590 202444 347596 202456
rect 347648 202444 347654 202496
rect 347700 202484 347728 202592
rect 347792 202552 347820 202660
rect 349982 202648 349988 202700
rect 350040 202688 350046 202700
rect 350442 202688 350448 202700
rect 350040 202660 350448 202688
rect 350040 202648 350046 202660
rect 350442 202648 350448 202660
rect 350500 202648 350506 202700
rect 351730 202648 351736 202700
rect 351788 202688 351794 202700
rect 353294 202688 353300 202700
rect 351788 202660 353300 202688
rect 351788 202648 351794 202660
rect 353294 202648 353300 202660
rect 353352 202648 353358 202700
rect 412910 202688 412916 202700
rect 353404 202660 412916 202688
rect 348326 202580 348332 202632
rect 348384 202620 348390 202632
rect 353404 202620 353432 202660
rect 412910 202648 412916 202660
rect 412968 202648 412974 202700
rect 413002 202648 413008 202700
rect 413060 202688 413066 202700
rect 417326 202688 417332 202700
rect 413060 202660 417332 202688
rect 413060 202648 413066 202660
rect 417326 202648 417332 202660
rect 417384 202648 417390 202700
rect 348384 202592 353432 202620
rect 348384 202580 348390 202592
rect 353478 202580 353484 202632
rect 353536 202620 353542 202632
rect 417142 202620 417148 202632
rect 353536 202592 417148 202620
rect 353536 202580 353542 202592
rect 417142 202580 417148 202592
rect 417200 202580 417206 202632
rect 416866 202552 416872 202564
rect 347792 202524 416872 202552
rect 416866 202512 416872 202524
rect 416924 202512 416930 202564
rect 412818 202484 412824 202496
rect 347700 202456 412824 202484
rect 412818 202444 412824 202456
rect 412876 202444 412882 202496
rect 412910 202444 412916 202496
rect 412968 202484 412974 202496
rect 417234 202484 417240 202496
rect 412968 202456 417240 202484
rect 412968 202444 412974 202456
rect 417234 202444 417240 202456
rect 417292 202444 417298 202496
rect 253934 202376 253940 202428
rect 253992 202416 253998 202428
rect 268010 202416 268016 202428
rect 253992 202388 268016 202416
rect 253992 202376 253998 202388
rect 268010 202376 268016 202388
rect 268068 202376 268074 202428
rect 299198 202376 299204 202428
rect 299256 202416 299262 202428
rect 306926 202416 306932 202428
rect 299256 202388 306932 202416
rect 299256 202376 299262 202388
rect 306926 202376 306932 202388
rect 306984 202376 306990 202428
rect 307018 202376 307024 202428
rect 307076 202416 307082 202428
rect 307570 202416 307576 202428
rect 307076 202388 307576 202416
rect 307076 202376 307082 202388
rect 307570 202376 307576 202388
rect 307628 202376 307634 202428
rect 310514 202376 310520 202428
rect 310572 202416 310578 202428
rect 311250 202416 311256 202428
rect 310572 202388 311256 202416
rect 310572 202376 310578 202388
rect 311250 202376 311256 202388
rect 311308 202376 311314 202428
rect 311342 202376 311348 202428
rect 311400 202416 311406 202428
rect 325694 202416 325700 202428
rect 311400 202388 325700 202416
rect 311400 202376 311406 202388
rect 325694 202376 325700 202388
rect 325752 202376 325758 202428
rect 332502 202376 332508 202428
rect 332560 202416 332566 202428
rect 415026 202416 415032 202428
rect 332560 202388 415032 202416
rect 332560 202376 332566 202388
rect 415026 202376 415032 202388
rect 415084 202376 415090 202428
rect 415762 202376 415768 202428
rect 415820 202416 415826 202428
rect 416682 202416 416688 202428
rect 415820 202388 416688 202416
rect 415820 202376 415826 202388
rect 416682 202376 416688 202388
rect 416740 202376 416746 202428
rect 266078 202348 266084 202360
rect 253860 202320 266084 202348
rect 266078 202308 266084 202320
rect 266136 202308 266142 202360
rect 266170 202308 266176 202360
rect 266228 202348 266234 202360
rect 269574 202348 269580 202360
rect 266228 202320 269580 202348
rect 266228 202308 266234 202320
rect 269574 202308 269580 202320
rect 269632 202308 269638 202360
rect 297542 202308 297548 202360
rect 297600 202348 297606 202360
rect 302234 202348 302240 202360
rect 297600 202320 302240 202348
rect 297600 202308 297606 202320
rect 302234 202308 302240 202320
rect 302292 202308 302298 202360
rect 305546 202308 305552 202360
rect 305604 202348 305610 202360
rect 305604 202320 375604 202348
rect 305604 202308 305610 202320
rect 140038 202240 140044 202292
rect 140096 202280 140102 202292
rect 178678 202280 178684 202292
rect 140096 202252 178684 202280
rect 140096 202240 140102 202252
rect 178678 202240 178684 202252
rect 178736 202240 178742 202292
rect 201402 202240 201408 202292
rect 201460 202280 201466 202292
rect 258534 202280 258540 202292
rect 201460 202252 258540 202280
rect 201460 202240 201466 202252
rect 258534 202240 258540 202252
rect 258592 202240 258598 202292
rect 269758 202280 269764 202292
rect 258828 202252 269764 202280
rect 103422 202172 103428 202224
rect 103480 202212 103486 202224
rect 142522 202212 142528 202224
rect 103480 202184 142528 202212
rect 103480 202172 103486 202184
rect 142522 202172 142528 202184
rect 142580 202172 142586 202224
rect 144178 202172 144184 202224
rect 144236 202212 144242 202224
rect 181254 202212 181260 202224
rect 144236 202184 181260 202212
rect 144236 202172 144242 202184
rect 181254 202172 181260 202184
rect 181312 202172 181318 202224
rect 199102 202172 199108 202224
rect 199160 202212 199166 202224
rect 256510 202212 256516 202224
rect 199160 202184 256516 202212
rect 199160 202172 199166 202184
rect 256510 202172 256516 202184
rect 256568 202172 256574 202224
rect 93762 202104 93768 202156
rect 93820 202144 93826 202156
rect 134702 202144 134708 202156
rect 93820 202116 134708 202144
rect 93820 202104 93826 202116
rect 134702 202104 134708 202116
rect 134760 202104 134766 202156
rect 141418 202104 141424 202156
rect 141476 202144 141482 202156
rect 180334 202144 180340 202156
rect 141476 202116 180340 202144
rect 141476 202104 141482 202116
rect 180334 202104 180340 202116
rect 180392 202104 180398 202156
rect 199286 202104 199292 202156
rect 199344 202144 199350 202156
rect 258828 202144 258856 202252
rect 269758 202240 269764 202252
rect 269816 202240 269822 202292
rect 292298 202240 292304 202292
rect 292356 202280 292362 202292
rect 375576 202280 375604 202320
rect 375650 202308 375656 202360
rect 375708 202348 375714 202360
rect 377306 202348 377312 202360
rect 375708 202320 377312 202348
rect 375708 202308 375714 202320
rect 377306 202308 377312 202320
rect 377364 202308 377370 202360
rect 410150 202308 410156 202360
rect 410208 202348 410214 202360
rect 411162 202348 411168 202360
rect 410208 202320 411168 202348
rect 410208 202308 410214 202320
rect 411162 202308 411168 202320
rect 411220 202308 411226 202360
rect 417142 202308 417148 202360
rect 417200 202348 417206 202360
rect 503898 202348 503904 202360
rect 417200 202320 503904 202348
rect 417200 202308 417206 202320
rect 503898 202308 503904 202320
rect 503956 202308 503962 202360
rect 378502 202280 378508 202292
rect 292356 202252 375512 202280
rect 375576 202252 378508 202280
rect 292356 202240 292362 202252
rect 258994 202172 259000 202224
rect 259052 202212 259058 202224
rect 266722 202212 266728 202224
rect 259052 202184 266728 202212
rect 259052 202172 259058 202184
rect 266722 202172 266728 202184
rect 266780 202172 266786 202224
rect 270954 202172 270960 202224
rect 271012 202212 271018 202224
rect 374362 202212 374368 202224
rect 271012 202184 374368 202212
rect 271012 202172 271018 202184
rect 374362 202172 374368 202184
rect 374420 202172 374426 202224
rect 374454 202172 374460 202224
rect 374512 202212 374518 202224
rect 375282 202212 375288 202224
rect 374512 202184 375288 202212
rect 374512 202172 374518 202184
rect 375282 202172 375288 202184
rect 375340 202172 375346 202224
rect 375484 202212 375512 202252
rect 378502 202240 378508 202252
rect 378560 202240 378566 202292
rect 411070 202240 411076 202292
rect 411128 202280 411134 202292
rect 503806 202280 503812 202292
rect 411128 202252 503812 202280
rect 411128 202240 411134 202252
rect 503806 202240 503812 202252
rect 503864 202240 503870 202292
rect 379698 202212 379704 202224
rect 375484 202184 379704 202212
rect 379698 202172 379704 202184
rect 379756 202172 379762 202224
rect 409230 202172 409236 202224
rect 409288 202212 409294 202224
rect 503714 202212 503720 202224
rect 409288 202184 503720 202212
rect 409288 202172 409294 202184
rect 503714 202172 503720 202184
rect 503772 202172 503778 202224
rect 199344 202116 258856 202144
rect 199344 202104 199350 202116
rect 258902 202104 258908 202156
rect 258960 202144 258966 202156
rect 268286 202144 268292 202156
rect 258960 202116 268292 202144
rect 258960 202104 258966 202116
rect 268286 202104 268292 202116
rect 268344 202104 268350 202156
rect 283558 202104 283564 202156
rect 283616 202144 283622 202156
rect 283616 202116 326384 202144
rect 283616 202104 283622 202116
rect 196894 202036 196900 202088
rect 196952 202076 196958 202088
rect 216858 202076 216864 202088
rect 196952 202048 216864 202076
rect 196952 202036 196958 202048
rect 216858 202036 216864 202048
rect 216916 202036 216922 202088
rect 217962 202036 217968 202088
rect 218020 202076 218026 202088
rect 218020 202048 239168 202076
rect 218020 202036 218026 202048
rect 195422 201968 195428 202020
rect 195480 202008 195486 202020
rect 223022 202008 223028 202020
rect 195480 201980 223028 202008
rect 195480 201968 195486 201980
rect 223022 201968 223028 201980
rect 223080 201968 223086 202020
rect 195882 201900 195888 201952
rect 195940 201940 195946 201952
rect 218054 201940 218060 201952
rect 195940 201912 218060 201940
rect 195940 201900 195946 201912
rect 218054 201900 218060 201912
rect 218112 201900 218118 201952
rect 220630 201900 220636 201952
rect 220688 201940 220694 201952
rect 227806 201940 227812 201952
rect 220688 201912 227812 201940
rect 220688 201900 220694 201912
rect 227806 201900 227812 201912
rect 227864 201900 227870 201952
rect 199654 201832 199660 201884
rect 199712 201872 199718 201884
rect 219526 201872 219532 201884
rect 199712 201844 219532 201872
rect 199712 201832 199718 201844
rect 219526 201832 219532 201844
rect 219584 201832 219590 201884
rect 196802 201764 196808 201816
rect 196860 201804 196866 201816
rect 218606 201804 218612 201816
rect 196860 201776 218612 201804
rect 196860 201764 196866 201776
rect 218606 201764 218612 201776
rect 218664 201764 218670 201816
rect 239140 201804 239168 202048
rect 239214 202036 239220 202088
rect 239272 202076 239278 202088
rect 240042 202076 240048 202088
rect 239272 202048 240048 202076
rect 239272 202036 239278 202048
rect 240042 202036 240048 202048
rect 240100 202036 240106 202088
rect 251818 202036 251824 202088
rect 251876 202076 251882 202088
rect 267734 202076 267740 202088
rect 251876 202048 267740 202076
rect 251876 202036 251882 202048
rect 267734 202036 267740 202048
rect 267792 202036 267798 202088
rect 297450 202036 297456 202088
rect 297508 202076 297514 202088
rect 303890 202076 303896 202088
rect 297508 202048 303896 202076
rect 297508 202036 297514 202048
rect 303890 202036 303896 202048
rect 303948 202036 303954 202088
rect 306926 202036 306932 202088
rect 306984 202076 306990 202088
rect 315298 202076 315304 202088
rect 306984 202048 315304 202076
rect 306984 202036 306990 202048
rect 315298 202036 315304 202048
rect 315356 202036 315362 202088
rect 246298 201968 246304 202020
rect 246356 202008 246362 202020
rect 246356 201980 248000 202008
rect 246356 201968 246362 201980
rect 243078 201900 243084 201952
rect 243136 201940 243142 201952
rect 247678 201940 247684 201952
rect 243136 201912 247684 201940
rect 243136 201900 243142 201912
rect 247678 201900 247684 201912
rect 247736 201900 247742 201952
rect 247972 201940 248000 201980
rect 253106 201968 253112 202020
rect 253164 202008 253170 202020
rect 253658 202008 253664 202020
rect 253164 201980 253664 202008
rect 253164 201968 253170 201980
rect 253658 201968 253664 201980
rect 253716 201968 253722 202020
rect 253750 201968 253756 202020
rect 253808 202008 253814 202020
rect 258718 202008 258724 202020
rect 253808 201980 258724 202008
rect 253808 201968 253814 201980
rect 258718 201968 258724 201980
rect 258776 201968 258782 202020
rect 258810 201968 258816 202020
rect 258868 202008 258874 202020
rect 266446 202008 266452 202020
rect 258868 201980 266452 202008
rect 258868 201968 258874 201980
rect 266446 201968 266452 201980
rect 266504 201968 266510 202020
rect 300486 201968 300492 202020
rect 300544 202008 300550 202020
rect 317138 202008 317144 202020
rect 300544 201980 317144 202008
rect 300544 201968 300550 201980
rect 317138 201968 317144 201980
rect 317196 201968 317202 202020
rect 320542 201968 320548 202020
rect 320600 202008 320606 202020
rect 321462 202008 321468 202020
rect 320600 201980 321468 202008
rect 320600 201968 320606 201980
rect 321462 201968 321468 201980
rect 321520 201968 321526 202020
rect 324038 201968 324044 202020
rect 324096 202008 324102 202020
rect 324958 202008 324964 202020
rect 324096 201980 324964 202008
rect 324096 201968 324102 201980
rect 324958 201968 324964 201980
rect 325016 201968 325022 202020
rect 326356 202008 326384 202116
rect 345750 202104 345756 202156
rect 345808 202144 345814 202156
rect 353478 202144 353484 202156
rect 345808 202116 353484 202144
rect 345808 202104 345814 202116
rect 353478 202104 353484 202116
rect 353536 202104 353542 202156
rect 353570 202104 353576 202156
rect 353628 202144 353634 202156
rect 354582 202144 354588 202156
rect 353628 202116 354588 202144
rect 353628 202104 353634 202116
rect 354582 202104 354588 202116
rect 354640 202104 354646 202156
rect 364886 202104 364892 202156
rect 364944 202144 364950 202156
rect 365530 202144 365536 202156
rect 364944 202116 365536 202144
rect 364944 202104 364950 202116
rect 365530 202104 365536 202116
rect 365588 202104 365594 202156
rect 366174 202104 366180 202156
rect 366232 202144 366238 202156
rect 367002 202144 367008 202156
rect 366232 202116 367008 202144
rect 366232 202104 366238 202116
rect 367002 202104 367008 202116
rect 367060 202104 367066 202156
rect 376478 202104 376484 202156
rect 376536 202144 376542 202156
rect 505738 202144 505744 202156
rect 376536 202116 505744 202144
rect 376536 202104 376542 202116
rect 505738 202104 505744 202116
rect 505796 202104 505802 202156
rect 357894 202036 357900 202088
rect 357952 202076 357958 202088
rect 357952 202048 414796 202076
rect 357952 202036 357958 202048
rect 334618 202008 334624 202020
rect 326356 201980 334624 202008
rect 334618 201968 334624 201980
rect 334676 201968 334682 202020
rect 366910 201968 366916 202020
rect 366968 202008 366974 202020
rect 414658 202008 414664 202020
rect 366968 201980 414664 202008
rect 366968 201968 366974 201980
rect 414658 201968 414664 201980
rect 414716 201968 414722 202020
rect 414768 202008 414796 202048
rect 414934 202036 414940 202088
rect 414992 202076 414998 202088
rect 417142 202076 417148 202088
rect 414992 202048 417148 202076
rect 414992 202036 414998 202048
rect 417142 202036 417148 202048
rect 417200 202036 417206 202088
rect 416958 202008 416964 202020
rect 414768 201980 416964 202008
rect 416958 201968 416964 201980
rect 417016 201968 417022 202020
rect 260834 201940 260840 201952
rect 247972 201912 260840 201940
rect 260834 201900 260840 201912
rect 260892 201900 260898 201952
rect 265342 201900 265348 201952
rect 265400 201940 265406 201952
rect 266814 201940 266820 201952
rect 265400 201912 266820 201940
rect 265400 201900 265406 201912
rect 266814 201900 266820 201912
rect 266872 201900 266878 201952
rect 266998 201900 267004 201952
rect 267056 201940 267062 201952
rect 268194 201940 268200 201952
rect 267056 201912 268200 201940
rect 267056 201900 267062 201912
rect 268194 201900 268200 201912
rect 268252 201900 268258 201952
rect 299198 201900 299204 201952
rect 299256 201940 299262 201952
rect 304258 201940 304264 201952
rect 299256 201912 304264 201940
rect 299256 201900 299262 201912
rect 304258 201900 304264 201912
rect 304316 201900 304322 201952
rect 315574 201940 315580 201952
rect 305932 201912 315580 201940
rect 239306 201832 239312 201884
rect 239364 201872 239370 201884
rect 247770 201872 247776 201884
rect 239364 201844 247776 201872
rect 239364 201832 239370 201844
rect 247770 201832 247776 201844
rect 247828 201832 247834 201884
rect 257062 201832 257068 201884
rect 257120 201872 257126 201884
rect 265986 201872 265992 201884
rect 257120 201844 265992 201872
rect 257120 201832 257126 201844
rect 265986 201832 265992 201844
rect 266044 201832 266050 201884
rect 266078 201832 266084 201884
rect 266136 201872 266142 201884
rect 270678 201872 270684 201884
rect 266136 201844 270684 201872
rect 266136 201832 266142 201844
rect 270678 201832 270684 201844
rect 270736 201832 270742 201884
rect 297266 201832 297272 201884
rect 297324 201872 297330 201884
rect 305546 201872 305552 201884
rect 297324 201844 305552 201872
rect 297324 201832 297330 201844
rect 305546 201832 305552 201844
rect 305604 201832 305610 201884
rect 246022 201804 246028 201816
rect 239140 201776 246028 201804
rect 246022 201764 246028 201776
rect 246080 201764 246086 201816
rect 256510 201764 256516 201816
rect 256568 201804 256574 201816
rect 259914 201804 259920 201816
rect 256568 201776 259920 201804
rect 256568 201764 256574 201776
rect 259914 201764 259920 201776
rect 259972 201764 259978 201816
rect 266446 201804 266452 201816
rect 260024 201776 266452 201804
rect 198734 201696 198740 201748
rect 198792 201736 198798 201748
rect 216030 201736 216036 201748
rect 198792 201708 216036 201736
rect 198792 201696 198798 201708
rect 216030 201696 216036 201708
rect 216088 201696 216094 201748
rect 250070 201696 250076 201748
rect 250128 201736 250134 201748
rect 250990 201736 250996 201748
rect 250128 201708 250996 201736
rect 250128 201696 250134 201708
rect 250990 201696 250996 201708
rect 251048 201696 251054 201748
rect 254854 201696 254860 201748
rect 254912 201736 254918 201748
rect 260024 201736 260052 201776
rect 266446 201764 266452 201776
rect 266504 201764 266510 201816
rect 270862 201804 270868 201816
rect 266786 201776 270868 201804
rect 254912 201708 260052 201736
rect 254912 201696 254918 201708
rect 262674 201696 262680 201748
rect 262732 201736 262738 201748
rect 265894 201736 265900 201748
rect 262732 201708 265900 201736
rect 262732 201696 262738 201708
rect 265894 201696 265900 201708
rect 265952 201696 265958 201748
rect 265986 201696 265992 201748
rect 266044 201736 266050 201748
rect 266786 201736 266814 201776
rect 270862 201764 270868 201776
rect 270920 201764 270926 201816
rect 300394 201764 300400 201816
rect 300452 201804 300458 201816
rect 305932 201804 305960 201912
rect 315574 201900 315580 201912
rect 315632 201900 315638 201952
rect 374362 201900 374368 201952
rect 374420 201940 374426 201952
rect 379974 201940 379980 201952
rect 374420 201912 379980 201940
rect 374420 201900 374426 201912
rect 379974 201900 379980 201912
rect 380032 201900 380038 201952
rect 412266 201900 412272 201952
rect 412324 201940 412330 201952
rect 457438 201940 457444 201952
rect 412324 201912 457444 201940
rect 412324 201900 412330 201912
rect 457438 201900 457444 201912
rect 457496 201900 457502 201952
rect 412818 201832 412824 201884
rect 412876 201872 412882 201884
rect 417050 201872 417056 201884
rect 412876 201844 417056 201872
rect 412876 201832 412882 201844
rect 417050 201832 417056 201844
rect 417108 201832 417114 201884
rect 300452 201776 305960 201804
rect 300452 201764 300458 201776
rect 307110 201764 307116 201816
rect 307168 201804 307174 201816
rect 313642 201804 313648 201816
rect 307168 201776 313648 201804
rect 307168 201764 307174 201776
rect 313642 201764 313648 201776
rect 313700 201764 313706 201816
rect 414658 201764 414664 201816
rect 414716 201804 414722 201816
rect 418798 201804 418804 201816
rect 414716 201776 418804 201804
rect 414716 201764 414722 201776
rect 418798 201764 418804 201776
rect 418856 201764 418862 201816
rect 266044 201708 266814 201736
rect 266044 201696 266050 201708
rect 268102 201696 268108 201748
rect 268160 201736 268166 201748
rect 270586 201736 270592 201748
rect 268160 201708 270592 201736
rect 268160 201696 268166 201708
rect 270586 201696 270592 201708
rect 270644 201696 270650 201748
rect 272242 201696 272248 201748
rect 272300 201736 272306 201748
rect 273162 201736 273168 201748
rect 272300 201708 273168 201736
rect 272300 201696 272306 201708
rect 273162 201696 273168 201708
rect 273220 201696 273226 201748
rect 273622 201696 273628 201748
rect 273680 201736 273686 201748
rect 274450 201736 274456 201748
rect 273680 201708 274456 201736
rect 273680 201696 273686 201708
rect 274450 201696 274456 201708
rect 274508 201696 274514 201748
rect 275278 201696 275284 201748
rect 275336 201736 275342 201748
rect 275830 201736 275836 201748
rect 275336 201708 275836 201736
rect 275336 201696 275342 201708
rect 275830 201696 275836 201708
rect 275888 201696 275894 201748
rect 279234 201696 279240 201748
rect 279292 201736 279298 201748
rect 280062 201736 280068 201748
rect 279292 201708 280068 201736
rect 279292 201696 279298 201708
rect 280062 201696 280068 201708
rect 280120 201696 280126 201748
rect 298370 201696 298376 201748
rect 298428 201736 298434 201748
rect 301038 201736 301044 201748
rect 298428 201708 301044 201736
rect 298428 201696 298434 201708
rect 301038 201696 301044 201708
rect 301096 201696 301102 201748
rect 311342 201736 311348 201748
rect 301148 201708 311348 201736
rect 198550 201628 198556 201680
rect 198608 201668 198614 201680
rect 212534 201668 212540 201680
rect 198608 201640 212540 201668
rect 198608 201628 198614 201640
rect 212534 201628 212540 201640
rect 212592 201628 212598 201680
rect 244642 201628 244648 201680
rect 244700 201668 244706 201680
rect 253842 201668 253848 201680
rect 244700 201640 253848 201668
rect 244700 201628 244706 201640
rect 253842 201628 253848 201640
rect 253900 201628 253906 201680
rect 258350 201628 258356 201680
rect 258408 201668 258414 201680
rect 266722 201668 266728 201680
rect 258408 201640 266728 201668
rect 258408 201628 258414 201640
rect 266722 201628 266728 201640
rect 266780 201628 266786 201680
rect 270770 201668 270776 201680
rect 266832 201640 270776 201668
rect 127618 201560 127624 201612
rect 127676 201600 127682 201612
rect 134150 201600 134156 201612
rect 127676 201572 134156 201600
rect 127676 201560 127682 201572
rect 134150 201560 134156 201572
rect 134208 201560 134214 201612
rect 198458 201560 198464 201612
rect 198516 201600 198522 201612
rect 211154 201600 211160 201612
rect 198516 201572 211160 201600
rect 198516 201560 198522 201572
rect 211154 201560 211160 201572
rect 211212 201560 211218 201612
rect 258718 201560 258724 201612
rect 258776 201600 258782 201612
rect 266354 201600 266360 201612
rect 258776 201572 266360 201600
rect 258776 201560 258782 201572
rect 266354 201560 266360 201572
rect 266412 201560 266418 201612
rect 266832 201600 266860 201640
rect 270770 201628 270776 201640
rect 270828 201628 270834 201680
rect 297358 201628 297364 201680
rect 297416 201668 297422 201680
rect 301148 201668 301176 201708
rect 311342 201696 311348 201708
rect 311400 201696 311406 201748
rect 297416 201640 301176 201668
rect 297416 201628 297422 201640
rect 301866 201628 301872 201680
rect 301924 201668 301930 201680
rect 312630 201668 312636 201680
rect 301924 201640 312636 201668
rect 301924 201628 301930 201640
rect 312630 201628 312636 201640
rect 312688 201628 312694 201680
rect 266556 201572 266860 201600
rect 198826 201492 198832 201544
rect 198884 201532 198890 201544
rect 211706 201532 211712 201544
rect 198884 201504 211712 201532
rect 198884 201492 198890 201504
rect 211706 201492 211712 201504
rect 211764 201492 211770 201544
rect 266446 201532 266452 201544
rect 258920 201504 266452 201532
rect 8018 201424 8024 201476
rect 8076 201464 8082 201476
rect 8110 201464 8116 201476
rect 8076 201436 8116 201464
rect 8076 201424 8082 201436
rect 8110 201424 8116 201436
rect 8168 201424 8174 201476
rect 252738 201424 252744 201476
rect 252796 201464 252802 201476
rect 258920 201464 258948 201504
rect 266446 201492 266452 201504
rect 266504 201492 266510 201544
rect 252796 201436 258948 201464
rect 252796 201424 252802 201436
rect 265894 201424 265900 201476
rect 265952 201464 265958 201476
rect 266556 201464 266584 201572
rect 267090 201560 267096 201612
rect 267148 201600 267154 201612
rect 270494 201600 270500 201612
rect 267148 201572 270500 201600
rect 267148 201560 267154 201572
rect 270494 201560 270500 201572
rect 270552 201560 270558 201612
rect 298738 201560 298744 201612
rect 298796 201600 298802 201612
rect 307294 201600 307300 201612
rect 298796 201572 307300 201600
rect 298796 201560 298802 201572
rect 307294 201560 307300 201572
rect 307352 201560 307358 201612
rect 266630 201492 266636 201544
rect 266688 201532 266694 201544
rect 268010 201532 268016 201544
rect 266688 201504 268016 201532
rect 266688 201492 266694 201504
rect 268010 201492 268016 201504
rect 268068 201492 268074 201544
rect 297634 201492 297640 201544
rect 297692 201532 297698 201544
rect 306926 201532 306932 201544
rect 297692 201504 306932 201532
rect 297692 201492 297698 201504
rect 306926 201492 306932 201504
rect 306984 201492 306990 201544
rect 355318 201492 355324 201544
rect 355376 201532 355382 201544
rect 355962 201532 355968 201544
rect 355376 201504 355968 201532
rect 355376 201492 355382 201504
rect 355962 201492 355968 201504
rect 356020 201492 356026 201544
rect 359642 201492 359648 201544
rect 359700 201532 359706 201544
rect 360102 201532 360108 201544
rect 359700 201504 360108 201532
rect 359700 201492 359706 201504
rect 360102 201492 360108 201504
rect 360160 201492 360166 201544
rect 360562 201492 360568 201544
rect 360620 201532 360626 201544
rect 361390 201532 361396 201544
rect 360620 201504 361396 201532
rect 360620 201492 360626 201504
rect 361390 201492 361396 201504
rect 361448 201492 361454 201544
rect 362310 201492 362316 201544
rect 362368 201532 362374 201544
rect 362770 201532 362776 201544
rect 362368 201504 362776 201532
rect 362368 201492 362374 201504
rect 362770 201492 362776 201504
rect 362828 201492 362834 201544
rect 400950 201492 400956 201544
rect 401008 201532 401014 201544
rect 401502 201532 401508 201544
rect 401008 201504 401508 201532
rect 401008 201492 401014 201504
rect 401502 201492 401508 201504
rect 401560 201492 401566 201544
rect 265952 201436 266584 201464
rect 265952 201424 265958 201436
rect 504174 201220 504180 201272
rect 504232 201260 504238 201272
rect 504450 201260 504456 201272
rect 504232 201232 504456 201260
rect 504232 201220 504238 201232
rect 504450 201220 504456 201232
rect 504508 201220 504514 201272
rect 4062 201152 4068 201204
rect 4120 201192 4126 201204
rect 436646 201192 436652 201204
rect 4120 201164 436652 201192
rect 4120 201152 4126 201164
rect 436646 201152 436652 201164
rect 436704 201152 436710 201204
rect 3878 201084 3884 201136
rect 3936 201124 3942 201136
rect 436554 201124 436560 201136
rect 3936 201096 436560 201124
rect 3936 201084 3942 201096
rect 436554 201084 436560 201096
rect 436612 201084 436618 201136
rect 2774 201016 2780 201068
rect 2832 201056 2838 201068
rect 436738 201056 436744 201068
rect 2832 201028 436744 201056
rect 2832 201016 2838 201028
rect 436738 201016 436744 201028
rect 436796 201016 436802 201068
rect 132402 200948 132408 201000
rect 132460 200988 132466 201000
rect 580718 200988 580724 201000
rect 132460 200960 580724 200988
rect 132460 200948 132466 200960
rect 580718 200948 580724 200960
rect 580776 200948 580782 201000
rect 131298 200880 131304 200932
rect 131356 200920 131362 200932
rect 580350 200920 580356 200932
rect 131356 200892 580356 200920
rect 131356 200880 131362 200892
rect 580350 200880 580356 200892
rect 580408 200880 580414 200932
rect 131390 200812 131396 200864
rect 131448 200852 131454 200864
rect 580626 200852 580632 200864
rect 131448 200824 580632 200852
rect 131448 200812 131454 200824
rect 580626 200812 580632 200824
rect 580684 200812 580690 200864
rect 131482 200744 131488 200796
rect 131540 200784 131546 200796
rect 580902 200784 580908 200796
rect 131540 200756 580908 200784
rect 131540 200744 131546 200756
rect 580902 200744 580908 200756
rect 580960 200744 580966 200796
rect 248690 200200 248696 200252
rect 248748 200240 248754 200252
rect 249380 200240 249386 200252
rect 248748 200212 249386 200240
rect 248748 200200 248754 200212
rect 249380 200200 249386 200212
rect 249438 200200 249444 200252
rect 254992 200200 254998 200252
rect 255050 200240 255056 200252
rect 258902 200240 258908 200252
rect 255050 200212 258908 200240
rect 255050 200200 255056 200212
rect 258902 200200 258908 200212
rect 258960 200200 258966 200252
rect 308536 200200 308542 200252
rect 308594 200240 308600 200252
rect 308766 200240 308772 200252
rect 308594 200212 308772 200240
rect 308594 200200 308600 200212
rect 308766 200200 308772 200212
rect 308824 200200 308830 200252
rect 133782 200132 133788 200184
rect 133840 200172 133846 200184
rect 579982 200172 579988 200184
rect 133840 200144 579988 200172
rect 133840 200132 133846 200144
rect 579982 200132 579988 200144
rect 580040 200132 580046 200184
rect 133506 200064 133512 200116
rect 133564 200104 133570 200116
rect 135254 200104 135260 200116
rect 133564 200076 135260 200104
rect 133564 200064 133570 200076
rect 135254 200064 135260 200076
rect 135312 200064 135318 200116
rect 238754 199860 238760 199912
rect 238812 199900 238818 199912
rect 239490 199900 239496 199912
rect 238812 199872 239496 199900
rect 238812 199860 238818 199872
rect 239490 199860 239496 199872
rect 239548 199860 239554 199912
rect 2774 199792 2780 199844
rect 2832 199832 2838 199844
rect 436278 199832 436284 199844
rect 2832 199804 436284 199832
rect 2832 199792 2838 199804
rect 436278 199792 436284 199804
rect 436336 199792 436342 199844
rect 3878 198704 3884 198756
rect 3936 198744 3942 198756
rect 131206 198744 131212 198756
rect 3936 198716 131212 198744
rect 3936 198704 3942 198716
rect 131206 198704 131212 198716
rect 131264 198704 131270 198756
rect 4062 197344 4068 197396
rect 4120 197384 4126 197396
rect 131206 197384 131212 197396
rect 4120 197356 131212 197384
rect 4120 197344 4126 197356
rect 131206 197344 131212 197356
rect 131264 197344 131270 197396
rect 131298 196324 131304 196376
rect 131356 196364 131362 196376
rect 131356 196336 131436 196364
rect 131356 196324 131362 196336
rect 14458 196052 14464 196104
rect 14516 196092 14522 196104
rect 131408 196092 131436 196336
rect 14516 196064 131436 196092
rect 14516 196052 14522 196064
rect 5350 195984 5356 196036
rect 5408 196024 5414 196036
rect 131206 196024 131212 196036
rect 5408 195996 131212 196024
rect 5408 195984 5414 195996
rect 131206 195984 131212 195996
rect 131264 195984 131270 196036
rect 122742 195848 122748 195900
rect 122800 195888 122806 195900
rect 122926 195888 122932 195900
rect 122800 195860 122932 195888
rect 122800 195848 122806 195860
rect 122926 195848 122932 195860
rect 122984 195848 122990 195900
rect 128354 195848 128360 195900
rect 128412 195888 128418 195900
rect 128538 195888 128544 195900
rect 128412 195860 128544 195888
rect 128412 195848 128418 195860
rect 128538 195848 128544 195860
rect 128596 195848 128602 195900
rect 128722 195576 128728 195628
rect 128780 195616 128786 195628
rect 129090 195616 129096 195628
rect 128780 195588 129096 195616
rect 128780 195576 128786 195588
rect 129090 195576 129096 195588
rect 129148 195576 129154 195628
rect 8938 194556 8944 194608
rect 8996 194596 9002 194608
rect 131206 194596 131212 194608
rect 8996 194568 131212 194596
rect 8996 194556 9002 194568
rect 131206 194556 131212 194568
rect 131264 194556 131270 194608
rect 6178 194420 6184 194472
rect 6236 194460 6242 194472
rect 131206 194460 131212 194472
rect 6236 194432 131212 194460
rect 6236 194420 6242 194432
rect 131206 194420 131212 194432
rect 131264 194420 131270 194472
rect 5166 193128 5172 193180
rect 5224 193168 5230 193180
rect 5224 193140 131344 193168
rect 5224 193128 5230 193140
rect 5258 193060 5264 193112
rect 5316 193100 5322 193112
rect 131206 193100 131212 193112
rect 5316 193072 131212 193100
rect 5316 193060 5322 193072
rect 131206 193060 131212 193072
rect 131264 193060 131270 193112
rect 131206 192788 131212 192840
rect 131264 192828 131270 192840
rect 131316 192828 131344 193140
rect 436278 192924 436284 192976
rect 436336 192964 436342 192976
rect 436830 192964 436836 192976
rect 436336 192936 436836 192964
rect 436336 192924 436342 192936
rect 436830 192924 436836 192936
rect 436888 192924 436894 192976
rect 131264 192800 131344 192828
rect 131264 192788 131270 192800
rect 4982 191768 4988 191820
rect 5040 191808 5046 191820
rect 131206 191808 131212 191820
rect 5040 191780 131212 191808
rect 5040 191768 5046 191780
rect 131206 191768 131212 191780
rect 131264 191768 131270 191820
rect 128722 191088 128728 191140
rect 128780 191128 128786 191140
rect 129090 191128 129096 191140
rect 128780 191100 129096 191128
rect 128780 191088 128786 191100
rect 129090 191088 129096 191100
rect 129148 191088 129154 191140
rect 3234 190408 3240 190460
rect 3292 190448 3298 190460
rect 131206 190448 131212 190460
rect 3292 190420 131212 190448
rect 3292 190408 3298 190420
rect 131206 190408 131212 190420
rect 131264 190408 131270 190460
rect 133506 189904 133512 189916
rect 133432 189876 133512 189904
rect 133432 189632 133460 189876
rect 133506 189864 133512 189876
rect 133564 189864 133570 189916
rect 133506 189728 133512 189780
rect 133564 189768 133570 189780
rect 133782 189768 133788 189780
rect 133564 189740 133788 189768
rect 133564 189728 133570 189740
rect 133782 189728 133788 189740
rect 133840 189728 133846 189780
rect 133782 189632 133788 189644
rect 133432 189604 133788 189632
rect 133782 189592 133788 189604
rect 133840 189592 133846 189644
rect 4890 188980 4896 189032
rect 4948 189020 4954 189032
rect 131206 189020 131212 189032
rect 4948 188992 131212 189020
rect 4948 188980 4954 188992
rect 131206 188980 131212 188992
rect 131264 188980 131270 189032
rect 4798 188844 4804 188896
rect 4856 188884 4862 188896
rect 4856 188856 9628 188884
rect 4856 188844 4862 188856
rect 9600 188816 9628 188856
rect 9674 188844 9680 188896
rect 9732 188844 9738 188896
rect 19242 188844 19248 188896
rect 19300 188884 19306 188896
rect 22094 188884 22100 188896
rect 19300 188856 22100 188884
rect 19300 188844 19306 188856
rect 22094 188844 22100 188856
rect 22152 188844 22158 188896
rect 22186 188844 22192 188896
rect 22244 188884 22250 188896
rect 22244 188856 28948 188884
rect 22244 188844 22250 188856
rect 9692 188816 9720 188844
rect 9600 188788 9720 188816
rect 28920 188816 28948 188856
rect 67634 188816 67640 188828
rect 28920 188788 31708 188816
rect 31680 188680 31708 188788
rect 60844 188788 67640 188816
rect 41506 188708 41512 188760
rect 41564 188748 41570 188760
rect 41564 188720 48360 188748
rect 41564 188708 41570 188720
rect 48332 188692 48360 188720
rect 60734 188708 60740 188760
rect 60792 188748 60798 188760
rect 60844 188748 60872 188788
rect 67634 188776 67640 188788
rect 67692 188776 67698 188828
rect 86954 188816 86960 188828
rect 81268 188788 86960 188816
rect 60792 188720 60872 188748
rect 60792 188708 60798 188720
rect 77202 188708 77208 188760
rect 77260 188748 77266 188760
rect 79962 188748 79968 188760
rect 77260 188720 79968 188748
rect 77260 188708 77266 188720
rect 79962 188708 79968 188720
rect 80020 188708 80026 188760
rect 80054 188708 80060 188760
rect 80112 188748 80118 188760
rect 81268 188748 81296 188788
rect 86954 188776 86960 188788
rect 87012 188776 87018 188828
rect 115934 188816 115940 188828
rect 108960 188788 115940 188816
rect 108960 188748 108988 188788
rect 115934 188776 115940 188788
rect 115992 188776 115998 188828
rect 80112 188720 81296 188748
rect 106200 188720 108988 188748
rect 80112 188708 80118 188720
rect 41322 188680 41328 188692
rect 31680 188652 41328 188680
rect 41322 188640 41328 188652
rect 41380 188640 41386 188692
rect 48314 188640 48320 188692
rect 48372 188640 48378 188692
rect 57882 188640 57888 188692
rect 57940 188680 57946 188692
rect 60642 188680 60648 188692
rect 57940 188652 60648 188680
rect 57940 188640 57946 188652
rect 60642 188640 60648 188652
rect 60700 188640 60706 188692
rect 96522 188640 96528 188692
rect 96580 188680 96586 188692
rect 99374 188680 99380 188692
rect 96580 188652 99380 188680
rect 96580 188640 96586 188652
rect 99374 188640 99380 188652
rect 99432 188640 99438 188692
rect 99466 188640 99472 188692
rect 99524 188680 99530 188692
rect 106200 188680 106228 188720
rect 125502 188708 125508 188760
rect 125560 188708 125566 188760
rect 99524 188652 106228 188680
rect 125520 188680 125548 188708
rect 125520 188652 131252 188680
rect 99524 188640 99530 188652
rect 131224 188624 131252 188652
rect 131206 188572 131212 188624
rect 131264 188572 131270 188624
rect 48314 188504 48320 188556
rect 48372 188544 48378 188556
rect 57882 188544 57888 188556
rect 48372 188516 57888 188544
rect 48372 188504 48378 188516
rect 57882 188504 57888 188516
rect 57940 188504 57946 188556
rect 3694 187620 3700 187672
rect 3752 187660 3758 187672
rect 131206 187660 131212 187672
rect 3752 187632 131212 187660
rect 3752 187620 3758 187632
rect 131206 187620 131212 187632
rect 131264 187620 131270 187672
rect 3510 186260 3516 186312
rect 3568 186300 3574 186312
rect 131206 186300 131212 186312
rect 3568 186272 131212 186300
rect 3568 186260 3574 186272
rect 131206 186260 131212 186272
rect 131264 186260 131270 186312
rect 132862 185172 132868 185224
rect 132920 185212 132926 185224
rect 133138 185212 133144 185224
rect 132920 185184 133144 185212
rect 132920 185172 132926 185184
rect 133138 185172 133144 185184
rect 133196 185172 133202 185224
rect 132862 184968 132868 185020
rect 132920 185008 132926 185020
rect 133046 185008 133052 185020
rect 132920 184980 133052 185008
rect 132920 184968 132926 184980
rect 133046 184968 133052 184980
rect 133104 184968 133110 185020
rect 8294 184832 8300 184884
rect 8352 184872 8358 184884
rect 131206 184872 131212 184884
rect 8352 184844 131212 184872
rect 8352 184832 8358 184844
rect 131206 184832 131212 184844
rect 131264 184832 131270 184884
rect 128354 183540 128360 183592
rect 128412 183580 128418 183592
rect 128538 183580 128544 183592
rect 128412 183552 128544 183580
rect 128412 183540 128418 183552
rect 128538 183540 128544 183552
rect 128596 183540 128602 183592
rect 72418 183472 72424 183524
rect 72476 183512 72482 183524
rect 131206 183512 131212 183524
rect 72476 183484 131212 183512
rect 72476 183472 72482 183484
rect 131206 183472 131212 183484
rect 131264 183472 131270 183524
rect 132586 181228 132592 181280
rect 132644 181268 132650 181280
rect 133230 181268 133236 181280
rect 132644 181240 133236 181268
rect 132644 181228 132650 181240
rect 133230 181228 133236 181240
rect 133288 181228 133294 181280
rect 3694 179460 3700 179512
rect 3752 179500 3758 179512
rect 8938 179500 8944 179512
rect 3752 179472 8944 179500
rect 3752 179460 3758 179472
rect 8938 179460 8944 179472
rect 8996 179460 9002 179512
rect 128722 177352 128728 177404
rect 128780 177392 128786 177404
rect 129090 177392 129096 177404
rect 128780 177364 129096 177392
rect 128780 177352 128786 177364
rect 129090 177352 129096 177364
rect 129148 177352 129154 177404
rect 122742 176712 122748 176724
rect 122668 176684 122748 176712
rect 122668 176588 122696 176684
rect 122742 176672 122748 176684
rect 122800 176672 122806 176724
rect 128538 176672 128544 176724
rect 128596 176672 128602 176724
rect 122650 176536 122656 176588
rect 122708 176536 122714 176588
rect 128556 176576 128584 176672
rect 128630 176576 128636 176588
rect 128556 176548 128636 176576
rect 128630 176536 128636 176548
rect 128688 176536 128694 176588
rect 128722 175584 128728 175636
rect 128780 175624 128786 175636
rect 129090 175624 129096 175636
rect 128780 175596 129096 175624
rect 128780 175584 128786 175596
rect 129090 175584 129096 175596
rect 129148 175584 129154 175636
rect 129642 175176 129648 175228
rect 129700 175216 129706 175228
rect 131206 175216 131212 175228
rect 129700 175188 131212 175216
rect 129700 175176 129706 175188
rect 131206 175176 131212 175188
rect 131264 175176 131270 175228
rect 129550 175108 129556 175160
rect 129608 175148 129614 175160
rect 132034 175148 132040 175160
rect 129608 175120 132040 175148
rect 129608 175108 129614 175120
rect 132034 175108 132040 175120
rect 132092 175108 132098 175160
rect 504450 173884 504456 173936
rect 504508 173924 504514 173936
rect 504634 173924 504640 173936
rect 504508 173896 504640 173924
rect 504508 173884 504514 173896
rect 504634 173884 504640 173896
rect 504692 173884 504698 173936
rect 128354 169056 128360 169108
rect 128412 169096 128418 169108
rect 128538 169096 128544 169108
rect 128412 169068 128544 169096
rect 128412 169056 128418 169068
rect 128538 169056 128544 169068
rect 128596 169056 128602 169108
rect 133046 168648 133052 168700
rect 133104 168648 133110 168700
rect 133064 168496 133092 168648
rect 133046 168444 133052 168496
rect 133104 168444 133110 168496
rect 130010 166812 130016 166864
rect 130068 166852 130074 166864
rect 132034 166852 132040 166864
rect 130068 166824 132040 166852
rect 130068 166812 130074 166824
rect 132034 166812 132040 166824
rect 132092 166812 132098 166864
rect 504174 164160 504180 164212
rect 504232 164200 504238 164212
rect 504358 164200 504364 164212
rect 504232 164172 504364 164200
rect 504232 164160 504238 164172
rect 504358 164160 504364 164172
rect 504416 164160 504422 164212
rect 128722 162120 128728 162172
rect 128780 162160 128786 162172
rect 129090 162160 129096 162172
rect 128780 162132 129096 162160
rect 128780 162120 128786 162132
rect 129090 162120 129096 162132
rect 129148 162120 129154 162172
rect 122558 161440 122564 161492
rect 122616 161480 122622 161492
rect 122742 161480 122748 161492
rect 122616 161452 122748 161480
rect 122616 161440 122622 161452
rect 122742 161440 122748 161452
rect 122800 161440 122806 161492
rect 4798 158720 4804 158772
rect 4856 158760 4862 158772
rect 131206 158760 131212 158772
rect 4856 158732 131212 158760
rect 4856 158720 4862 158732
rect 131206 158720 131212 158732
rect 131264 158720 131270 158772
rect 4154 155932 4160 155984
rect 4212 155972 4218 155984
rect 131206 155972 131212 155984
rect 4212 155944 131212 155972
rect 4212 155932 4218 155944
rect 131206 155932 131212 155944
rect 131264 155932 131270 155984
rect 3050 155864 3056 155916
rect 3108 155904 3114 155916
rect 3108 155876 131252 155904
rect 3108 155864 3114 155876
rect 131224 155848 131252 155876
rect 131206 155796 131212 155848
rect 131264 155796 131270 155848
rect 436094 155592 436100 155644
rect 436152 155632 436158 155644
rect 438118 155632 438124 155644
rect 436152 155604 438124 155632
rect 436152 155592 436158 155604
rect 438118 155592 438124 155604
rect 438176 155592 438182 155644
rect 2866 154504 2872 154556
rect 2924 154544 2930 154556
rect 131206 154544 131212 154556
rect 2924 154516 131212 154544
rect 2924 154504 2930 154516
rect 131206 154504 131212 154516
rect 131264 154504 131270 154556
rect 2958 153144 2964 153196
rect 3016 153184 3022 153196
rect 131206 153184 131212 153196
rect 3016 153156 131212 153184
rect 3016 153144 3022 153156
rect 131206 153144 131212 153156
rect 131264 153144 131270 153196
rect 5074 153076 5080 153128
rect 5132 153116 5138 153128
rect 5132 153088 6868 153116
rect 5132 153076 5138 153088
rect 6840 153048 6868 153088
rect 6914 153076 6920 153128
rect 6972 153076 6978 153128
rect 31680 153088 70348 153116
rect 6932 153048 6960 153076
rect 31680 153048 31708 153088
rect 6840 153020 6960 153048
rect 22204 153020 31708 153048
rect 70320 153048 70348 153088
rect 82814 153076 82820 153128
rect 82872 153076 82878 153128
rect 82906 153076 82912 153128
rect 82964 153116 82970 153128
rect 82964 153088 93900 153116
rect 82964 153076 82970 153088
rect 82832 153048 82860 153076
rect 70320 153020 71912 153048
rect 16482 152940 16488 152992
rect 16540 152980 16546 152992
rect 16540 152952 21036 152980
rect 16540 152940 16546 152952
rect 21008 152912 21036 152952
rect 22204 152912 22232 153020
rect 71884 152980 71912 153020
rect 80164 153020 82860 153048
rect 93872 153048 93900 153088
rect 93872 153020 108988 153048
rect 80164 152980 80192 153020
rect 71884 152952 80192 152980
rect 108960 152980 108988 153020
rect 116302 152980 116308 152992
rect 108960 152952 116308 152980
rect 116302 152940 116308 152952
rect 116360 152940 116366 152992
rect 21008 152884 22232 152912
rect 116302 152804 116308 152856
rect 116360 152844 116366 152856
rect 131206 152844 131212 152856
rect 116360 152816 131212 152844
rect 116360 152804 116366 152816
rect 131206 152804 131212 152816
rect 131264 152804 131270 152856
rect 437382 151920 437388 151972
rect 437440 151960 437446 151972
rect 442258 151960 442264 151972
rect 437440 151932 442264 151960
rect 437440 151920 437446 151932
rect 442258 151920 442264 151932
rect 442316 151920 442322 151972
rect 3142 151716 3148 151768
rect 3200 151756 3206 151768
rect 131206 151756 131212 151768
rect 3200 151728 131212 151756
rect 3200 151716 3206 151728
rect 131206 151716 131212 151728
rect 131264 151716 131270 151768
rect 3326 150356 3332 150408
rect 3384 150396 3390 150408
rect 131206 150396 131212 150408
rect 3384 150368 131212 150396
rect 3384 150356 3390 150368
rect 131206 150356 131212 150368
rect 131264 150356 131270 150408
rect 437014 150288 437020 150340
rect 437072 150328 437078 150340
rect 440878 150328 440884 150340
rect 437072 150300 440884 150328
rect 437072 150288 437078 150300
rect 440878 150288 440884 150300
rect 440936 150288 440942 150340
rect 128722 149812 128728 149864
rect 128780 149852 128786 149864
rect 129090 149852 129096 149864
rect 128780 149824 129096 149852
rect 128780 149812 128786 149824
rect 129090 149812 129096 149824
rect 129148 149812 129154 149864
rect 3970 148996 3976 149048
rect 4028 149036 4034 149048
rect 131206 149036 131212 149048
rect 4028 149008 131212 149036
rect 4028 148996 4034 149008
rect 131206 148996 131212 149008
rect 131264 148996 131270 149048
rect 115934 148860 115940 148912
rect 115992 148860 115998 148912
rect 436186 148860 436192 148912
rect 436244 148900 436250 148912
rect 439498 148900 439504 148912
rect 436244 148872 439504 148900
rect 436244 148860 436250 148872
rect 439498 148860 439504 148872
rect 439556 148860 439562 148912
rect 70394 148792 70400 148844
rect 70452 148832 70458 148844
rect 84194 148832 84200 148844
rect 70452 148804 74488 148832
rect 70452 148792 70458 148804
rect 22186 148724 22192 148776
rect 22244 148764 22250 148776
rect 22244 148736 26280 148764
rect 22244 148724 22250 148736
rect 26252 148708 26280 148736
rect 41506 148724 41512 148776
rect 41564 148764 41570 148776
rect 50982 148764 50988 148776
rect 41564 148736 50988 148764
rect 41564 148724 41570 148736
rect 50982 148724 50988 148736
rect 51040 148724 51046 148776
rect 56594 148724 56600 148776
rect 56652 148764 56658 148776
rect 64874 148764 64880 148776
rect 56652 148736 64880 148764
rect 56652 148724 56658 148736
rect 64874 148724 64880 148736
rect 64932 148724 64938 148776
rect 74460 148764 74488 148804
rect 80164 148804 84200 148832
rect 79962 148764 79968 148776
rect 74460 148736 79968 148764
rect 79962 148724 79968 148736
rect 80020 148724 80026 148776
rect 80054 148724 80060 148776
rect 80112 148764 80118 148776
rect 80164 148764 80192 148804
rect 84194 148792 84200 148804
rect 84252 148792 84258 148844
rect 115952 148832 115980 148860
rect 108960 148804 115980 148832
rect 108960 148764 108988 148804
rect 80112 148736 80192 148764
rect 103440 148736 108988 148764
rect 80112 148724 80118 148736
rect 3786 148656 3792 148708
rect 3844 148696 3850 148708
rect 22002 148696 22008 148708
rect 3844 148668 22008 148696
rect 3844 148656 3850 148668
rect 22002 148656 22008 148668
rect 22060 148656 22066 148708
rect 26234 148656 26240 148708
rect 26292 148656 26298 148708
rect 35802 148656 35808 148708
rect 35860 148696 35866 148708
rect 41322 148696 41328 148708
rect 35860 148668 41328 148696
rect 35860 148656 35866 148668
rect 41322 148656 41328 148668
rect 41380 148656 41386 148708
rect 51074 148656 51080 148708
rect 51132 148696 51138 148708
rect 56502 148696 56508 148708
rect 51132 148668 56508 148696
rect 51132 148656 51138 148668
rect 56502 148656 56508 148668
rect 56560 148656 56566 148708
rect 93762 148656 93768 148708
rect 93820 148696 93826 148708
rect 99374 148696 99380 148708
rect 93820 148668 99380 148696
rect 93820 148656 93826 148668
rect 99374 148656 99380 148668
rect 99432 148656 99438 148708
rect 99466 148656 99472 148708
rect 99524 148696 99530 148708
rect 103440 148696 103468 148736
rect 99524 148668 103468 148696
rect 99524 148656 99530 148668
rect 116026 148588 116032 148640
rect 116084 148628 116090 148640
rect 131206 148628 131212 148640
rect 116084 148600 131212 148628
rect 116084 148588 116090 148600
rect 131206 148588 131212 148600
rect 131264 148588 131270 148640
rect 26234 148520 26240 148572
rect 26292 148560 26298 148572
rect 35802 148560 35808 148572
rect 26292 148532 35808 148560
rect 26292 148520 26298 148532
rect 35802 148520 35808 148532
rect 35860 148520 35866 148572
rect 130930 148180 130936 148232
rect 130988 148220 130994 148232
rect 131206 148220 131212 148232
rect 130988 148192 131212 148220
rect 130988 148180 130994 148192
rect 131206 148180 131212 148192
rect 131264 148180 131270 148232
rect 3602 147568 3608 147620
rect 3660 147608 3666 147620
rect 132218 147608 132224 147620
rect 3660 147580 132224 147608
rect 3660 147568 3666 147580
rect 132218 147568 132224 147580
rect 132276 147568 132282 147620
rect 132310 147568 132316 147620
rect 132368 147568 132374 147620
rect 122558 147500 122564 147552
rect 122616 147540 122622 147552
rect 122742 147540 122748 147552
rect 122616 147512 122748 147540
rect 122616 147500 122622 147512
rect 122742 147500 122748 147512
rect 122800 147500 122806 147552
rect 132328 147540 132356 147568
rect 132236 147512 132356 147540
rect 132236 146600 132264 147512
rect 132218 146548 132224 146600
rect 132276 146548 132282 146600
rect 130930 146344 130936 146396
rect 130988 146384 130994 146396
rect 131114 146384 131120 146396
rect 130988 146356 131120 146384
rect 130988 146344 130994 146356
rect 131114 146344 131120 146356
rect 131172 146344 131178 146396
rect 3418 146208 3424 146260
rect 3476 146248 3482 146260
rect 131114 146248 131120 146260
rect 3476 146220 131120 146248
rect 3476 146208 3482 146220
rect 131114 146208 131120 146220
rect 131172 146208 131178 146260
rect 436094 146208 436100 146260
rect 436152 146248 436158 146260
rect 438210 146248 438216 146260
rect 436152 146220 438216 146248
rect 436152 146208 436158 146220
rect 438210 146208 438216 146220
rect 438268 146208 438274 146260
rect 24762 144848 24768 144900
rect 24820 144888 24826 144900
rect 131114 144888 131120 144900
rect 24820 144860 115980 144888
rect 24820 144848 24826 144860
rect 115952 144820 115980 144860
rect 122668 144860 131120 144888
rect 122668 144820 122696 144860
rect 131114 144848 131120 144860
rect 131172 144848 131178 144900
rect 437382 144848 437388 144900
rect 437440 144888 437446 144900
rect 580258 144888 580264 144900
rect 437440 144860 580264 144888
rect 437440 144848 437446 144860
rect 580258 144848 580264 144860
rect 580316 144848 580322 144900
rect 115952 144792 122696 144820
rect 131022 144440 131028 144492
rect 131080 144440 131086 144492
rect 131040 144152 131068 144440
rect 131022 144100 131028 144152
rect 131080 144100 131086 144152
rect 128814 143488 128820 143540
rect 128872 143528 128878 143540
rect 129090 143528 129096 143540
rect 128872 143500 129096 143528
rect 128872 143488 128878 143500
rect 129090 143488 129096 143500
rect 129148 143488 129154 143540
rect 436094 142060 436100 142112
rect 436152 142100 436158 142112
rect 438302 142100 438308 142112
rect 436152 142072 438308 142100
rect 436152 142060 436158 142072
rect 438302 142060 438308 142072
rect 438360 142060 438366 142112
rect 437382 140700 437388 140752
rect 437440 140740 437446 140752
rect 580442 140740 580448 140752
rect 437440 140712 580448 140740
rect 437440 140700 437446 140712
rect 580442 140700 580448 140712
rect 580500 140700 580506 140752
rect 122558 137980 122564 138032
rect 122616 137980 122622 138032
rect 122576 137884 122604 137980
rect 437382 137912 437388 137964
rect 437440 137952 437446 137964
rect 580534 137952 580540 137964
rect 437440 137924 580540 137952
rect 437440 137912 437446 137924
rect 580534 137912 580540 137924
rect 580592 137912 580598 137964
rect 122650 137884 122656 137896
rect 122576 137856 122656 137884
rect 122650 137844 122656 137856
rect 122708 137844 122714 137896
rect 437014 136552 437020 136604
rect 437072 136592 437078 136604
rect 504450 136592 504456 136604
rect 437072 136564 504456 136592
rect 437072 136552 437078 136564
rect 504450 136552 504456 136564
rect 504508 136552 504514 136604
rect 2774 136348 2780 136400
rect 2832 136388 2838 136400
rect 5350 136388 5356 136400
rect 2832 136360 5356 136388
rect 2832 136348 2838 136360
rect 5350 136348 5356 136360
rect 5408 136348 5414 136400
rect 128630 135192 128636 135244
rect 128688 135232 128694 135244
rect 128722 135232 128728 135244
rect 128688 135204 128728 135232
rect 128688 135192 128694 135204
rect 128722 135192 128728 135204
rect 128780 135192 128786 135244
rect 128814 135192 128820 135244
rect 128872 135232 128878 135244
rect 129090 135232 129096 135244
rect 128872 135204 129096 135232
rect 128872 135192 128878 135204
rect 129090 135192 129096 135204
rect 129148 135192 129154 135244
rect 132862 135192 132868 135244
rect 132920 135192 132926 135244
rect 132880 135164 132908 135192
rect 132954 135164 132960 135176
rect 132880 135136 132960 135164
rect 132954 135124 132960 135136
rect 133012 135124 133018 135176
rect 437382 133832 437388 133884
rect 437440 133872 437446 133884
rect 580810 133872 580816 133884
rect 437440 133844 580816 133872
rect 437440 133832 437446 133844
rect 580810 133832 580816 133844
rect 580868 133832 580874 133884
rect 436830 132404 436836 132456
rect 436888 132444 436894 132456
rect 580166 132444 580172 132456
rect 436888 132416 580172 132444
rect 436888 132404 436894 132416
rect 580166 132404 580172 132416
rect 580224 132404 580230 132456
rect 128814 130364 128820 130416
rect 128872 130404 128878 130416
rect 129090 130404 129096 130416
rect 128872 130376 129096 130404
rect 128872 130364 128878 130376
rect 129090 130364 129096 130376
rect 129148 130364 129154 130416
rect 437382 129684 437388 129736
rect 437440 129724 437446 129736
rect 580074 129724 580080 129736
rect 437440 129696 580080 129724
rect 437440 129684 437446 129696
rect 580074 129684 580080 129696
rect 580132 129684 580138 129736
rect 128722 128324 128728 128376
rect 128780 128324 128786 128376
rect 128630 128256 128636 128308
rect 128688 128296 128694 128308
rect 128740 128296 128768 128324
rect 128688 128268 128768 128296
rect 128688 128256 128694 128268
rect 436094 128256 436100 128308
rect 436152 128296 436158 128308
rect 580626 128296 580632 128308
rect 436152 128268 580632 128296
rect 436152 128256 436158 128268
rect 580626 128256 580632 128268
rect 580684 128256 580690 128308
rect 128722 125536 128728 125588
rect 128780 125536 128786 125588
rect 128814 125536 128820 125588
rect 128872 125576 128878 125588
rect 129090 125576 129096 125588
rect 128872 125548 129096 125576
rect 128872 125536 128878 125548
rect 129090 125536 129096 125548
rect 129148 125536 129154 125588
rect 129182 125536 129188 125588
rect 129240 125536 129246 125588
rect 128740 125440 128768 125536
rect 129200 125452 129228 125536
rect 129090 125440 129096 125452
rect 128740 125412 129096 125440
rect 129090 125400 129096 125412
rect 129148 125400 129154 125452
rect 129182 125400 129188 125452
rect 129240 125400 129246 125452
rect 134058 120776 134064 120828
rect 134116 120816 134122 120828
rect 580902 120816 580908 120828
rect 134116 120788 580908 120816
rect 134116 120776 134122 120788
rect 580902 120776 580908 120788
rect 580960 120776 580966 120828
rect 133966 120708 133972 120760
rect 134024 120748 134030 120760
rect 580350 120748 580356 120760
rect 134024 120720 580356 120748
rect 134024 120708 134030 120720
rect 580350 120708 580356 120720
rect 580408 120708 580414 120760
rect 132402 120640 132408 120692
rect 132460 120680 132466 120692
rect 580258 120680 580264 120692
rect 132460 120652 580264 120680
rect 132460 120640 132466 120652
rect 580258 120640 580264 120652
rect 580316 120640 580322 120692
rect 3234 120572 3240 120624
rect 3292 120612 3298 120624
rect 436462 120612 436468 120624
rect 3292 120584 436468 120612
rect 3292 120572 3298 120584
rect 436462 120572 436468 120584
rect 436520 120572 436526 120624
rect 187786 119756 187792 119808
rect 187844 119796 187850 119808
rect 188752 119796 188758 119808
rect 187844 119768 188758 119796
rect 187844 119756 187850 119768
rect 188752 119756 188758 119768
rect 188810 119756 188816 119808
rect 205174 119756 205180 119808
rect 205232 119796 205238 119808
rect 210188 119796 210194 119808
rect 205232 119768 210194 119796
rect 205232 119756 205238 119768
rect 210188 119756 210194 119768
rect 210246 119756 210252 119808
rect 130194 119348 130200 119400
rect 130252 119388 130258 119400
rect 139394 119388 139400 119400
rect 130252 119360 139400 119388
rect 130252 119348 130258 119360
rect 139394 119348 139400 119360
rect 139452 119348 139458 119400
rect 143626 119348 143632 119400
rect 143684 119388 143690 119400
rect 144362 119388 144368 119400
rect 143684 119360 144368 119388
rect 143684 119348 143690 119360
rect 144362 119348 144368 119360
rect 144420 119348 144426 119400
rect 130838 119076 130844 119128
rect 130896 119116 130902 119128
rect 142246 119116 142252 119128
rect 130896 119088 142252 119116
rect 130896 119076 130902 119088
rect 142246 119076 142252 119088
rect 142304 119116 142310 119128
rect 142522 119116 142528 119128
rect 142304 119088 142528 119116
rect 142304 119076 142310 119088
rect 142522 119076 142528 119088
rect 142580 119076 142586 119128
rect 137186 118940 137192 118992
rect 137244 118980 137250 118992
rect 138290 118980 138296 118992
rect 137244 118952 138296 118980
rect 137244 118940 137250 118952
rect 138290 118940 138296 118952
rect 138348 118940 138354 118992
rect 129458 118872 129464 118924
rect 129516 118912 129522 118924
rect 145006 118912 145012 118924
rect 129516 118884 145012 118912
rect 129516 118872 129522 118884
rect 145006 118872 145012 118884
rect 145064 118872 145070 118924
rect 131022 118804 131028 118856
rect 131080 118844 131086 118856
rect 147766 118844 147772 118856
rect 131080 118816 147772 118844
rect 131080 118804 131086 118816
rect 147766 118804 147772 118816
rect 147824 118804 147830 118856
rect 129366 118736 129372 118788
rect 129424 118776 129430 118788
rect 149054 118776 149060 118788
rect 129424 118748 149060 118776
rect 129424 118736 129430 118748
rect 149054 118736 149060 118748
rect 149112 118736 149118 118788
rect 128262 118668 128268 118720
rect 128320 118708 128326 118720
rect 154666 118708 154672 118720
rect 128320 118680 154672 118708
rect 128320 118668 128326 118680
rect 154666 118668 154672 118680
rect 154724 118708 154730 118720
rect 155310 118708 155316 118720
rect 154724 118680 155316 118708
rect 154724 118668 154730 118680
rect 155310 118668 155316 118680
rect 155368 118668 155374 118720
rect 69842 118600 69848 118652
rect 69900 118640 69906 118652
rect 70302 118640 70308 118652
rect 69900 118612 70308 118640
rect 69900 118600 69906 118612
rect 70302 118600 70308 118612
rect 70360 118640 70366 118652
rect 138198 118640 138204 118652
rect 70360 118612 138204 118640
rect 70360 118600 70366 118612
rect 138198 118600 138204 118612
rect 138256 118600 138262 118652
rect 138290 118600 138296 118652
rect 138348 118640 138354 118652
rect 143074 118640 143080 118652
rect 138348 118612 143080 118640
rect 138348 118600 138354 118612
rect 143074 118600 143080 118612
rect 143132 118600 143138 118652
rect 146754 118600 146760 118652
rect 146812 118640 146818 118652
rect 157334 118640 157340 118652
rect 146812 118612 157340 118640
rect 146812 118600 146818 118612
rect 157334 118600 157340 118612
rect 157392 118600 157398 118652
rect 170398 118600 170404 118652
rect 170456 118640 170462 118652
rect 198182 118640 198188 118652
rect 170456 118612 198188 118640
rect 170456 118600 170462 118612
rect 198182 118600 198188 118612
rect 198240 118600 198246 118652
rect 200022 118600 200028 118652
rect 200080 118640 200086 118652
rect 236178 118640 236184 118652
rect 200080 118612 236184 118640
rect 200080 118600 200086 118612
rect 236178 118600 236184 118612
rect 236236 118600 236242 118652
rect 239398 118600 239404 118652
rect 239456 118640 239462 118652
rect 249794 118640 249800 118652
rect 239456 118612 249800 118640
rect 239456 118600 239462 118612
rect 249794 118600 249800 118612
rect 249852 118600 249858 118652
rect 249886 118600 249892 118652
rect 249944 118640 249950 118652
rect 258258 118640 258264 118652
rect 249944 118612 258264 118640
rect 249944 118600 249950 118612
rect 258258 118600 258264 118612
rect 258316 118600 258322 118652
rect 298646 118600 298652 118652
rect 298704 118640 298710 118652
rect 318978 118640 318984 118652
rect 298704 118612 318984 118640
rect 298704 118600 298710 118612
rect 318978 118600 318984 118612
rect 319036 118600 319042 118652
rect 349430 118600 349436 118652
rect 349488 118640 349494 118652
rect 416958 118640 416964 118652
rect 349488 118612 416964 118640
rect 349488 118600 349494 118612
rect 416958 118600 416964 118612
rect 417016 118600 417022 118652
rect 424778 118600 424784 118652
rect 424836 118640 424842 118652
rect 493318 118640 493324 118652
rect 424836 118612 493324 118640
rect 424836 118600 424842 118612
rect 493318 118600 493324 118612
rect 493376 118600 493382 118652
rect 97902 118532 97908 118584
rect 97960 118572 97966 118584
rect 181070 118572 181076 118584
rect 97960 118544 181076 118572
rect 97960 118532 97966 118544
rect 181070 118532 181076 118544
rect 181128 118532 181134 118584
rect 195882 118532 195888 118584
rect 195940 118572 195946 118584
rect 234706 118572 234712 118584
rect 195940 118544 234712 118572
rect 195940 118532 195946 118544
rect 234706 118532 234712 118544
rect 234764 118532 234770 118584
rect 240042 118532 240048 118584
rect 240100 118572 240106 118584
rect 256970 118572 256976 118584
rect 240100 118544 256976 118572
rect 240100 118532 240106 118544
rect 256970 118532 256976 118544
rect 257028 118532 257034 118584
rect 301130 118532 301136 118584
rect 301188 118572 301194 118584
rect 323118 118572 323124 118584
rect 301188 118544 323124 118572
rect 301188 118532 301194 118544
rect 323118 118532 323124 118544
rect 323176 118532 323182 118584
rect 364058 118532 364064 118584
rect 364116 118572 364122 118584
rect 380158 118572 380164 118584
rect 364116 118544 380164 118572
rect 364116 118532 364122 118544
rect 380158 118532 380164 118544
rect 380216 118532 380222 118584
rect 408218 118532 408224 118584
rect 408276 118572 408282 118584
rect 478138 118572 478144 118584
rect 408276 118544 478144 118572
rect 408276 118532 408282 118544
rect 478138 118532 478144 118544
rect 478196 118532 478202 118584
rect 82722 118464 82728 118516
rect 82780 118504 82786 118516
rect 164510 118504 164516 118516
rect 82780 118476 164516 118504
rect 82780 118464 82786 118476
rect 164510 118464 164516 118476
rect 164568 118464 164574 118516
rect 188982 118464 188988 118516
rect 189040 118504 189046 118516
rect 230658 118504 230664 118516
rect 189040 118476 230664 118504
rect 189040 118464 189046 118476
rect 230658 118464 230664 118476
rect 230716 118464 230722 118516
rect 237282 118464 237288 118516
rect 237340 118504 237346 118516
rect 255314 118504 255320 118516
rect 237340 118476 255320 118504
rect 237340 118464 237346 118476
rect 255314 118464 255320 118476
rect 255372 118464 255378 118516
rect 299290 118464 299296 118516
rect 299348 118504 299354 118516
rect 320358 118504 320364 118516
rect 299348 118476 320364 118504
rect 299348 118464 299354 118476
rect 320358 118464 320364 118476
rect 320416 118464 320422 118516
rect 342162 118464 342168 118516
rect 342220 118504 342226 118516
rect 400950 118504 400956 118516
rect 342220 118476 400956 118504
rect 342220 118464 342226 118476
rect 400950 118464 400956 118476
rect 401008 118464 401014 118516
rect 404262 118464 404268 118516
rect 404320 118504 404326 118516
rect 475378 118504 475384 118516
rect 404320 118476 475384 118504
rect 404320 118464 404326 118476
rect 475378 118464 475384 118476
rect 475436 118464 475442 118516
rect 120718 118396 120724 118448
rect 120776 118436 120782 118448
rect 125686 118436 125692 118448
rect 120776 118408 125692 118436
rect 120776 118396 120782 118408
rect 125686 118396 125692 118408
rect 125744 118436 125750 118448
rect 170030 118436 170036 118448
rect 125744 118408 170036 118436
rect 125744 118396 125750 118408
rect 170030 118396 170036 118408
rect 170088 118396 170094 118448
rect 186222 118396 186228 118448
rect 186280 118436 186286 118448
rect 229462 118436 229468 118448
rect 186280 118408 229468 118436
rect 186280 118396 186286 118408
rect 229462 118396 229468 118408
rect 229520 118396 229526 118448
rect 235902 118396 235908 118448
rect 235960 118436 235966 118448
rect 254578 118436 254584 118448
rect 235960 118408 254584 118436
rect 235960 118396 235966 118408
rect 254578 118396 254584 118408
rect 254636 118396 254642 118448
rect 302142 118396 302148 118448
rect 302200 118436 302206 118448
rect 325878 118436 325884 118448
rect 302200 118408 325884 118436
rect 302200 118396 302206 118408
rect 325878 118396 325884 118408
rect 325936 118396 325942 118448
rect 335998 118396 336004 118448
rect 336056 118436 336062 118448
rect 348418 118436 348424 118448
rect 336056 118408 348424 118436
rect 336056 118396 336062 118408
rect 348418 118396 348424 118408
rect 348476 118396 348482 118448
rect 369670 118396 369676 118448
rect 369728 118436 369734 118448
rect 374638 118436 374644 118448
rect 369728 118408 374644 118436
rect 369728 118396 369734 118408
rect 374638 118396 374644 118408
rect 374696 118396 374702 118448
rect 417418 118396 417424 118448
rect 417476 118436 417482 118448
rect 422846 118436 422852 118448
rect 417476 118408 422852 118436
rect 417476 118396 417482 118408
rect 422846 118396 422852 118408
rect 422904 118396 422910 118448
rect 431770 118396 431776 118448
rect 431828 118436 431834 118448
rect 500218 118436 500224 118448
rect 431828 118408 500224 118436
rect 431828 118396 431834 118408
rect 500218 118396 500224 118408
rect 500276 118396 500282 118448
rect 71590 118328 71596 118380
rect 71648 118368 71654 118380
rect 88334 118368 88340 118380
rect 71648 118340 88340 118368
rect 71648 118328 71654 118340
rect 88334 118328 88340 118340
rect 88392 118328 88398 118380
rect 110322 118328 110328 118380
rect 110380 118368 110386 118380
rect 145558 118368 145564 118380
rect 110380 118340 145564 118368
rect 110380 118328 110386 118340
rect 145558 118328 145564 118340
rect 145616 118328 145622 118380
rect 146846 118328 146852 118380
rect 146904 118368 146910 118380
rect 153470 118368 153476 118380
rect 146904 118340 153476 118368
rect 146904 118328 146910 118340
rect 153470 118328 153476 118340
rect 153528 118328 153534 118380
rect 182174 118328 182180 118380
rect 182232 118368 182238 118380
rect 187786 118368 187792 118380
rect 182232 118340 187792 118368
rect 182232 118328 182238 118340
rect 187786 118328 187792 118340
rect 187844 118328 187850 118380
rect 194502 118328 194508 118380
rect 194560 118368 194566 118380
rect 233234 118368 233240 118380
rect 194560 118340 233240 118368
rect 194560 118328 194566 118340
rect 233234 118328 233240 118340
rect 233292 118328 233298 118380
rect 238110 118368 238116 118380
rect 233344 118340 238116 118368
rect 56502 118260 56508 118312
rect 56560 118300 56566 118312
rect 125870 118300 125876 118312
rect 56560 118272 125876 118300
rect 56560 118260 56566 118272
rect 125870 118260 125876 118272
rect 125928 118300 125934 118312
rect 126882 118300 126888 118312
rect 125928 118272 126888 118300
rect 125928 118260 125934 118272
rect 126882 118260 126888 118272
rect 126940 118260 126946 118312
rect 128906 118260 128912 118312
rect 128964 118300 128970 118312
rect 135438 118300 135444 118312
rect 128964 118272 135444 118300
rect 128964 118260 128970 118272
rect 135438 118260 135444 118272
rect 135496 118300 135502 118312
rect 137186 118300 137192 118312
rect 135496 118272 137192 118300
rect 135496 118260 135502 118272
rect 137186 118260 137192 118272
rect 137244 118260 137250 118312
rect 137278 118260 137284 118312
rect 137336 118300 137342 118312
rect 182910 118300 182916 118312
rect 137336 118272 182916 118300
rect 137336 118260 137342 118272
rect 182910 118260 182916 118272
rect 182968 118260 182974 118312
rect 183462 118260 183468 118312
rect 183520 118300 183526 118312
rect 227714 118300 227720 118312
rect 183520 118272 227720 118300
rect 183520 118260 183526 118272
rect 227714 118260 227720 118272
rect 227772 118260 227778 118312
rect 231118 118260 231124 118312
rect 231176 118300 231182 118312
rect 233344 118300 233372 118340
rect 238110 118328 238116 118340
rect 238168 118328 238174 118380
rect 238662 118328 238668 118380
rect 238720 118368 238726 118380
rect 256694 118368 256700 118380
rect 238720 118340 256700 118368
rect 238720 118328 238726 118340
rect 256694 118328 256700 118340
rect 256752 118328 256758 118380
rect 260742 118328 260748 118380
rect 260800 118368 260806 118380
rect 267734 118368 267740 118380
rect 260800 118340 267740 118368
rect 260800 118328 260806 118340
rect 267734 118328 267740 118340
rect 267792 118328 267798 118380
rect 304166 118328 304172 118380
rect 304224 118368 304230 118380
rect 330018 118368 330024 118380
rect 304224 118340 330024 118368
rect 304224 118328 304230 118340
rect 330018 118328 330024 118340
rect 330076 118328 330082 118380
rect 338482 118328 338488 118380
rect 338540 118368 338546 118380
rect 396258 118368 396264 118380
rect 338540 118340 396264 118368
rect 338540 118328 338546 118340
rect 396258 118328 396264 118340
rect 396316 118328 396322 118380
rect 400858 118328 400864 118380
rect 400916 118368 400922 118380
rect 473998 118368 474004 118380
rect 400916 118340 474004 118368
rect 400916 118328 400922 118340
rect 473998 118328 474004 118340
rect 474056 118328 474062 118380
rect 231176 118272 233372 118300
rect 231176 118260 231182 118272
rect 237190 118260 237196 118312
rect 237248 118300 237254 118312
rect 255774 118300 255780 118312
rect 237248 118272 255780 118300
rect 237248 118260 237254 118272
rect 255774 118260 255780 118272
rect 255832 118260 255838 118312
rect 256602 118260 256608 118312
rect 256660 118300 256666 118312
rect 265526 118300 265532 118312
rect 256660 118272 265532 118300
rect 256660 118260 256666 118272
rect 265526 118260 265532 118272
rect 265584 118260 265590 118312
rect 306006 118260 306012 118312
rect 306064 118300 306070 118312
rect 332870 118300 332876 118312
rect 306064 118272 332876 118300
rect 306064 118260 306070 118272
rect 332870 118260 332876 118272
rect 332928 118260 332934 118312
rect 337838 118260 337844 118312
rect 337896 118300 337902 118312
rect 351178 118300 351184 118312
rect 337896 118272 351184 118300
rect 337896 118260 337902 118272
rect 351178 118260 351184 118272
rect 351236 118260 351242 118312
rect 362310 118260 362316 118312
rect 362368 118300 362374 118312
rect 442994 118300 443000 118312
rect 362368 118272 443000 118300
rect 362368 118260 362374 118272
rect 442994 118260 443000 118272
rect 443052 118260 443058 118312
rect 31662 118192 31668 118244
rect 31720 118232 31726 118244
rect 107562 118232 107568 118244
rect 31720 118204 107568 118232
rect 31720 118192 31726 118204
rect 107562 118192 107568 118204
rect 107620 118192 107626 118244
rect 113082 118192 113088 118244
rect 113140 118232 113146 118244
rect 175550 118232 175556 118244
rect 113140 118204 175556 118232
rect 113140 118192 113146 118204
rect 175550 118192 175556 118204
rect 175608 118192 175614 118244
rect 184842 118192 184848 118244
rect 184900 118232 184906 118244
rect 229186 118232 229192 118244
rect 184900 118204 229192 118232
rect 184900 118192 184906 118204
rect 229186 118192 229192 118204
rect 229244 118192 229250 118244
rect 233142 118192 233148 118244
rect 233200 118232 233206 118244
rect 253290 118232 253296 118244
rect 233200 118204 253296 118232
rect 233200 118192 233206 118204
rect 253290 118192 253296 118204
rect 253348 118192 253354 118244
rect 253842 118192 253848 118244
rect 253900 118232 253906 118244
rect 263686 118232 263692 118244
rect 253900 118204 263692 118232
rect 253900 118192 253906 118204
rect 263686 118192 263692 118204
rect 263744 118192 263750 118244
rect 300486 118192 300492 118244
rect 300544 118232 300550 118244
rect 300544 118204 307064 118232
rect 300544 118192 300550 118204
rect 28902 118124 28908 118176
rect 28960 118164 28966 118176
rect 114462 118164 114468 118176
rect 28960 118136 114468 118164
rect 28960 118124 28966 118136
rect 114462 118124 114468 118136
rect 114520 118124 114526 118176
rect 129274 118124 129280 118176
rect 129332 118164 129338 118176
rect 177390 118164 177396 118176
rect 129332 118136 177396 118164
rect 129332 118124 129338 118136
rect 177390 118124 177396 118136
rect 177448 118124 177454 118176
rect 179322 118124 179328 118176
rect 179380 118164 179386 118176
rect 225782 118164 225788 118176
rect 179380 118136 225788 118164
rect 179380 118124 179386 118136
rect 225782 118124 225788 118136
rect 225840 118124 225846 118176
rect 234522 118124 234528 118176
rect 234580 118164 234586 118176
rect 253934 118164 253940 118176
rect 234580 118136 253940 118164
rect 234580 118124 234586 118136
rect 253934 118124 253940 118136
rect 253992 118124 253998 118176
rect 257982 118124 257988 118176
rect 258040 118164 258046 118176
rect 266354 118164 266360 118176
rect 258040 118136 266360 118164
rect 258040 118124 258046 118136
rect 266354 118124 266360 118136
rect 266412 118124 266418 118176
rect 267642 118124 267648 118176
rect 267700 118164 267706 118176
rect 271046 118164 271052 118176
rect 267700 118136 271052 118164
rect 267700 118124 267706 118136
rect 271046 118124 271052 118136
rect 271104 118124 271110 118176
rect 291102 118124 291108 118176
rect 291160 118164 291166 118176
rect 305178 118164 305184 118176
rect 291160 118136 305184 118164
rect 291160 118124 291166 118136
rect 305178 118124 305184 118136
rect 305236 118124 305242 118176
rect 307036 118164 307064 118204
rect 307662 118192 307668 118244
rect 307720 118232 307726 118244
rect 336918 118232 336924 118244
rect 307720 118204 336924 118232
rect 307720 118192 307726 118204
rect 336918 118192 336924 118204
rect 336976 118192 336982 118244
rect 339402 118192 339408 118244
rect 339460 118232 339466 118244
rect 353938 118232 353944 118244
rect 339460 118204 353944 118232
rect 339460 118192 339466 118204
rect 353938 118192 353944 118204
rect 353996 118192 354002 118244
rect 356790 118192 356796 118244
rect 356848 118232 356854 118244
rect 356848 118204 365116 118232
rect 356848 118192 356854 118204
rect 307036 118136 308168 118164
rect 23382 118056 23388 118108
rect 23440 118096 23446 118108
rect 110322 118096 110328 118108
rect 23440 118068 110328 118096
rect 23440 118056 23446 118068
rect 110322 118056 110328 118068
rect 110380 118056 110386 118108
rect 115198 118056 115204 118108
rect 115256 118096 115262 118108
rect 126974 118096 126980 118108
rect 115256 118068 126980 118096
rect 115256 118056 115262 118068
rect 126974 118056 126980 118068
rect 127032 118056 127038 118108
rect 128170 118056 128176 118108
rect 128228 118096 128234 118108
rect 133138 118096 133144 118108
rect 128228 118068 133144 118096
rect 128228 118056 128234 118068
rect 133138 118056 133144 118068
rect 133196 118056 133202 118108
rect 133230 118056 133236 118108
rect 133288 118096 133294 118108
rect 173894 118096 173900 118108
rect 133288 118068 173900 118096
rect 133288 118056 133294 118068
rect 173894 118056 173900 118068
rect 173952 118056 173958 118108
rect 176562 118056 176568 118108
rect 176620 118096 176626 118108
rect 223942 118096 223948 118108
rect 176620 118068 223948 118096
rect 176620 118056 176626 118068
rect 223942 118056 223948 118068
rect 224000 118056 224006 118108
rect 231762 118056 231768 118108
rect 231820 118096 231826 118108
rect 252738 118096 252744 118108
rect 231820 118068 252744 118096
rect 231820 118056 231826 118068
rect 252738 118056 252744 118068
rect 252796 118056 252802 118108
rect 255222 118056 255228 118108
rect 255280 118096 255286 118108
rect 264974 118096 264980 118108
rect 255280 118068 264980 118096
rect 255280 118056 255286 118068
rect 264974 118056 264980 118068
rect 265032 118056 265038 118108
rect 293126 118056 293132 118108
rect 293184 118096 293190 118108
rect 307938 118096 307944 118108
rect 293184 118068 307944 118096
rect 293184 118056 293190 118068
rect 307938 118056 307944 118068
rect 307996 118056 308002 118108
rect 60642 117988 60648 118040
rect 60700 118028 60706 118040
rect 82722 118028 82728 118040
rect 60700 118000 82728 118028
rect 60700 117988 60706 118000
rect 82722 117988 82728 118000
rect 82780 117988 82786 118040
rect 88334 117988 88340 118040
rect 88392 118028 88398 118040
rect 179414 118028 179420 118040
rect 88392 118000 179420 118028
rect 88392 117988 88398 118000
rect 179414 117988 179420 118000
rect 179472 117988 179478 118040
rect 182082 117988 182088 118040
rect 182140 118028 182146 118040
rect 226978 118028 226984 118040
rect 182140 118000 226984 118028
rect 182140 117988 182146 118000
rect 226978 117988 226984 118000
rect 227036 117988 227042 118040
rect 229002 117988 229008 118040
rect 229060 118028 229066 118040
rect 251266 118028 251272 118040
rect 229060 118000 251272 118028
rect 229060 117988 229066 118000
rect 251266 117988 251272 118000
rect 251324 117988 251330 118040
rect 253750 117988 253756 118040
rect 253808 118028 253814 118040
rect 264330 118028 264336 118040
rect 253808 118000 264336 118028
rect 253808 117988 253814 118000
rect 264330 117988 264336 118000
rect 264388 117988 264394 118040
rect 266262 117988 266268 118040
rect 266320 118028 266326 118040
rect 270494 118028 270500 118040
rect 266320 118000 270500 118028
rect 266320 117988 266326 118000
rect 270494 117988 270500 118000
rect 270552 117988 270558 118040
rect 294966 117988 294972 118040
rect 295024 118028 295030 118040
rect 295024 118000 306144 118028
rect 295024 117988 295030 118000
rect 9582 117920 9588 117972
rect 9640 117960 9646 117972
rect 69842 117960 69848 117972
rect 9640 117932 69848 117960
rect 9640 117920 9646 117932
rect 69842 117920 69848 117932
rect 69900 117920 69906 117972
rect 122834 117920 122840 117972
rect 122892 117960 122898 117972
rect 122892 117932 166396 117960
rect 122892 117920 122898 117932
rect 107562 117852 107568 117904
rect 107620 117892 107626 117904
rect 149882 117892 149888 117904
rect 107620 117864 149888 117892
rect 107620 117852 107626 117864
rect 149882 117852 149888 117864
rect 149940 117852 149946 117904
rect 96522 117784 96528 117836
rect 96580 117824 96586 117836
rect 99190 117824 99196 117836
rect 96580 117796 99196 117824
rect 96580 117784 96586 117796
rect 99190 117784 99196 117796
rect 99248 117784 99254 117836
rect 122098 117784 122104 117836
rect 122156 117824 122162 117836
rect 122650 117824 122656 117836
rect 122156 117796 122656 117824
rect 122156 117784 122162 117796
rect 122650 117784 122656 117796
rect 122708 117824 122714 117836
rect 160830 117824 160836 117836
rect 122708 117796 160836 117824
rect 122708 117784 122714 117796
rect 160830 117784 160836 117796
rect 160888 117784 160894 117836
rect 71682 117716 71688 117768
rect 71740 117756 71746 117768
rect 73798 117756 73804 117768
rect 71740 117728 73804 117756
rect 71740 117716 71746 117728
rect 73798 117716 73804 117728
rect 73856 117756 73862 117768
rect 79962 117756 79968 117768
rect 73856 117728 79968 117756
rect 73856 117716 73862 117728
rect 79962 117716 79968 117728
rect 80020 117716 80026 117768
rect 99466 117716 99472 117768
rect 99524 117756 99530 117768
rect 122834 117756 122840 117768
rect 99524 117728 108988 117756
rect 99524 117716 99530 117728
rect 80146 117648 80152 117700
rect 80204 117688 80210 117700
rect 86954 117688 86960 117700
rect 80204 117660 86960 117688
rect 80204 117648 80210 117660
rect 86954 117648 86960 117660
rect 87012 117648 87018 117700
rect 108960 117688 108988 117728
rect 109052 117728 122840 117756
rect 109052 117688 109080 117728
rect 122834 117716 122840 117728
rect 122892 117716 122898 117768
rect 126882 117716 126888 117768
rect 126940 117756 126946 117768
rect 162854 117756 162860 117768
rect 126940 117728 162860 117756
rect 126940 117716 126946 117728
rect 162854 117716 162860 117728
rect 162912 117716 162918 117768
rect 108960 117660 109080 117688
rect 127618 117648 127624 117700
rect 127676 117688 127682 117700
rect 128170 117688 128176 117700
rect 127676 117660 128176 117688
rect 127676 117648 127682 117660
rect 128170 117648 128176 117660
rect 128228 117648 128234 117700
rect 129090 117648 129096 117700
rect 129148 117688 129154 117700
rect 129366 117688 129372 117700
rect 129148 117660 129372 117688
rect 129148 117648 129154 117660
rect 129366 117648 129372 117660
rect 129424 117688 129430 117700
rect 137278 117688 137284 117700
rect 129424 117660 137284 117688
rect 129424 117648 129430 117660
rect 137278 117648 137284 117660
rect 137336 117648 137342 117700
rect 137388 117660 137600 117688
rect 130470 117580 130476 117632
rect 130528 117620 130534 117632
rect 137388 117620 137416 117660
rect 130528 117592 137416 117620
rect 137572 117620 137600 117660
rect 137646 117648 137652 117700
rect 137704 117688 137710 117700
rect 166258 117688 166264 117700
rect 137704 117660 166264 117688
rect 137704 117648 137710 117660
rect 166258 117648 166264 117660
rect 166316 117648 166322 117700
rect 158990 117620 158996 117632
rect 137572 117592 158996 117620
rect 130528 117580 130534 117592
rect 158990 117580 158996 117592
rect 159048 117580 159054 117632
rect 166368 117620 166396 117932
rect 177942 117920 177948 117972
rect 178000 117960 178006 117972
rect 225138 117960 225144 117972
rect 178000 117932 225144 117960
rect 178000 117920 178006 117932
rect 225138 117920 225144 117932
rect 225196 117920 225202 117972
rect 226242 117920 226248 117972
rect 226300 117960 226306 117972
rect 239398 117960 239404 117972
rect 226300 117932 239404 117960
rect 226300 117920 226306 117932
rect 239398 117920 239404 117932
rect 239456 117920 239462 117972
rect 241698 117960 241704 117972
rect 239508 117932 241704 117960
rect 197262 117852 197268 117904
rect 197320 117892 197326 117904
rect 234982 117892 234988 117904
rect 197320 117864 234988 117892
rect 197320 117852 197326 117864
rect 234982 117852 234988 117864
rect 235040 117852 235046 117904
rect 238110 117852 238116 117904
rect 238168 117892 238174 117904
rect 239508 117892 239536 117932
rect 241698 117920 241704 117932
rect 241756 117920 241762 117972
rect 251082 117920 251088 117972
rect 251140 117960 251146 117972
rect 262490 117960 262496 117972
rect 251140 117932 262496 117960
rect 251140 117920 251146 117932
rect 262490 117920 262496 117932
rect 262548 117920 262554 117972
rect 264882 117920 264888 117972
rect 264940 117960 264946 117972
rect 269850 117960 269856 117972
rect 264940 117932 269856 117960
rect 264940 117920 264946 117932
rect 269850 117920 269856 117932
rect 269908 117920 269914 117972
rect 279050 117920 279056 117972
rect 279108 117960 279114 117972
rect 280338 117960 280344 117972
rect 279108 117932 280344 117960
rect 279108 117920 279114 117932
rect 280338 117920 280344 117932
rect 280396 117920 280402 117972
rect 280890 117920 280896 117972
rect 280948 117960 280954 117972
rect 281442 117960 281448 117972
rect 280948 117932 281448 117960
rect 280948 117920 280954 117932
rect 281442 117920 281448 117932
rect 281500 117920 281506 117972
rect 238168 117864 239536 117892
rect 238168 117852 238174 117864
rect 241422 117852 241428 117904
rect 241480 117892 241486 117904
rect 257614 117892 257620 117904
rect 241480 117864 257620 117892
rect 241480 117852 241486 117864
rect 257614 117852 257620 117864
rect 257672 117852 257678 117904
rect 263502 117852 263508 117904
rect 263560 117892 263566 117904
rect 268654 117892 268660 117904
rect 263560 117864 268660 117892
rect 263560 117852 263566 117864
rect 268654 117852 268660 117864
rect 268712 117852 268718 117904
rect 296530 117852 296536 117904
rect 296588 117892 296594 117904
rect 306116 117892 306144 118000
rect 308140 117960 308168 118136
rect 316678 118124 316684 118176
rect 316736 118164 316742 118176
rect 339678 118164 339684 118176
rect 316736 118136 339684 118164
rect 316736 118124 316742 118136
rect 339678 118124 339684 118136
rect 339736 118124 339742 118176
rect 359274 118124 359280 118176
rect 359332 118164 359338 118176
rect 360102 118164 360108 118176
rect 359332 118136 360108 118164
rect 359332 118124 359338 118136
rect 360102 118124 360108 118136
rect 360160 118124 360166 118176
rect 316586 118056 316592 118108
rect 316644 118096 316650 118108
rect 343910 118096 343916 118108
rect 316644 118068 343916 118096
rect 316644 118056 316650 118068
rect 343910 118056 343916 118068
rect 343968 118056 343974 118108
rect 354950 118056 354956 118108
rect 355008 118096 355014 118108
rect 364978 118096 364984 118108
rect 355008 118068 364984 118096
rect 355008 118056 355014 118068
rect 364978 118056 364984 118068
rect 365036 118056 365042 118108
rect 365088 118096 365116 118204
rect 365990 118192 365996 118244
rect 366048 118232 366054 118244
rect 449894 118232 449900 118244
rect 366048 118204 449900 118232
rect 366048 118192 366054 118204
rect 449894 118192 449900 118204
rect 449952 118192 449958 118244
rect 374638 118124 374644 118176
rect 374696 118164 374702 118176
rect 456794 118164 456800 118176
rect 374696 118136 456800 118164
rect 374696 118124 374702 118136
rect 456794 118124 456800 118136
rect 456852 118124 456858 118176
rect 365088 118068 372292 118096
rect 313182 117988 313188 118040
rect 313240 118028 313246 118040
rect 347958 118028 347964 118040
rect 313240 118000 347964 118028
rect 313240 117988 313246 118000
rect 347958 117988 347964 118000
rect 348016 117988 348022 118040
rect 372264 118028 372292 118068
rect 373350 118056 373356 118108
rect 373408 118096 373414 118108
rect 463694 118096 463700 118108
rect 373408 118068 463700 118096
rect 373408 118056 373414 118068
rect 463694 118056 463700 118068
rect 463752 118056 463758 118108
rect 374638 118028 374644 118040
rect 372264 118000 374644 118028
rect 374638 117988 374644 118000
rect 374696 117988 374702 118040
rect 377030 117988 377036 118040
rect 377088 118028 377094 118040
rect 470594 118028 470600 118040
rect 377088 118000 470600 118028
rect 377088 117988 377094 118000
rect 470594 117988 470600 118000
rect 470652 117988 470658 118040
rect 321738 117960 321744 117972
rect 308140 117932 321744 117960
rect 321738 117920 321744 117932
rect 321796 117920 321802 117972
rect 380710 117920 380716 117972
rect 380768 117960 380774 117972
rect 477494 117960 477500 117972
rect 380768 117932 477500 117960
rect 380768 117920 380774 117932
rect 477494 117920 477500 117932
rect 477552 117920 477558 117972
rect 311894 117892 311900 117904
rect 296588 117864 302372 117892
rect 306116 117864 311900 117892
rect 296588 117852 296594 117864
rect 167730 117784 167736 117836
rect 167788 117824 167794 117836
rect 189074 117824 189080 117836
rect 167788 117796 189080 117824
rect 167788 117784 167794 117796
rect 189074 117784 189080 117796
rect 189132 117784 189138 117836
rect 213822 117784 213828 117836
rect 213880 117824 213886 117836
rect 243630 117824 243636 117836
rect 213880 117796 243636 117824
rect 213880 117784 213886 117796
rect 243630 117784 243636 117796
rect 243688 117784 243694 117836
rect 245746 117784 245752 117836
rect 245804 117824 245810 117836
rect 260006 117824 260012 117836
rect 245804 117796 260012 117824
rect 245804 117784 245810 117796
rect 260006 117784 260012 117796
rect 260064 117784 260070 117836
rect 263410 117784 263416 117836
rect 263468 117824 263474 117836
rect 269206 117824 269212 117836
rect 263468 117796 269212 117824
rect 263468 117784 263474 117796
rect 269206 117784 269212 117796
rect 269264 117784 269270 117836
rect 296162 117784 296168 117836
rect 296220 117824 296226 117836
rect 296220 117796 302280 117824
rect 296220 117784 296226 117796
rect 191098 117716 191104 117768
rect 191156 117756 191162 117768
rect 205174 117756 205180 117768
rect 191156 117728 205180 117756
rect 191156 117716 191162 117728
rect 205174 117716 205180 117728
rect 205232 117716 205238 117768
rect 217962 117716 217968 117768
rect 218020 117756 218026 117768
rect 245654 117756 245660 117768
rect 218020 117728 245660 117756
rect 218020 117716 218026 117728
rect 245654 117716 245660 117728
rect 245712 117716 245718 117768
rect 246942 117716 246948 117768
rect 247000 117756 247006 117768
rect 260834 117756 260840 117768
rect 247000 117728 260840 117756
rect 247000 117716 247006 117728
rect 260834 117716 260840 117728
rect 260892 117716 260898 117768
rect 262122 117716 262128 117768
rect 262180 117756 262186 117768
rect 268010 117756 268016 117768
rect 262180 117728 268016 117756
rect 262180 117716 262186 117728
rect 268010 117716 268016 117728
rect 268068 117716 268074 117768
rect 277854 117716 277860 117768
rect 277912 117756 277918 117768
rect 278682 117756 278688 117768
rect 277912 117728 278688 117756
rect 277912 117716 277918 117728
rect 278682 117716 278688 117728
rect 278740 117716 278746 117768
rect 169018 117648 169024 117700
rect 169076 117688 169082 117700
rect 192662 117688 192668 117700
rect 169076 117660 192668 117688
rect 169076 117648 169082 117660
rect 192662 117648 192668 117660
rect 192720 117648 192726 117700
rect 213178 117648 213184 117700
rect 213236 117688 213242 117700
rect 232498 117688 232504 117700
rect 213236 117660 232504 117688
rect 213236 117648 213242 117660
rect 232498 117648 232504 117660
rect 232556 117648 232562 117700
rect 233878 117648 233884 117700
rect 233936 117688 233942 117700
rect 244274 117688 244280 117700
rect 233936 117660 244280 117688
rect 233936 117648 233942 117660
rect 244274 117648 244280 117660
rect 244332 117648 244338 117700
rect 245562 117648 245568 117700
rect 245620 117688 245626 117700
rect 259454 117688 259460 117700
rect 245620 117660 259460 117688
rect 245620 117648 245626 117660
rect 259454 117648 259460 117660
rect 259512 117648 259518 117700
rect 302252 117688 302280 117796
rect 302344 117756 302372 117864
rect 311894 117852 311900 117864
rect 311952 117852 311958 117904
rect 314562 117852 314568 117904
rect 314620 117892 314626 117904
rect 322198 117892 322204 117904
rect 314620 117864 322204 117892
rect 314620 117852 314626 117864
rect 322198 117852 322204 117864
rect 322256 117852 322262 117904
rect 331858 117892 331864 117904
rect 322308 117864 331864 117892
rect 316402 117784 316408 117836
rect 316460 117824 316466 117836
rect 322308 117824 322336 117864
rect 331858 117852 331864 117864
rect 331916 117852 331922 117904
rect 345842 117852 345848 117904
rect 345900 117892 345906 117904
rect 407758 117892 407764 117904
rect 345900 117864 407764 117892
rect 345900 117852 345906 117864
rect 407758 117852 407764 117864
rect 407816 117852 407822 117904
rect 420822 117852 420828 117904
rect 420880 117892 420886 117904
rect 489178 117892 489184 117904
rect 420880 117864 489184 117892
rect 420880 117852 420886 117864
rect 489178 117852 489184 117864
rect 489236 117852 489242 117904
rect 316460 117796 322336 117824
rect 316460 117784 316466 117796
rect 331122 117784 331128 117836
rect 331180 117824 331186 117836
rect 337378 117824 337384 117836
rect 331180 117796 337384 117824
rect 331180 117784 331186 117796
rect 337378 117784 337384 117796
rect 337436 117784 337442 117836
rect 369688 117796 369992 117824
rect 314654 117756 314660 117768
rect 302344 117728 314660 117756
rect 314654 117716 314660 117728
rect 314712 117716 314718 117768
rect 315206 117716 315212 117768
rect 315264 117756 315270 117768
rect 315942 117756 315948 117768
rect 315264 117728 315948 117756
rect 315264 117716 315270 117728
rect 315942 117716 315948 117728
rect 316000 117716 316006 117768
rect 320726 117716 320732 117768
rect 320784 117756 320790 117768
rect 321370 117756 321376 117768
rect 320784 117728 321376 117756
rect 320784 117716 320790 117728
rect 321370 117716 321376 117728
rect 321428 117716 321434 117768
rect 321922 117716 321928 117768
rect 321980 117756 321986 117768
rect 357986 117756 357992 117768
rect 321980 117728 357992 117756
rect 321980 117716 321986 117728
rect 357986 117716 357992 117728
rect 358044 117716 358050 117768
rect 302252 117660 303476 117688
rect 171870 117620 171876 117632
rect 166368 117592 171876 117620
rect 171870 117580 171876 117592
rect 171928 117580 171934 117632
rect 196618 117580 196624 117632
rect 196676 117620 196682 117632
rect 211706 117620 211712 117632
rect 196676 117592 211712 117620
rect 196676 117580 196682 117592
rect 211706 117580 211712 117592
rect 211764 117580 211770 117632
rect 224218 117580 224224 117632
rect 224276 117620 224282 117632
rect 236822 117620 236828 117632
rect 224276 117592 236828 117620
rect 224276 117580 224282 117592
rect 236822 117580 236828 117592
rect 236880 117580 236886 117632
rect 237282 117580 237288 117632
rect 237340 117620 237346 117632
rect 240410 117620 240416 117632
rect 237340 117592 240416 117620
rect 237340 117580 237346 117592
rect 240410 117580 240416 117592
rect 240468 117580 240474 117632
rect 244182 117580 244188 117632
rect 244240 117620 244246 117632
rect 258810 117620 258816 117632
rect 244240 117592 258816 117620
rect 244240 117580 244246 117592
rect 258810 117580 258816 117592
rect 258868 117580 258874 117632
rect 259270 117580 259276 117632
rect 259328 117620 259334 117632
rect 263134 117620 263140 117632
rect 259328 117592 263140 117620
rect 259328 117580 259334 117592
rect 263134 117580 263140 117592
rect 263192 117580 263198 117632
rect 86954 117512 86960 117564
rect 87012 117552 87018 117564
rect 96522 117552 96528 117564
rect 87012 117524 96528 117552
rect 87012 117512 87018 117524
rect 96522 117512 96528 117524
rect 96580 117512 96586 117564
rect 128814 117512 128820 117564
rect 128872 117552 128878 117564
rect 137646 117552 137652 117564
rect 128872 117524 137652 117552
rect 128872 117512 128878 117524
rect 137646 117512 137652 117524
rect 137704 117512 137710 117564
rect 138658 117512 138664 117564
rect 138716 117552 138722 117564
rect 139394 117552 139400 117564
rect 138716 117524 139400 117552
rect 138716 117512 138722 117524
rect 139394 117512 139400 117524
rect 139452 117552 139458 117564
rect 146754 117552 146760 117564
rect 139452 117524 146760 117552
rect 139452 117512 139458 117524
rect 146754 117512 146760 117524
rect 146812 117512 146818 117564
rect 235258 117512 235264 117564
rect 235316 117552 235322 117564
rect 247770 117552 247776 117564
rect 235316 117524 247776 117552
rect 235316 117512 235322 117524
rect 247770 117512 247776 117524
rect 247828 117512 247834 117564
rect 248322 117512 248328 117564
rect 248380 117552 248386 117564
rect 261294 117552 261300 117564
rect 248380 117524 261300 117552
rect 248380 117512 248386 117524
rect 261294 117512 261300 117524
rect 261352 117512 261358 117564
rect 67542 117444 67548 117496
rect 67600 117484 67606 117496
rect 71038 117484 71044 117496
rect 67600 117456 71044 117484
rect 67600 117444 67606 117456
rect 71038 117444 71044 117456
rect 71096 117484 71102 117496
rect 168374 117484 168380 117496
rect 71096 117456 168380 117484
rect 71096 117444 71102 117456
rect 168374 117444 168380 117456
rect 168432 117444 168438 117496
rect 229738 117444 229744 117496
rect 229796 117484 229802 117496
rect 238846 117484 238852 117496
rect 229796 117456 238852 117484
rect 229796 117444 229802 117456
rect 238846 117444 238852 117456
rect 238904 117444 238910 117496
rect 240226 117484 240232 117496
rect 238956 117456 240232 117484
rect 114462 117376 114468 117428
rect 114520 117416 114526 117428
rect 148042 117416 148048 117428
rect 114520 117388 148048 117416
rect 114520 117376 114526 117388
rect 148042 117376 148048 117388
rect 148100 117376 148106 117428
rect 182174 117376 182180 117428
rect 182232 117416 182238 117428
rect 186498 117416 186504 117428
rect 182232 117388 186504 117416
rect 182232 117376 182238 117388
rect 186498 117376 186504 117388
rect 186556 117376 186562 117428
rect 232498 117376 232504 117428
rect 232556 117416 232562 117428
rect 232556 117388 237420 117416
rect 232556 117376 232562 117388
rect 92382 117308 92388 117360
rect 92440 117348 92446 117360
rect 97902 117348 97908 117360
rect 92440 117320 97908 117348
rect 92440 117308 92446 117320
rect 97902 117308 97908 117320
rect 97960 117308 97966 117360
rect 109678 117308 109684 117360
rect 109736 117348 109742 117360
rect 113082 117348 113088 117360
rect 109736 117320 113088 117348
rect 109736 117308 109742 117320
rect 113082 117308 113088 117320
rect 113140 117308 113146 117360
rect 133138 117308 133144 117360
rect 133196 117348 133202 117360
rect 190454 117348 190460 117360
rect 133196 117320 190460 117348
rect 133196 117308 133202 117320
rect 190454 117308 190460 117320
rect 190512 117308 190518 117360
rect 190546 117308 190552 117360
rect 190604 117348 190610 117360
rect 192110 117348 192116 117360
rect 190604 117320 192116 117348
rect 190604 117308 190610 117320
rect 192110 117308 192116 117320
rect 192168 117308 192174 117360
rect 225598 117308 225604 117360
rect 225656 117348 225662 117360
rect 231302 117348 231308 117360
rect 225656 117320 231308 117348
rect 225656 117308 225662 117320
rect 231302 117308 231308 117320
rect 231360 117308 231366 117360
rect 232590 117308 232596 117360
rect 232648 117348 232654 117360
rect 237282 117348 237288 117360
rect 232648 117320 237288 117348
rect 232648 117308 232654 117320
rect 237282 117308 237288 117320
rect 237340 117308 237346 117360
rect 237392 117348 237420 117388
rect 238956 117348 238984 117456
rect 240226 117444 240232 117456
rect 240284 117444 240290 117496
rect 243538 117444 243544 117496
rect 243596 117484 243602 117496
rect 249058 117484 249064 117496
rect 243596 117456 249064 117484
rect 243596 117444 243602 117456
rect 249058 117444 249064 117456
rect 249116 117444 249122 117496
rect 249702 117444 249708 117496
rect 249760 117484 249766 117496
rect 262214 117484 262220 117496
rect 249760 117456 262220 117484
rect 249760 117444 249766 117456
rect 262214 117444 262220 117456
rect 262272 117444 262278 117496
rect 271782 117444 271788 117496
rect 271840 117484 271846 117496
rect 273254 117484 273260 117496
rect 271840 117456 273260 117484
rect 271840 117444 271846 117456
rect 273254 117444 273260 117456
rect 273312 117444 273318 117496
rect 303448 117484 303476 117660
rect 305362 117648 305368 117700
rect 305420 117688 305426 117700
rect 312630 117688 312636 117700
rect 305420 117660 312636 117688
rect 305420 117648 305426 117660
rect 312630 117648 312636 117660
rect 312688 117648 312694 117700
rect 312722 117648 312728 117700
rect 312780 117688 312786 117700
rect 319346 117688 319352 117700
rect 312780 117660 319352 117688
rect 312780 117648 312786 117660
rect 319346 117648 319352 117660
rect 319404 117648 319410 117700
rect 320082 117648 320088 117700
rect 320140 117688 320146 117700
rect 320140 117660 324544 117688
rect 320140 117648 320146 117660
rect 308490 117580 308496 117632
rect 308548 117620 308554 117632
rect 308950 117620 308956 117632
rect 308548 117592 308956 117620
rect 308548 117580 308554 117592
rect 308950 117580 308956 117592
rect 309008 117580 309014 117632
rect 311526 117580 311532 117632
rect 311584 117620 311590 117632
rect 316586 117620 316592 117632
rect 311584 117592 316592 117620
rect 311584 117580 311590 117592
rect 316586 117580 316592 117592
rect 316644 117580 316650 117632
rect 324516 117620 324544 117660
rect 360470 117648 360476 117700
rect 360528 117688 360534 117700
rect 369688 117688 369716 117796
rect 360528 117660 369716 117688
rect 369964 117688 369992 117796
rect 422846 117784 422852 117836
rect 422904 117824 422910 117836
rect 486418 117824 486424 117836
rect 422904 117796 486424 117824
rect 422904 117784 422910 117796
rect 486418 117784 486424 117796
rect 486476 117784 486482 117836
rect 394694 117716 394700 117768
rect 394752 117716 394758 117768
rect 394878 117716 394884 117768
rect 394936 117756 394942 117768
rect 394936 117728 404400 117756
rect 394936 117716 394942 117728
rect 380250 117688 380256 117700
rect 369964 117660 380256 117688
rect 360528 117648 360534 117660
rect 380250 117648 380256 117660
rect 380308 117648 380314 117700
rect 393222 117648 393228 117700
rect 393280 117688 393286 117700
rect 394712 117688 394740 117716
rect 404372 117700 404400 117728
rect 411898 117716 411904 117768
rect 411956 117756 411962 117768
rect 480898 117756 480904 117768
rect 411956 117728 480904 117756
rect 411956 117716 411962 117728
rect 480898 117716 480904 117728
rect 480956 117716 480962 117768
rect 393280 117660 394740 117688
rect 393280 117648 393286 117660
rect 404354 117648 404360 117700
rect 404412 117648 404418 117700
rect 415302 117648 415308 117700
rect 415360 117688 415366 117700
rect 482278 117688 482284 117700
rect 415360 117660 482284 117688
rect 415360 117648 415366 117660
rect 482278 117648 482284 117660
rect 482336 117648 482342 117700
rect 331950 117620 331956 117632
rect 324516 117592 331956 117620
rect 331950 117580 331956 117592
rect 332008 117580 332014 117632
rect 353110 117580 353116 117632
rect 353168 117620 353174 117632
rect 425330 117620 425336 117632
rect 353168 117592 425336 117620
rect 353168 117580 353174 117592
rect 425330 117580 425336 117592
rect 425388 117580 425394 117632
rect 428458 117580 428464 117632
rect 428516 117620 428522 117632
rect 496078 117620 496084 117632
rect 428516 117592 496084 117620
rect 428516 117580 428522 117592
rect 496078 117580 496084 117592
rect 496136 117580 496142 117632
rect 307202 117512 307208 117564
rect 307260 117552 307266 117564
rect 307260 117524 307892 117552
rect 307260 117512 307266 117524
rect 307864 117484 307892 117524
rect 309686 117512 309692 117564
rect 309744 117552 309750 117564
rect 316678 117552 316684 117564
rect 309744 117524 316684 117552
rect 309744 117512 309750 117524
rect 316678 117512 316684 117524
rect 316736 117512 316742 117564
rect 419258 117512 419264 117564
rect 419316 117552 419322 117564
rect 420178 117552 420184 117564
rect 419316 117524 420184 117552
rect 419316 117512 419322 117524
rect 420178 117512 420184 117524
rect 420236 117512 420242 117564
rect 430298 117512 430304 117564
rect 430356 117552 430362 117564
rect 431218 117552 431224 117564
rect 430356 117524 431224 117552
rect 430356 117512 430362 117524
rect 431218 117512 431224 117524
rect 431276 117512 431282 117564
rect 314102 117484 314108 117496
rect 303448 117456 307800 117484
rect 307864 117456 314108 117484
rect 242158 117376 242164 117428
rect 242216 117416 242222 117428
rect 247218 117416 247224 117428
rect 242216 117388 247224 117416
rect 242216 117376 242222 117388
rect 247218 117376 247224 117388
rect 247276 117376 247282 117428
rect 269022 117376 269028 117428
rect 269080 117416 269086 117428
rect 271874 117416 271880 117428
rect 269080 117388 271880 117416
rect 269080 117376 269086 117388
rect 271874 117376 271880 117388
rect 271932 117376 271938 117428
rect 272518 117376 272524 117428
rect 272576 117416 272582 117428
rect 273530 117416 273536 117428
rect 272576 117388 273536 117416
rect 272576 117376 272582 117388
rect 273530 117376 273536 117388
rect 273588 117376 273594 117428
rect 284570 117376 284576 117428
rect 284628 117416 284634 117428
rect 285490 117416 285496 117428
rect 284628 117388 285496 117416
rect 284628 117376 284634 117388
rect 285490 117376 285496 117388
rect 285548 117376 285554 117428
rect 303430 117376 303436 117428
rect 303488 117416 303494 117428
rect 305638 117416 305644 117428
rect 303488 117388 305644 117416
rect 303488 117376 303494 117388
rect 305638 117376 305644 117388
rect 305696 117376 305702 117428
rect 237392 117320 238984 117348
rect 239398 117308 239404 117360
rect 239456 117348 239462 117360
rect 242250 117348 242256 117360
rect 239456 117320 242256 117348
rect 239456 117308 239462 117320
rect 242250 117308 242256 117320
rect 242308 117308 242314 117360
rect 242802 117308 242808 117360
rect 242860 117348 242866 117360
rect 249886 117348 249892 117360
rect 242860 117320 249892 117348
rect 242860 117308 242866 117320
rect 249886 117308 249892 117320
rect 249944 117308 249950 117360
rect 250438 117308 250444 117360
rect 250496 117348 250502 117360
rect 251450 117348 251456 117360
rect 250496 117320 251456 117348
rect 250496 117308 250502 117320
rect 251450 117308 251456 117320
rect 251508 117308 251514 117360
rect 252462 117308 252468 117360
rect 252520 117348 252526 117360
rect 259270 117348 259276 117360
rect 252520 117320 259276 117348
rect 252520 117308 252526 117320
rect 259270 117308 259276 117320
rect 259328 117308 259334 117360
rect 259362 117308 259368 117360
rect 259420 117348 259426 117360
rect 266814 117348 266820 117360
rect 259420 117320 266820 117348
rect 259420 117308 259426 117320
rect 266814 117308 266820 117320
rect 266872 117308 266878 117360
rect 271138 117308 271144 117360
rect 271196 117348 271202 117360
rect 272334 117348 272340 117360
rect 271196 117320 272340 117348
rect 271196 117308 271202 117320
rect 272334 117308 272340 117320
rect 272392 117308 272398 117360
rect 273162 117308 273168 117360
rect 273220 117348 273226 117360
rect 274174 117348 274180 117360
rect 273220 117320 274180 117348
rect 273220 117308 273226 117320
rect 274174 117308 274180 117320
rect 274232 117308 274238 117360
rect 279694 117308 279700 117360
rect 279752 117348 279758 117360
rect 280062 117348 280068 117360
rect 279752 117320 280068 117348
rect 279752 117308 279758 117320
rect 280062 117308 280068 117320
rect 280120 117308 280126 117360
rect 282086 117308 282092 117360
rect 282144 117348 282150 117360
rect 282822 117348 282828 117360
rect 282144 117320 282828 117348
rect 282144 117308 282150 117320
rect 282822 117308 282828 117320
rect 282880 117308 282886 117360
rect 283374 117308 283380 117360
rect 283432 117348 283438 117360
rect 284018 117348 284024 117360
rect 283432 117320 284024 117348
rect 283432 117308 283438 117320
rect 284018 117308 284024 117320
rect 284076 117308 284082 117360
rect 285214 117308 285220 117360
rect 285272 117348 285278 117360
rect 285582 117348 285588 117360
rect 285272 117320 285588 117348
rect 285272 117308 285278 117320
rect 285582 117308 285588 117320
rect 285640 117308 285646 117360
rect 286410 117308 286416 117360
rect 286468 117348 286474 117360
rect 286962 117348 286968 117360
rect 286468 117320 286968 117348
rect 286468 117308 286474 117320
rect 286962 117308 286968 117320
rect 287020 117308 287026 117360
rect 287606 117308 287612 117360
rect 287664 117348 287670 117360
rect 288342 117348 288348 117360
rect 287664 117320 288348 117348
rect 287664 117308 287670 117320
rect 288342 117308 288348 117320
rect 288400 117308 288406 117360
rect 288894 117308 288900 117360
rect 288952 117348 288958 117360
rect 289538 117348 289544 117360
rect 288952 117320 289544 117348
rect 288952 117308 288958 117320
rect 289538 117308 289544 117320
rect 289596 117308 289602 117360
rect 290090 117308 290096 117360
rect 290148 117348 290154 117360
rect 290734 117348 290740 117360
rect 290148 117320 290740 117348
rect 290148 117308 290154 117320
rect 290734 117308 290740 117320
rect 290792 117308 290798 117360
rect 291930 117308 291936 117360
rect 291988 117348 291994 117360
rect 292390 117348 292396 117360
rect 291988 117320 292396 117348
rect 291988 117308 291994 117320
rect 292390 117308 292396 117320
rect 292448 117308 292454 117360
rect 294322 117308 294328 117360
rect 294380 117348 294386 117360
rect 295242 117348 295248 117360
rect 294380 117320 295248 117348
rect 294380 117308 294386 117320
rect 295242 117308 295248 117320
rect 295300 117308 295306 117360
rect 295610 117308 295616 117360
rect 295668 117348 295674 117360
rect 296622 117348 296628 117360
rect 295668 117320 296628 117348
rect 295668 117308 295674 117320
rect 296622 117308 296628 117320
rect 296680 117308 296686 117360
rect 297450 117308 297456 117360
rect 297508 117348 297514 117360
rect 297910 117348 297916 117360
rect 297508 117320 297916 117348
rect 297508 117308 297514 117320
rect 297910 117308 297916 117320
rect 297968 117308 297974 117360
rect 299842 117308 299848 117360
rect 299900 117348 299906 117360
rect 300762 117348 300768 117360
rect 299900 117320 300768 117348
rect 299900 117308 299906 117320
rect 300762 117308 300768 117320
rect 300820 117308 300826 117360
rect 301682 117308 301688 117360
rect 301740 117348 301746 117360
rect 302878 117348 302884 117360
rect 301740 117320 302884 117348
rect 301740 117308 301746 117320
rect 302878 117308 302884 117320
rect 302936 117308 302942 117360
rect 302970 117308 302976 117360
rect 303028 117348 303034 117360
rect 303522 117348 303528 117360
rect 303028 117320 303528 117348
rect 303028 117308 303034 117320
rect 303522 117308 303528 117320
rect 303580 117308 303586 117360
rect 306650 117308 306656 117360
rect 306708 117348 306714 117360
rect 307662 117348 307668 117360
rect 306708 117320 307668 117348
rect 306708 117308 306714 117320
rect 307662 117308 307668 117320
rect 307720 117308 307726 117360
rect 307772 117348 307800 117456
rect 314102 117444 314108 117456
rect 314160 117444 314166 117496
rect 327442 117444 327448 117496
rect 327500 117484 327506 117496
rect 334618 117484 334624 117496
rect 327500 117456 334624 117484
rect 327500 117444 327506 117456
rect 334618 117444 334624 117456
rect 334676 117444 334682 117496
rect 336642 117444 336648 117496
rect 336700 117484 336706 117496
rect 341150 117484 341156 117496
rect 336700 117456 341156 117484
rect 336700 117444 336706 117456
rect 341150 117444 341156 117456
rect 341208 117444 341214 117496
rect 380250 117444 380256 117496
rect 380308 117484 380314 117496
rect 383654 117484 383660 117496
rect 380308 117456 383660 117484
rect 380308 117444 380314 117456
rect 383654 117444 383660 117456
rect 383712 117444 383718 117496
rect 413738 117444 413744 117496
rect 413796 117484 413802 117496
rect 414658 117484 414664 117496
rect 413796 117456 414664 117484
rect 413796 117444 413802 117456
rect 414658 117444 414664 117456
rect 414716 117444 414722 117496
rect 426342 117444 426348 117496
rect 426400 117484 426406 117496
rect 429838 117484 429844 117496
rect 426400 117456 429844 117484
rect 426400 117444 426406 117456
rect 429838 117444 429844 117456
rect 429896 117444 429902 117496
rect 310882 117376 310888 117428
rect 310940 117416 310946 117428
rect 315298 117416 315304 117428
rect 310940 117388 315304 117416
rect 310940 117376 310946 117388
rect 315298 117376 315304 117388
rect 315356 117376 315362 117428
rect 332962 117376 332968 117428
rect 333020 117416 333026 117428
rect 333882 117416 333888 117428
rect 333020 117388 333888 117416
rect 333020 117376 333026 117388
rect 333882 117376 333888 117388
rect 333940 117376 333946 117428
rect 334802 117376 334808 117428
rect 334860 117416 334866 117428
rect 338758 117416 338764 117428
rect 334860 117388 338764 117416
rect 334860 117376 334866 117388
rect 338758 117376 338764 117388
rect 338816 117376 338822 117428
rect 340322 117376 340328 117428
rect 340380 117416 340386 117428
rect 342898 117416 342904 117428
rect 340380 117388 342904 117416
rect 340380 117376 340386 117388
rect 342898 117376 342904 117388
rect 342956 117376 342962 117428
rect 344002 117376 344008 117428
rect 344060 117416 344066 117428
rect 345658 117416 345664 117428
rect 344060 117388 345664 117416
rect 344060 117376 344066 117388
rect 345658 117376 345664 117388
rect 345716 117376 345722 117428
rect 347590 117376 347596 117428
rect 347648 117416 347654 117428
rect 349798 117416 349804 117428
rect 347648 117388 349804 117416
rect 347648 117376 347654 117388
rect 349798 117376 349804 117388
rect 349856 117376 349862 117428
rect 367830 117376 367836 117428
rect 367888 117416 367894 117428
rect 369118 117416 369124 117428
rect 367888 117388 369124 117416
rect 367888 117376 367894 117388
rect 369118 117376 369124 117388
rect 369176 117376 369182 117428
rect 371510 117376 371516 117428
rect 371568 117416 371574 117428
rect 377398 117416 377404 117428
rect 371568 117388 377404 117416
rect 371568 117376 371574 117388
rect 377398 117376 377404 117388
rect 377456 117376 377462 117428
rect 399662 117376 399668 117428
rect 399720 117416 399726 117428
rect 400122 117416 400128 117428
rect 399720 117388 400128 117416
rect 399720 117376 399726 117388
rect 400122 117376 400128 117388
rect 400180 117376 400186 117428
rect 421742 117376 421748 117428
rect 421800 117416 421806 117428
rect 422202 117416 422208 117428
rect 421800 117388 422208 117416
rect 421800 117376 421806 117388
rect 422202 117376 422208 117388
rect 422260 117376 422266 117428
rect 312538 117348 312544 117360
rect 307772 117320 312544 117348
rect 312538 117308 312544 117320
rect 312596 117308 312602 117360
rect 313918 117308 313924 117360
rect 313976 117348 313982 117360
rect 314562 117348 314568 117360
rect 313976 117320 314568 117348
rect 313976 117308 313982 117320
rect 314562 117308 314568 117320
rect 314620 117308 314626 117360
rect 318242 117308 318248 117360
rect 318300 117348 318306 117360
rect 318702 117348 318708 117360
rect 318300 117320 318708 117348
rect 318300 117308 318306 117320
rect 318702 117308 318708 117320
rect 318760 117308 318766 117360
rect 319438 117308 319444 117360
rect 319496 117348 319502 117360
rect 320082 117348 320088 117360
rect 319496 117320 320088 117348
rect 319496 117308 319502 117320
rect 320082 117308 320088 117320
rect 320140 117308 320146 117360
rect 322566 117308 322572 117360
rect 322624 117348 322630 117360
rect 322842 117348 322848 117360
rect 322624 117320 322848 117348
rect 322624 117308 322630 117320
rect 322842 117308 322848 117320
rect 322900 117308 322906 117360
rect 323762 117308 323768 117360
rect 323820 117348 323826 117360
rect 324222 117348 324228 117360
rect 323820 117320 324228 117348
rect 323820 117308 323826 117320
rect 324222 117308 324228 117320
rect 324280 117308 324286 117360
rect 324958 117308 324964 117360
rect 325016 117348 325022 117360
rect 325510 117348 325516 117360
rect 325016 117320 325516 117348
rect 325016 117308 325022 117320
rect 325510 117308 325516 117320
rect 325568 117308 325574 117360
rect 326246 117308 326252 117360
rect 326304 117348 326310 117360
rect 326982 117348 326988 117360
rect 326304 117320 326988 117348
rect 326304 117308 326310 117320
rect 326982 117308 326988 117320
rect 327040 117308 327046 117360
rect 328086 117308 328092 117360
rect 328144 117348 328150 117360
rect 328362 117348 328368 117360
rect 328144 117320 328368 117348
rect 328144 117308 328150 117320
rect 328362 117308 328368 117320
rect 328420 117308 328426 117360
rect 329282 117308 329288 117360
rect 329340 117348 329346 117360
rect 329742 117348 329748 117360
rect 329340 117320 329748 117348
rect 329340 117308 329346 117320
rect 329742 117308 329748 117320
rect 329800 117308 329806 117360
rect 330478 117308 330484 117360
rect 330536 117348 330542 117360
rect 331122 117348 331128 117360
rect 330536 117320 331128 117348
rect 330536 117308 330542 117320
rect 331122 117308 331128 117320
rect 331180 117308 331186 117360
rect 331674 117308 331680 117360
rect 331732 117348 331738 117360
rect 332502 117348 332508 117360
rect 331732 117320 332508 117348
rect 331732 117308 331738 117320
rect 332502 117308 332508 117320
rect 332560 117308 332566 117360
rect 333514 117308 333520 117360
rect 333572 117348 333578 117360
rect 333790 117348 333796 117360
rect 333572 117320 333796 117348
rect 333572 117308 333578 117320
rect 333790 117308 333796 117320
rect 333848 117308 333854 117360
rect 337194 117308 337200 117360
rect 337252 117348 337258 117360
rect 338022 117348 338028 117360
rect 337252 117320 338028 117348
rect 337252 117308 337258 117320
rect 338022 117308 338028 117320
rect 338080 117308 338086 117360
rect 341518 117308 341524 117360
rect 341576 117348 341582 117360
rect 342162 117348 342168 117360
rect 341576 117320 342168 117348
rect 341576 117308 341582 117320
rect 342162 117308 342168 117320
rect 342220 117308 342226 117360
rect 342714 117308 342720 117360
rect 342772 117348 342778 117360
rect 343542 117348 343548 117360
rect 342772 117320 343548 117348
rect 342772 117308 342778 117320
rect 343542 117308 343548 117320
rect 343600 117308 343606 117360
rect 344554 117308 344560 117360
rect 344612 117348 344618 117360
rect 344922 117348 344928 117360
rect 344612 117320 344928 117348
rect 344612 117308 344618 117320
rect 344922 117308 344928 117320
rect 344980 117308 344986 117360
rect 347038 117308 347044 117360
rect 347096 117348 347102 117360
rect 347682 117348 347688 117360
rect 347096 117320 347688 117348
rect 347096 117308 347102 117320
rect 347682 117308 347688 117320
rect 347740 117308 347746 117360
rect 348234 117308 348240 117360
rect 348292 117348 348298 117360
rect 349062 117348 349068 117360
rect 348292 117320 349068 117348
rect 348292 117308 348298 117320
rect 349062 117308 349068 117320
rect 349120 117308 349126 117360
rect 350074 117308 350080 117360
rect 350132 117348 350138 117360
rect 350442 117348 350448 117360
rect 350132 117320 350448 117348
rect 350132 117308 350138 117320
rect 350442 117308 350448 117320
rect 350500 117308 350506 117360
rect 351270 117308 351276 117360
rect 351328 117348 351334 117360
rect 352466 117348 352472 117360
rect 351328 117320 352472 117348
rect 351328 117308 351334 117320
rect 352466 117308 352472 117320
rect 352524 117308 352530 117360
rect 352558 117308 352564 117360
rect 352616 117348 352622 117360
rect 353202 117348 353208 117360
rect 352616 117320 353208 117348
rect 352616 117308 352622 117320
rect 353202 117308 353208 117320
rect 353260 117308 353266 117360
rect 353754 117308 353760 117360
rect 353812 117348 353818 117360
rect 354582 117348 354588 117360
rect 353812 117320 354588 117348
rect 353812 117308 353818 117320
rect 354582 117308 354588 117320
rect 354640 117308 354646 117360
rect 355594 117308 355600 117360
rect 355652 117348 355658 117360
rect 355962 117348 355968 117360
rect 355652 117320 355968 117348
rect 355652 117308 355658 117320
rect 355962 117308 355968 117320
rect 356020 117308 356026 117360
rect 358078 117308 358084 117360
rect 358136 117348 358142 117360
rect 358630 117348 358636 117360
rect 358136 117320 358636 117348
rect 358136 117308 358142 117320
rect 358630 117308 358636 117320
rect 358688 117308 358694 117360
rect 361114 117308 361120 117360
rect 361172 117348 361178 117360
rect 361482 117348 361488 117360
rect 361172 117320 361488 117348
rect 361172 117308 361178 117320
rect 361482 117308 361488 117320
rect 361540 117308 361546 117360
rect 363598 117308 363604 117360
rect 363656 117348 363662 117360
rect 364242 117348 364248 117360
rect 363656 117320 364248 117348
rect 363656 117308 363662 117320
rect 364242 117308 364248 117320
rect 364300 117308 364306 117360
rect 364794 117308 364800 117360
rect 364852 117348 364858 117360
rect 365622 117348 365628 117360
rect 364852 117320 365628 117348
rect 364852 117308 364858 117320
rect 365622 117308 365628 117320
rect 365680 117308 365686 117360
rect 366634 117308 366640 117360
rect 366692 117348 366698 117360
rect 367002 117348 367008 117360
rect 366692 117320 367008 117348
rect 366692 117308 366698 117320
rect 367002 117308 367008 117320
rect 367060 117308 367066 117360
rect 369026 117308 369032 117360
rect 369084 117348 369090 117360
rect 369762 117348 369768 117360
rect 369084 117320 369768 117348
rect 369084 117308 369090 117320
rect 369762 117308 369768 117320
rect 369820 117308 369826 117360
rect 370314 117308 370320 117360
rect 370372 117348 370378 117360
rect 371142 117348 371148 117360
rect 370372 117320 371148 117348
rect 370372 117308 370378 117320
rect 371142 117308 371148 117320
rect 371200 117308 371206 117360
rect 372154 117308 372160 117360
rect 372212 117348 372218 117360
rect 372522 117348 372528 117360
rect 372212 117320 372528 117348
rect 372212 117308 372218 117320
rect 372522 117308 372528 117320
rect 372580 117308 372586 117360
rect 374546 117308 374552 117360
rect 374604 117348 374610 117360
rect 375190 117348 375196 117360
rect 374604 117320 375196 117348
rect 374604 117308 374610 117320
rect 375190 117308 375196 117320
rect 375248 117308 375254 117360
rect 375834 117308 375840 117360
rect 375892 117348 375898 117360
rect 376662 117348 376668 117360
rect 375892 117320 376668 117348
rect 375892 117308 375898 117320
rect 376662 117308 376668 117320
rect 376720 117308 376726 117360
rect 377674 117308 377680 117360
rect 377732 117348 377738 117360
rect 378042 117348 378048 117360
rect 377732 117320 378048 117348
rect 377732 117308 377738 117320
rect 378042 117308 378048 117320
rect 378100 117308 378106 117360
rect 378870 117308 378876 117360
rect 378928 117348 378934 117360
rect 379422 117348 379428 117360
rect 378928 117320 379428 117348
rect 378928 117308 378934 117320
rect 379422 117308 379428 117320
rect 379480 117308 379486 117360
rect 380066 117308 380072 117360
rect 380124 117348 380130 117360
rect 380802 117348 380808 117360
rect 380124 117320 380808 117348
rect 380124 117308 380130 117320
rect 380802 117308 380808 117320
rect 380860 117308 380866 117360
rect 381354 117308 381360 117360
rect 381412 117348 381418 117360
rect 382182 117348 382188 117360
rect 381412 117320 382188 117348
rect 381412 117308 381418 117320
rect 382182 117308 382188 117320
rect 382240 117308 382246 117360
rect 382550 117308 382556 117360
rect 382608 117348 382614 117360
rect 383562 117348 383568 117360
rect 382608 117320 383568 117348
rect 382608 117308 382614 117320
rect 383562 117308 383568 117320
rect 383620 117308 383626 117360
rect 384390 117308 384396 117360
rect 384448 117348 384454 117360
rect 384850 117348 384856 117360
rect 384448 117320 384856 117348
rect 384448 117308 384454 117320
rect 384850 117308 384856 117320
rect 384908 117308 384914 117360
rect 385586 117308 385592 117360
rect 385644 117348 385650 117360
rect 386322 117348 386328 117360
rect 385644 117320 386328 117348
rect 385644 117308 385650 117320
rect 386322 117308 386328 117320
rect 386380 117308 386386 117360
rect 386782 117308 386788 117360
rect 386840 117348 386846 117360
rect 387610 117348 387616 117360
rect 386840 117320 387616 117348
rect 386840 117308 386846 117320
rect 387610 117308 387616 117320
rect 387668 117308 387674 117360
rect 388070 117308 388076 117360
rect 388128 117348 388134 117360
rect 388898 117348 388904 117360
rect 388128 117320 388904 117348
rect 388128 117308 388134 117320
rect 388898 117308 388904 117320
rect 388956 117308 388962 117360
rect 389910 117308 389916 117360
rect 389968 117348 389974 117360
rect 390370 117348 390376 117360
rect 389968 117320 390376 117348
rect 389968 117308 389974 117320
rect 390370 117308 390376 117320
rect 390428 117308 390434 117360
rect 391106 117308 391112 117360
rect 391164 117348 391170 117360
rect 391842 117348 391848 117360
rect 391164 117320 391848 117348
rect 391164 117308 391170 117320
rect 391842 117308 391848 117320
rect 391900 117308 391906 117360
rect 392302 117308 392308 117360
rect 392360 117348 392366 117360
rect 393130 117348 393136 117360
rect 392360 117320 393136 117348
rect 392360 117308 392366 117320
rect 393130 117308 393136 117320
rect 393188 117308 393194 117360
rect 393590 117308 393596 117360
rect 393648 117348 393654 117360
rect 394418 117348 394424 117360
rect 393648 117320 394424 117348
rect 393648 117308 393654 117320
rect 394418 117308 394424 117320
rect 394476 117308 394482 117360
rect 395430 117308 395436 117360
rect 395488 117348 395494 117360
rect 395890 117348 395896 117360
rect 395488 117320 395896 117348
rect 395488 117308 395494 117320
rect 395890 117308 395896 117320
rect 395948 117308 395954 117360
rect 396626 117308 396632 117360
rect 396684 117348 396690 117360
rect 397362 117348 397368 117360
rect 396684 117320 397368 117348
rect 396684 117308 396690 117320
rect 397362 117308 397368 117320
rect 397420 117308 397426 117360
rect 397822 117308 397828 117360
rect 397880 117348 397886 117360
rect 398650 117348 398656 117360
rect 397880 117320 398656 117348
rect 397880 117308 397886 117320
rect 398650 117308 398656 117320
rect 398708 117308 398714 117360
rect 399110 117308 399116 117360
rect 399168 117348 399174 117360
rect 399938 117348 399944 117360
rect 399168 117320 399944 117348
rect 399168 117308 399174 117320
rect 399938 117308 399944 117320
rect 399996 117308 400002 117360
rect 402146 117308 402152 117360
rect 402204 117348 402210 117360
rect 402790 117348 402796 117360
rect 402204 117320 402796 117348
rect 402204 117308 402210 117320
rect 402790 117308 402796 117320
rect 402848 117308 402854 117360
rect 403342 117308 403348 117360
rect 403400 117348 403406 117360
rect 404262 117348 404268 117360
rect 403400 117320 404268 117348
rect 403400 117308 403406 117320
rect 404262 117308 404268 117320
rect 404320 117308 404326 117360
rect 405182 117308 405188 117360
rect 405240 117348 405246 117360
rect 405642 117348 405648 117360
rect 405240 117320 405648 117348
rect 405240 117308 405246 117320
rect 405642 117308 405648 117320
rect 405700 117308 405706 117360
rect 406378 117308 406384 117360
rect 406436 117348 406442 117360
rect 407022 117348 407028 117360
rect 406436 117320 407028 117348
rect 406436 117308 406442 117320
rect 407022 117308 407028 117320
rect 407080 117308 407086 117360
rect 407666 117308 407672 117360
rect 407724 117348 407730 117360
rect 408402 117348 408408 117360
rect 407724 117320 408408 117348
rect 407724 117308 407730 117320
rect 408402 117308 408408 117320
rect 408460 117308 408466 117360
rect 408862 117308 408868 117360
rect 408920 117348 408926 117360
rect 409690 117348 409696 117360
rect 408920 117320 409696 117348
rect 408920 117308 408926 117320
rect 409690 117308 409696 117320
rect 409748 117308 409754 117360
rect 410702 117308 410708 117360
rect 410760 117348 410766 117360
rect 411162 117348 411168 117360
rect 410760 117320 411168 117348
rect 410760 117308 410766 117320
rect 411162 117308 411168 117320
rect 411220 117308 411226 117360
rect 413186 117308 413192 117360
rect 413244 117348 413250 117360
rect 413922 117348 413928 117360
rect 413244 117320 413928 117348
rect 413244 117308 413250 117320
rect 413922 117308 413928 117320
rect 413980 117308 413986 117360
rect 414382 117308 414388 117360
rect 414440 117348 414446 117360
rect 415302 117348 415308 117360
rect 414440 117320 415308 117348
rect 414440 117308 414446 117320
rect 415302 117308 415308 117320
rect 415360 117308 415366 117360
rect 416222 117308 416228 117360
rect 416280 117348 416286 117360
rect 416682 117348 416688 117360
rect 416280 117320 416688 117348
rect 416280 117308 416286 117320
rect 416682 117308 416688 117320
rect 416740 117308 416746 117360
rect 418614 117308 418620 117360
rect 418672 117348 418678 117360
rect 419442 117348 419448 117360
rect 418672 117320 419448 117348
rect 418672 117308 418678 117320
rect 419442 117308 419448 117320
rect 419500 117308 419506 117360
rect 419902 117308 419908 117360
rect 419960 117348 419966 117360
rect 420822 117348 420828 117360
rect 419960 117320 420828 117348
rect 419960 117308 419966 117320
rect 420822 117308 420828 117320
rect 420880 117308 420886 117360
rect 422938 117308 422944 117360
rect 422996 117348 423002 117360
rect 423582 117348 423588 117360
rect 422996 117320 423588 117348
rect 422996 117308 423002 117320
rect 423582 117308 423588 117320
rect 423640 117308 423646 117360
rect 424134 117308 424140 117360
rect 424192 117348 424198 117360
rect 424962 117348 424968 117360
rect 424192 117320 424968 117348
rect 424192 117308 424198 117320
rect 424962 117308 424968 117320
rect 425020 117308 425026 117360
rect 425422 117308 425428 117360
rect 425480 117348 425486 117360
rect 426342 117348 426348 117360
rect 425480 117320 426348 117348
rect 425480 117308 425486 117320
rect 426342 117308 426348 117320
rect 426400 117308 426406 117360
rect 427262 117308 427268 117360
rect 427320 117348 427326 117360
rect 427722 117348 427728 117360
rect 427320 117320 427728 117348
rect 427320 117308 427326 117320
rect 427722 117308 427728 117320
rect 427780 117308 427786 117360
rect 429654 117308 429660 117360
rect 429712 117348 429718 117360
rect 430482 117348 430488 117360
rect 429712 117320 430488 117348
rect 429712 117308 429718 117320
rect 430482 117308 430488 117320
rect 430540 117308 430546 117360
rect 430942 117308 430948 117360
rect 431000 117348 431006 117360
rect 431862 117348 431868 117360
rect 431000 117320 431868 117348
rect 431000 117308 431006 117320
rect 431862 117308 431868 117320
rect 431920 117308 431926 117360
rect 432782 117308 432788 117360
rect 432840 117348 432846 117360
rect 433242 117348 433248 117360
rect 432840 117320 433248 117348
rect 432840 117308 432846 117320
rect 433242 117308 433248 117320
rect 433300 117308 433306 117360
rect 433978 117308 433984 117360
rect 434036 117348 434042 117360
rect 439498 117348 439504 117360
rect 434036 117320 439504 117348
rect 434036 117308 434042 117320
rect 439498 117308 439504 117320
rect 439556 117308 439562 117360
rect 133782 117240 133788 117292
rect 133840 117280 133846 117292
rect 190564 117280 190592 117308
rect 133840 117252 190592 117280
rect 133840 117240 133846 117252
rect 130286 117172 130292 117224
rect 130344 117212 130350 117224
rect 133874 117212 133880 117224
rect 130344 117184 133880 117212
rect 130344 117172 130350 117184
rect 133874 117172 133880 117184
rect 133932 117172 133938 117224
rect 143442 117172 143448 117224
rect 143500 117212 143506 117224
rect 154482 117212 154488 117224
rect 143500 117184 154488 117212
rect 143500 117172 143506 117184
rect 154482 117172 154488 117184
rect 154540 117172 154546 117224
rect 171134 117212 171140 117224
rect 162780 117184 171140 117212
rect 133874 117036 133880 117088
rect 133932 117076 133938 117088
rect 143442 117076 143448 117088
rect 133932 117048 143448 117076
rect 133932 117036 133938 117048
rect 143442 117036 143448 117048
rect 143500 117036 143506 117088
rect 161382 117036 161388 117088
rect 161440 117076 161446 117088
rect 162780 117076 162808 117184
rect 171134 117172 171140 117184
rect 171192 117172 171198 117224
rect 182174 117212 182180 117224
rect 182100 117184 182180 117212
rect 161440 117048 162808 117076
rect 161440 117036 161446 117048
rect 180702 117036 180708 117088
rect 180760 117076 180766 117088
rect 182100 117076 182128 117184
rect 182174 117172 182180 117184
rect 182232 117172 182238 117224
rect 404354 117172 404360 117224
rect 404412 117212 404418 117224
rect 410518 117212 410524 117224
rect 404412 117184 410524 117212
rect 404412 117172 404418 117184
rect 410518 117172 410524 117184
rect 410576 117172 410582 117224
rect 180760 117048 182128 117076
rect 180760 117036 180766 117048
rect 154482 116900 154488 116952
rect 154540 116940 154546 116952
rect 161382 116940 161388 116952
rect 154540 116912 161388 116940
rect 154540 116900 154546 116912
rect 161382 116900 161388 116912
rect 161440 116900 161446 116952
rect 208486 116628 208492 116680
rect 208544 116668 208550 116680
rect 209222 116668 209228 116680
rect 208544 116640 209228 116668
rect 208544 116628 208550 116640
rect 209222 116628 209228 116640
rect 209280 116628 209286 116680
rect 205634 116560 205640 116612
rect 205692 116600 205698 116612
rect 206186 116600 206192 116612
rect 205692 116572 206192 116600
rect 205692 116560 205698 116572
rect 206186 116560 206192 116572
rect 206244 116560 206250 116612
rect 208394 116560 208400 116612
rect 208452 116600 208458 116612
rect 208670 116600 208676 116612
rect 208452 116572 208676 116600
rect 208452 116560 208458 116572
rect 208670 116560 208676 116572
rect 208728 116560 208734 116612
rect 212534 116560 212540 116612
rect 212592 116600 212598 116612
rect 212902 116600 212908 116612
rect 212592 116572 212908 116600
rect 212592 116560 212598 116572
rect 212902 116560 212908 116572
rect 212960 116560 212966 116612
rect 214006 116560 214012 116612
rect 214064 116600 214070 116612
rect 214742 116600 214748 116612
rect 214064 116572 214748 116600
rect 214064 116560 214070 116572
rect 214742 116560 214748 116572
rect 214800 116560 214806 116612
rect 420270 115948 420276 116000
rect 420328 115988 420334 116000
rect 420454 115988 420460 116000
rect 420328 115960 420460 115988
rect 420328 115948 420334 115960
rect 420454 115948 420460 115960
rect 420512 115948 420518 116000
rect 128722 115880 128728 115932
rect 128780 115920 128786 115932
rect 128998 115920 129004 115932
rect 128780 115892 129004 115920
rect 128780 115880 128786 115892
rect 128998 115880 129004 115892
rect 129056 115880 129062 115932
rect 143626 115880 143632 115932
rect 143684 115920 143690 115932
rect 143718 115920 143724 115932
rect 143684 115892 143724 115920
rect 143684 115880 143690 115892
rect 143718 115880 143724 115892
rect 143776 115880 143782 115932
rect 144914 115880 144920 115932
rect 144972 115920 144978 115932
rect 145282 115920 145288 115932
rect 144972 115892 145288 115920
rect 144972 115880 144978 115892
rect 145282 115880 145288 115892
rect 145340 115880 145346 115932
rect 168466 115880 168472 115932
rect 168524 115920 168530 115932
rect 168558 115920 168564 115932
rect 168524 115892 168564 115920
rect 168524 115880 168530 115892
rect 168558 115880 168564 115892
rect 168616 115880 168622 115932
rect 238938 115880 238944 115932
rect 238996 115920 239002 115932
rect 239122 115920 239128 115932
rect 238996 115892 239128 115920
rect 238996 115880 239002 115892
rect 239122 115880 239128 115892
rect 239180 115880 239186 115932
rect 248230 115880 248236 115932
rect 248288 115920 248294 115932
rect 248322 115920 248328 115932
rect 248288 115892 248328 115920
rect 248288 115880 248294 115892
rect 248322 115880 248328 115892
rect 248380 115880 248386 115932
rect 253750 115880 253756 115932
rect 253808 115920 253814 115932
rect 253934 115920 253940 115932
rect 253808 115892 253940 115920
rect 253808 115880 253814 115892
rect 253934 115880 253940 115892
rect 253992 115880 253998 115932
rect 314010 115880 314016 115932
rect 314068 115920 314074 115932
rect 314102 115920 314108 115932
rect 314068 115892 314108 115920
rect 314068 115880 314074 115892
rect 314102 115880 314108 115892
rect 314160 115880 314166 115932
rect 339678 115880 339684 115932
rect 339736 115920 339742 115932
rect 339862 115920 339868 115932
rect 339736 115892 339868 115920
rect 339736 115880 339742 115892
rect 339862 115880 339868 115892
rect 339920 115880 339926 115932
rect 341242 115880 341248 115932
rect 341300 115920 341306 115932
rect 341426 115920 341432 115932
rect 341300 115892 341432 115920
rect 341300 115880 341306 115892
rect 341426 115880 341432 115892
rect 341484 115880 341490 115932
rect 343910 115880 343916 115932
rect 343968 115920 343974 115932
rect 344094 115920 344100 115932
rect 343968 115892 344100 115920
rect 343968 115880 343974 115892
rect 344094 115880 344100 115892
rect 344152 115880 344158 115932
rect 409322 114588 409328 114640
rect 409380 114628 409386 114640
rect 409598 114628 409604 114640
rect 409380 114600 409604 114628
rect 409380 114588 409386 114600
rect 409598 114588 409604 114600
rect 409656 114588 409662 114640
rect 147950 114520 147956 114572
rect 148008 114560 148014 114572
rect 148594 114560 148600 114572
rect 148008 114532 148600 114560
rect 148008 114520 148014 114532
rect 148594 114520 148600 114532
rect 148652 114520 148658 114572
rect 157426 114520 157432 114572
rect 157484 114560 157490 114572
rect 157794 114560 157800 114572
rect 157484 114532 157800 114560
rect 157484 114520 157490 114532
rect 157794 114520 157800 114532
rect 157852 114520 157858 114572
rect 179598 114520 179604 114572
rect 179656 114560 179662 114572
rect 179966 114560 179972 114572
rect 179656 114532 179972 114560
rect 179656 114520 179662 114532
rect 179966 114520 179972 114532
rect 180024 114520 180030 114572
rect 245378 114520 245384 114572
rect 245436 114560 245442 114572
rect 245746 114560 245752 114572
rect 245436 114532 245752 114560
rect 245436 114520 245442 114532
rect 245746 114520 245752 114532
rect 245804 114520 245810 114572
rect 250070 114520 250076 114572
rect 250128 114560 250134 114572
rect 250346 114560 250352 114572
rect 250128 114532 250352 114560
rect 250128 114520 250134 114532
rect 250346 114520 250352 114532
rect 250404 114520 250410 114572
rect 276106 114520 276112 114572
rect 276164 114560 276170 114572
rect 276198 114560 276204 114572
rect 276164 114532 276204 114560
rect 276164 114520 276170 114532
rect 276198 114520 276204 114532
rect 276256 114520 276262 114572
rect 382918 114520 382924 114572
rect 382976 114560 382982 114572
rect 383102 114560 383108 114572
rect 382976 114532 383108 114560
rect 382976 114520 382982 114532
rect 383102 114520 383108 114532
rect 383160 114520 383166 114572
rect 403710 114520 403716 114572
rect 403768 114560 403774 114572
rect 403894 114560 403900 114572
rect 403768 114532 403900 114560
rect 403768 114520 403774 114532
rect 403894 114520 403900 114532
rect 403952 114520 403958 114572
rect 161658 114452 161664 114504
rect 161716 114492 161722 114504
rect 161842 114492 161848 114504
rect 161716 114464 161848 114492
rect 161716 114452 161722 114464
rect 161842 114452 161848 114464
rect 161900 114452 161906 114504
rect 185026 114452 185032 114504
rect 185084 114492 185090 114504
rect 185118 114492 185124 114504
rect 185084 114464 185124 114492
rect 185084 114452 185090 114464
rect 185118 114452 185124 114464
rect 185176 114452 185182 114504
rect 189074 114452 189080 114504
rect 189132 114492 189138 114504
rect 189258 114492 189264 114504
rect 189132 114464 189264 114492
rect 189132 114452 189138 114464
rect 189258 114452 189264 114464
rect 189316 114452 189322 114504
rect 409414 114452 409420 114504
rect 409472 114492 409478 114504
rect 409598 114492 409604 114504
rect 409472 114464 409604 114492
rect 409472 114452 409478 114464
rect 409598 114452 409604 114464
rect 409656 114452 409662 114504
rect 425974 114452 425980 114504
rect 426032 114452 426038 114504
rect 431586 114452 431592 114504
rect 431644 114492 431650 114504
rect 431678 114492 431684 114504
rect 431644 114464 431684 114492
rect 431644 114452 431650 114464
rect 431678 114452 431684 114464
rect 431736 114452 431742 114504
rect 147950 114384 147956 114436
rect 148008 114424 148014 114436
rect 148226 114424 148232 114436
rect 148008 114396 148232 114424
rect 148008 114384 148014 114396
rect 148226 114384 148232 114396
rect 148284 114384 148290 114436
rect 425992 114424 426020 114452
rect 426158 114424 426164 114436
rect 425992 114396 426164 114424
rect 426158 114384 426164 114396
rect 426216 114384 426222 114436
rect 133874 113840 133880 113892
rect 133932 113880 133938 113892
rect 134518 113880 134524 113892
rect 133932 113852 134524 113880
rect 133932 113840 133938 113852
rect 134518 113840 134524 113852
rect 134576 113840 134582 113892
rect 135254 113840 135260 113892
rect 135312 113880 135318 113892
rect 135714 113880 135720 113892
rect 135312 113852 135720 113880
rect 135312 113840 135318 113852
rect 135714 113840 135720 113852
rect 135772 113840 135778 113892
rect 136726 113840 136732 113892
rect 136784 113880 136790 113892
rect 137002 113880 137008 113892
rect 136784 113852 137008 113880
rect 136784 113840 136790 113852
rect 137002 113840 137008 113852
rect 137060 113840 137066 113892
rect 139486 113840 139492 113892
rect 139544 113880 139550 113892
rect 140038 113880 140044 113892
rect 139544 113852 140044 113880
rect 139544 113840 139550 113852
rect 140038 113840 140044 113852
rect 140096 113840 140102 113892
rect 166994 113840 167000 113892
rect 167052 113880 167058 113892
rect 167638 113880 167644 113892
rect 167052 113852 167644 113880
rect 167052 113840 167058 113852
rect 167638 113840 167644 113852
rect 167696 113840 167702 113892
rect 169846 113840 169852 113892
rect 169904 113880 169910 113892
rect 170674 113880 170680 113892
rect 169904 113852 170680 113880
rect 169904 113840 169910 113852
rect 170674 113840 170680 113852
rect 170732 113840 170738 113892
rect 178034 113840 178040 113892
rect 178092 113880 178098 113892
rect 178586 113880 178592 113892
rect 178092 113852 178592 113880
rect 178092 113840 178098 113852
rect 178586 113840 178592 113852
rect 178644 113840 178650 113892
rect 186314 113840 186320 113892
rect 186372 113880 186378 113892
rect 187142 113880 187148 113892
rect 186372 113852 187148 113880
rect 186372 113840 186378 113852
rect 187142 113840 187148 113852
rect 187200 113840 187206 113892
rect 194594 113840 194600 113892
rect 194652 113880 194658 113892
rect 195146 113880 195152 113892
rect 194652 113852 195152 113880
rect 194652 113840 194658 113852
rect 195146 113840 195152 113852
rect 195204 113840 195210 113892
rect 201494 113840 201500 113892
rect 201552 113880 201558 113892
rect 201862 113880 201868 113892
rect 201552 113852 201868 113880
rect 201552 113840 201558 113852
rect 201862 113840 201868 113852
rect 201920 113840 201926 113892
rect 136634 113772 136640 113824
rect 136692 113812 136698 113824
rect 137554 113812 137560 113824
rect 136692 113784 137560 113812
rect 136692 113772 136698 113784
rect 137554 113772 137560 113784
rect 137612 113772 137618 113824
rect 222194 113704 222200 113756
rect 222252 113744 222258 113756
rect 222654 113744 222660 113756
rect 222252 113716 222660 113744
rect 222252 113704 222258 113716
rect 222654 113704 222660 113716
rect 222712 113704 222718 113756
rect 233418 113160 233424 113212
rect 233476 113200 233482 113212
rect 233694 113200 233700 113212
rect 233476 113172 233700 113200
rect 233476 113160 233482 113172
rect 233694 113160 233700 113172
rect 233752 113160 233758 113212
rect 414750 113160 414756 113212
rect 414808 113200 414814 113212
rect 415210 113200 415216 113212
rect 414808 113172 415216 113200
rect 414808 113160 414814 113172
rect 415210 113160 415216 113172
rect 415268 113160 415274 113212
rect 175366 111732 175372 111784
rect 175424 111772 175430 111784
rect 176194 111772 176200 111784
rect 175424 111744 176200 111772
rect 175424 111732 175430 111744
rect 176194 111732 176200 111744
rect 176252 111732 176258 111784
rect 436922 111732 436928 111784
rect 436980 111772 436986 111784
rect 579798 111772 579804 111784
rect 436980 111744 579804 111772
rect 436980 111732 436986 111744
rect 579798 111732 579804 111744
rect 579856 111732 579862 111784
rect 200114 111460 200120 111512
rect 200172 111500 200178 111512
rect 200666 111500 200672 111512
rect 200172 111472 200672 111500
rect 200172 111460 200178 111472
rect 200666 111460 200672 111472
rect 200724 111460 200730 111512
rect 198734 110576 198740 110628
rect 198792 110616 198798 110628
rect 199470 110616 199476 110628
rect 198792 110588 199476 110616
rect 198792 110576 198798 110588
rect 199470 110576 199476 110588
rect 199528 110576 199534 110628
rect 245746 109964 245752 110016
rect 245804 110004 245810 110016
rect 246574 110004 246580 110016
rect 245804 109976 246580 110004
rect 245804 109964 245810 109976
rect 246574 109964 246580 109976
rect 246632 109964 246638 110016
rect 153286 109760 153292 109812
rect 153344 109800 153350 109812
rect 154114 109800 154120 109812
rect 153344 109772 154120 109800
rect 153344 109760 153350 109772
rect 154114 109760 154120 109772
rect 154172 109760 154178 109812
rect 172514 109080 172520 109132
rect 172572 109120 172578 109132
rect 173066 109120 173072 109132
rect 172572 109092 173072 109120
rect 172572 109080 172578 109092
rect 173066 109080 173072 109092
rect 173124 109080 173130 109132
rect 179598 109080 179604 109132
rect 179656 109080 179662 109132
rect 190730 109120 190736 109132
rect 190656 109092 190736 109120
rect 159082 109052 159088 109064
rect 159008 109024 159088 109052
rect 159008 108996 159036 109024
rect 159082 109012 159088 109024
rect 159140 109012 159146 109064
rect 168558 109052 168564 109064
rect 168484 109024 168564 109052
rect 168484 108996 168512 109024
rect 168558 109012 168564 109024
rect 168616 109012 168622 109064
rect 179616 108996 179644 109080
rect 190656 108996 190684 109092
rect 190730 109080 190736 109092
rect 190788 109080 190794 109132
rect 196066 109080 196072 109132
rect 196124 109080 196130 109132
rect 383102 109080 383108 109132
rect 383160 109080 383166 109132
rect 196084 108996 196112 109080
rect 314102 109052 314108 109064
rect 314028 109024 314108 109052
rect 314028 108996 314056 109024
rect 314102 109012 314108 109024
rect 314160 109012 314166 109064
rect 383120 108996 383148 109080
rect 388806 109012 388812 109064
rect 388864 109052 388870 109064
rect 388990 109052 388996 109064
rect 388864 109024 388996 109052
rect 388864 109012 388870 109024
rect 388990 109012 388996 109024
rect 389048 109012 389054 109064
rect 394326 109012 394332 109064
rect 394384 109052 394390 109064
rect 394510 109052 394516 109064
rect 394384 109024 394516 109052
rect 394384 109012 394390 109024
rect 394510 109012 394516 109024
rect 394568 109012 394574 109064
rect 403894 109012 403900 109064
rect 403952 109052 403958 109064
rect 403952 109024 404032 109052
rect 403952 109012 403958 109024
rect 404004 108996 404032 109024
rect 3234 108944 3240 108996
rect 3292 108984 3298 108996
rect 131206 108984 131212 108996
rect 3292 108956 131212 108984
rect 3292 108944 3298 108956
rect 131206 108944 131212 108956
rect 131264 108944 131270 108996
rect 158990 108944 158996 108996
rect 159048 108944 159054 108996
rect 168466 108944 168472 108996
rect 168524 108944 168530 108996
rect 179598 108944 179604 108996
rect 179656 108944 179662 108996
rect 190638 108944 190644 108996
rect 190696 108944 190702 108996
rect 196066 108944 196072 108996
rect 196124 108944 196130 108996
rect 314010 108944 314016 108996
rect 314068 108944 314074 108996
rect 383102 108944 383108 108996
rect 383160 108944 383166 108996
rect 403986 108944 403992 108996
rect 404044 108944 404050 108996
rect 217042 106468 217048 106480
rect 216968 106440 217048 106468
rect 216968 106344 216996 106440
rect 217042 106428 217048 106440
rect 217100 106428 217106 106480
rect 317046 106360 317052 106412
rect 317104 106400 317110 106412
rect 317230 106400 317236 106412
rect 317104 106372 317236 106400
rect 317104 106360 317110 106372
rect 317230 106360 317236 106372
rect 317288 106360 317294 106412
rect 143626 106292 143632 106344
rect 143684 106332 143690 106344
rect 143718 106332 143724 106344
rect 143684 106304 143724 106332
rect 143684 106292 143690 106304
rect 143718 106292 143724 106304
rect 143776 106292 143782 106344
rect 216950 106292 216956 106344
rect 217008 106292 217014 106344
rect 245378 106292 245384 106344
rect 245436 106332 245442 106344
rect 245470 106332 245476 106344
rect 245436 106304 245476 106332
rect 245436 106292 245442 106304
rect 245470 106292 245476 106304
rect 245528 106292 245534 106344
rect 248230 106292 248236 106344
rect 248288 106332 248294 106344
rect 248322 106332 248328 106344
rect 248288 106304 248328 106332
rect 248288 106292 248294 106304
rect 248322 106292 248328 106304
rect 248380 106292 248386 106344
rect 253750 106292 253756 106344
rect 253808 106332 253814 106344
rect 253934 106332 253940 106344
rect 253808 106304 253940 106332
rect 253808 106292 253814 106304
rect 253934 106292 253940 106304
rect 253992 106292 253998 106344
rect 339678 106292 339684 106344
rect 339736 106332 339742 106344
rect 339862 106332 339868 106344
rect 339736 106304 339868 106332
rect 339736 106292 339742 106304
rect 339862 106292 339868 106304
rect 339920 106292 339926 106344
rect 343910 106292 343916 106344
rect 343968 106332 343974 106344
rect 344094 106332 344100 106344
rect 343968 106304 344100 106332
rect 343968 106292 343974 106304
rect 344094 106292 344100 106304
rect 344152 106292 344158 106344
rect 415210 106292 415216 106344
rect 415268 106292 415274 106344
rect 431678 106292 431684 106344
rect 431736 106292 431742 106344
rect 140774 106224 140780 106276
rect 140832 106264 140838 106276
rect 140958 106264 140964 106276
rect 140832 106236 140964 106264
rect 140832 106224 140838 106236
rect 140958 106224 140964 106236
rect 141016 106224 141022 106276
rect 156138 106224 156144 106276
rect 156196 106264 156202 106276
rect 156506 106264 156512 106276
rect 156196 106236 156512 106264
rect 156196 106224 156202 106236
rect 156506 106224 156512 106236
rect 156564 106224 156570 106276
rect 251266 106224 251272 106276
rect 251324 106264 251330 106276
rect 251450 106264 251456 106276
rect 251324 106236 251456 106264
rect 251324 106224 251330 106236
rect 251450 106224 251456 106236
rect 251508 106224 251514 106276
rect 341426 106224 341432 106276
rect 341484 106264 341490 106276
rect 341518 106264 341524 106276
rect 341484 106236 341524 106264
rect 341484 106224 341490 106236
rect 341518 106224 341524 106236
rect 341576 106224 341582 106276
rect 400582 106224 400588 106276
rect 400640 106264 400646 106276
rect 400858 106264 400864 106276
rect 400640 106236 400864 106264
rect 400640 106224 400646 106236
rect 400858 106224 400864 106236
rect 400916 106224 400922 106276
rect 403986 106224 403992 106276
rect 404044 106264 404050 106276
rect 404078 106264 404084 106276
rect 404044 106236 404084 106264
rect 404044 106224 404050 106236
rect 404078 106224 404084 106236
rect 404136 106224 404142 106276
rect 415228 106208 415256 106292
rect 431586 106224 431592 106276
rect 431644 106264 431650 106276
rect 431696 106264 431724 106292
rect 431644 106236 431724 106264
rect 431644 106224 431650 106236
rect 415210 106156 415216 106208
rect 415268 106156 415274 106208
rect 189074 104932 189080 104984
rect 189132 104972 189138 104984
rect 189166 104972 189172 104984
rect 189132 104944 189172 104972
rect 189132 104932 189138 104944
rect 189166 104932 189172 104944
rect 189224 104932 189230 104984
rect 161658 104864 161664 104916
rect 161716 104904 161722 104916
rect 161842 104904 161848 104916
rect 161716 104876 161848 104904
rect 161716 104864 161722 104876
rect 161842 104864 161848 104876
rect 161900 104864 161906 104916
rect 218238 104864 218244 104916
rect 218296 104904 218302 104916
rect 218330 104904 218336 104916
rect 218296 104876 218336 104904
rect 218296 104864 218302 104876
rect 218330 104864 218336 104876
rect 218388 104864 218394 104916
rect 233326 104864 233332 104916
rect 233384 104904 233390 104916
rect 233510 104904 233516 104916
rect 233384 104876 233516 104904
rect 233384 104864 233390 104876
rect 233510 104864 233516 104876
rect 233568 104864 233574 104916
rect 409322 104864 409328 104916
rect 409380 104904 409386 104916
rect 409414 104904 409420 104916
rect 409380 104876 409420 104904
rect 409380 104864 409386 104876
rect 409414 104864 409420 104876
rect 409472 104864 409478 104916
rect 140958 104796 140964 104848
rect 141016 104836 141022 104848
rect 141142 104836 141148 104848
rect 141016 104808 141148 104836
rect 141016 104796 141022 104808
rect 141142 104796 141148 104808
rect 141200 104796 141206 104848
rect 143626 104796 143632 104848
rect 143684 104836 143690 104848
rect 143902 104836 143908 104848
rect 143684 104808 143908 104836
rect 143684 104796 143690 104808
rect 143902 104796 143908 104808
rect 143960 104796 143966 104848
rect 148042 104796 148048 104848
rect 148100 104836 148106 104848
rect 148226 104836 148232 104848
rect 148100 104808 148232 104836
rect 148100 104796 148106 104808
rect 148226 104796 148232 104808
rect 148284 104796 148290 104848
rect 152090 104796 152096 104848
rect 152148 104836 152154 104848
rect 152182 104836 152188 104848
rect 152148 104808 152188 104836
rect 152148 104796 152154 104808
rect 152182 104796 152188 104808
rect 152240 104796 152246 104848
rect 221274 104796 221280 104848
rect 221332 104836 221338 104848
rect 221458 104836 221464 104848
rect 221332 104808 221464 104836
rect 221332 104796 221338 104808
rect 221458 104796 221464 104808
rect 221516 104796 221522 104848
rect 253566 104796 253572 104848
rect 253624 104836 253630 104848
rect 253750 104836 253756 104848
rect 253624 104808 253756 104836
rect 253624 104796 253630 104808
rect 253750 104796 253756 104808
rect 253808 104796 253814 104848
rect 275922 104796 275928 104848
rect 275980 104836 275986 104848
rect 276106 104836 276112 104848
rect 275980 104808 276112 104836
rect 275980 104796 275986 104808
rect 276106 104796 276112 104808
rect 276164 104796 276170 104848
rect 316862 104796 316868 104848
rect 316920 104836 316926 104848
rect 317046 104836 317052 104848
rect 316920 104808 317052 104836
rect 316920 104796 316926 104808
rect 317046 104796 317052 104808
rect 317104 104796 317110 104848
rect 420546 104796 420552 104848
rect 420604 104836 420610 104848
rect 420638 104836 420644 104848
rect 420604 104808 420644 104836
rect 420604 104796 420610 104808
rect 420638 104796 420644 104808
rect 420696 104796 420702 104848
rect 425974 104796 425980 104848
rect 426032 104836 426038 104848
rect 426158 104836 426164 104848
rect 426032 104808 426164 104836
rect 426032 104796 426038 104808
rect 426158 104796 426164 104808
rect 426216 104796 426222 104848
rect 431402 104796 431408 104848
rect 431460 104836 431466 104848
rect 431678 104836 431684 104848
rect 431460 104808 431684 104836
rect 431460 104796 431466 104808
rect 431678 104796 431684 104808
rect 431736 104796 431742 104848
rect 179598 103436 179604 103488
rect 179656 103476 179662 103488
rect 179690 103476 179696 103488
rect 179656 103448 179696 103476
rect 179656 103436 179662 103448
rect 179690 103436 179696 103448
rect 179748 103436 179754 103488
rect 189166 103436 189172 103488
rect 189224 103476 189230 103488
rect 189534 103476 189540 103488
rect 189224 103448 189540 103476
rect 189224 103436 189230 103448
rect 189534 103436 189540 103448
rect 189592 103436 189598 103488
rect 233326 103436 233332 103488
rect 233384 103476 233390 103488
rect 233510 103476 233516 103488
rect 233384 103448 233516 103476
rect 233384 103436 233390 103448
rect 233510 103436 233516 103448
rect 233568 103436 233574 103488
rect 414934 103436 414940 103488
rect 414992 103476 414998 103488
rect 415118 103476 415124 103488
rect 414992 103448 415124 103476
rect 414992 103436 414998 103448
rect 415118 103436 415124 103448
rect 415176 103436 415182 103488
rect 133138 99424 133144 99476
rect 133196 99424 133202 99476
rect 138106 99424 138112 99476
rect 138164 99424 138170 99476
rect 162946 99424 162952 99476
rect 163004 99424 163010 99476
rect 216950 99424 216956 99476
rect 217008 99424 217014 99476
rect 227898 99464 227904 99476
rect 227824 99436 227904 99464
rect 133156 99340 133184 99424
rect 138124 99340 138152 99424
rect 162964 99340 162992 99424
rect 168374 99356 168380 99408
rect 168432 99396 168438 99408
rect 168558 99396 168564 99408
rect 168432 99368 168564 99396
rect 168432 99356 168438 99368
rect 168558 99356 168564 99368
rect 168616 99356 168622 99408
rect 179598 99356 179604 99408
rect 179656 99396 179662 99408
rect 179656 99368 179736 99396
rect 179656 99356 179662 99368
rect 179708 99340 179736 99368
rect 216968 99340 216996 99424
rect 227824 99340 227852 99436
rect 227898 99424 227904 99436
rect 227956 99424 227962 99476
rect 383286 99464 383292 99476
rect 383212 99436 383292 99464
rect 249886 99356 249892 99408
rect 249944 99356 249950 99408
rect 313918 99356 313924 99408
rect 313976 99396 313982 99408
rect 314102 99396 314108 99408
rect 313976 99368 314108 99396
rect 313976 99356 313982 99368
rect 314102 99356 314108 99368
rect 314160 99356 314166 99408
rect 133138 99288 133144 99340
rect 133196 99288 133202 99340
rect 138106 99288 138112 99340
rect 138164 99288 138170 99340
rect 162946 99288 162952 99340
rect 163004 99288 163010 99340
rect 179690 99288 179696 99340
rect 179748 99288 179754 99340
rect 216950 99288 216956 99340
rect 217008 99288 217014 99340
rect 227806 99288 227812 99340
rect 227864 99288 227870 99340
rect 249904 99328 249932 99356
rect 383212 99340 383240 99436
rect 383286 99424 383292 99436
rect 383344 99424 383350 99476
rect 249978 99328 249984 99340
rect 249904 99300 249984 99328
rect 249978 99288 249984 99300
rect 250036 99288 250042 99340
rect 383194 99288 383200 99340
rect 383252 99288 383258 99340
rect 173802 98676 173808 98728
rect 173860 98716 173866 98728
rect 173986 98716 173992 98728
rect 173860 98688 173992 98716
rect 173860 98676 173866 98688
rect 173986 98676 173992 98688
rect 174044 98676 174050 98728
rect 251266 96636 251272 96688
rect 251324 96676 251330 96688
rect 251450 96676 251456 96688
rect 251324 96648 251456 96676
rect 251324 96636 251330 96648
rect 251450 96636 251456 96648
rect 251508 96636 251514 96688
rect 341518 96636 341524 96688
rect 341576 96636 341582 96688
rect 400582 96636 400588 96688
rect 400640 96676 400646 96688
rect 400766 96676 400772 96688
rect 400640 96648 400772 96676
rect 400640 96636 400646 96648
rect 400766 96636 400772 96648
rect 400824 96636 400830 96688
rect 168374 96568 168380 96620
rect 168432 96608 168438 96620
rect 168558 96608 168564 96620
rect 168432 96580 168564 96608
rect 168432 96568 168438 96580
rect 168558 96568 168564 96580
rect 168616 96568 168622 96620
rect 180978 96568 180984 96620
rect 181036 96608 181042 96620
rect 181162 96608 181168 96620
rect 181036 96580 181168 96608
rect 181036 96568 181042 96580
rect 181162 96568 181168 96580
rect 181220 96568 181226 96620
rect 186038 96568 186044 96620
rect 186096 96608 186102 96620
rect 186222 96608 186228 96620
rect 186096 96580 186228 96608
rect 186096 96568 186102 96580
rect 186222 96568 186228 96580
rect 186280 96568 186286 96620
rect 203058 96568 203064 96620
rect 203116 96608 203122 96620
rect 203242 96608 203248 96620
rect 203116 96580 203248 96608
rect 203116 96568 203122 96580
rect 203242 96568 203248 96580
rect 203300 96568 203306 96620
rect 204622 96568 204628 96620
rect 204680 96608 204686 96620
rect 204806 96608 204812 96620
rect 204680 96580 204812 96608
rect 204680 96568 204686 96580
rect 204806 96568 204812 96580
rect 204864 96568 204870 96620
rect 209958 96568 209964 96620
rect 210016 96608 210022 96620
rect 210142 96608 210148 96620
rect 210016 96580 210148 96608
rect 210016 96568 210022 96580
rect 210142 96568 210148 96580
rect 210200 96568 210206 96620
rect 274450 96568 274456 96620
rect 274508 96608 274514 96620
rect 274726 96608 274732 96620
rect 274508 96580 274732 96608
rect 274508 96568 274514 96580
rect 274726 96568 274732 96580
rect 274784 96568 274790 96620
rect 341426 96568 341432 96620
rect 341484 96608 341490 96620
rect 341536 96608 341564 96636
rect 341484 96580 341564 96608
rect 341484 96568 341490 96580
rect 343910 96568 343916 96620
rect 343968 96608 343974 96620
rect 344094 96608 344100 96620
rect 343968 96580 344100 96608
rect 343968 96568 343974 96580
rect 344094 96568 344100 96580
rect 344152 96568 344158 96620
rect 382918 96568 382924 96620
rect 382976 96608 382982 96620
rect 383194 96608 383200 96620
rect 382976 96580 383200 96608
rect 382976 96568 382982 96580
rect 383194 96568 383200 96580
rect 383252 96568 383258 96620
rect 403710 96568 403716 96620
rect 403768 96608 403774 96620
rect 403986 96608 403992 96620
rect 403768 96580 403992 96608
rect 403768 96568 403774 96580
rect 403986 96568 403992 96580
rect 404044 96568 404050 96620
rect 190638 96500 190644 96552
rect 190696 96540 190702 96552
rect 190730 96540 190736 96552
rect 190696 96512 190736 96540
rect 190696 96500 190702 96512
rect 190730 96500 190736 96512
rect 190788 96500 190794 96552
rect 148042 95208 148048 95260
rect 148100 95248 148106 95260
rect 148226 95248 148232 95260
rect 148100 95220 148232 95248
rect 148100 95208 148106 95220
rect 148226 95208 148232 95220
rect 148284 95208 148290 95260
rect 150710 95208 150716 95260
rect 150768 95248 150774 95260
rect 150986 95248 150992 95260
rect 150768 95220 150992 95248
rect 150768 95208 150774 95220
rect 150986 95208 150992 95220
rect 151044 95208 151050 95260
rect 151814 95208 151820 95260
rect 151872 95248 151878 95260
rect 152090 95248 152096 95260
rect 151872 95220 152096 95248
rect 151872 95208 151878 95220
rect 152090 95208 152096 95220
rect 152148 95208 152154 95260
rect 215570 95208 215576 95260
rect 215628 95248 215634 95260
rect 215938 95248 215944 95260
rect 215628 95220 215944 95248
rect 215628 95208 215634 95220
rect 215938 95208 215944 95220
rect 215996 95208 216002 95260
rect 216950 95208 216956 95260
rect 217008 95248 217014 95260
rect 217042 95248 217048 95260
rect 217008 95220 217048 95248
rect 217008 95208 217014 95220
rect 217042 95208 217048 95220
rect 217100 95208 217106 95260
rect 218330 95208 218336 95260
rect 218388 95248 218394 95260
rect 218422 95248 218428 95260
rect 218388 95220 218428 95248
rect 218388 95208 218394 95220
rect 218422 95208 218428 95220
rect 218480 95208 218486 95260
rect 233510 95208 233516 95260
rect 233568 95208 233574 95260
rect 253566 95208 253572 95260
rect 253624 95248 253630 95260
rect 253750 95248 253756 95260
rect 253624 95220 253756 95248
rect 253624 95208 253630 95220
rect 253750 95208 253756 95220
rect 253808 95208 253814 95260
rect 275922 95208 275928 95260
rect 275980 95248 275986 95260
rect 276014 95248 276020 95260
rect 275980 95220 276020 95248
rect 275980 95208 275986 95220
rect 276014 95208 276020 95220
rect 276072 95208 276078 95260
rect 316862 95208 316868 95260
rect 316920 95248 316926 95260
rect 317046 95248 317052 95260
rect 316920 95220 317052 95248
rect 316920 95208 316926 95220
rect 317046 95208 317052 95220
rect 317104 95208 317110 95260
rect 341426 95208 341432 95260
rect 341484 95248 341490 95260
rect 341518 95248 341524 95260
rect 341484 95220 341524 95248
rect 341484 95208 341490 95220
rect 341518 95208 341524 95220
rect 341576 95208 341582 95260
rect 409322 95208 409328 95260
rect 409380 95248 409386 95260
rect 409598 95248 409604 95260
rect 409380 95220 409604 95248
rect 409380 95208 409386 95220
rect 409598 95208 409604 95220
rect 409656 95208 409662 95260
rect 420546 95208 420552 95260
rect 420604 95248 420610 95260
rect 420730 95248 420736 95260
rect 420604 95220 420736 95248
rect 420604 95208 420610 95220
rect 420730 95208 420736 95220
rect 420788 95208 420794 95260
rect 185946 95140 185952 95192
rect 186004 95180 186010 95192
rect 186038 95180 186044 95192
rect 186004 95152 186044 95180
rect 186004 95140 186010 95152
rect 186038 95140 186044 95152
rect 186096 95140 186102 95192
rect 233528 95124 233556 95208
rect 431402 95140 431408 95192
rect 431460 95180 431466 95192
rect 431494 95180 431500 95192
rect 431460 95152 431500 95180
rect 431460 95140 431466 95152
rect 431494 95140 431500 95152
rect 431552 95140 431558 95192
rect 189350 95072 189356 95124
rect 189408 95112 189414 95124
rect 189534 95112 189540 95124
rect 189408 95084 189540 95112
rect 189408 95072 189414 95084
rect 189534 95072 189540 95084
rect 189592 95072 189598 95124
rect 233510 95072 233516 95124
rect 233568 95072 233574 95124
rect 276014 95072 276020 95124
rect 276072 95112 276078 95124
rect 276290 95112 276296 95124
rect 276072 95084 276296 95112
rect 276072 95072 276078 95084
rect 276290 95072 276296 95084
rect 276348 95072 276354 95124
rect 173802 93848 173808 93900
rect 173860 93888 173866 93900
rect 173986 93888 173992 93900
rect 173860 93860 173992 93888
rect 173860 93848 173866 93860
rect 173986 93848 173992 93860
rect 174044 93848 174050 93900
rect 3418 93780 3424 93832
rect 3476 93820 3482 93832
rect 14458 93820 14464 93832
rect 3476 93792 14464 93820
rect 3476 93780 3482 93792
rect 14458 93780 14464 93792
rect 14516 93780 14522 93832
rect 150526 91740 150532 91792
rect 150584 91780 150590 91792
rect 150710 91780 150716 91792
rect 150584 91752 150716 91780
rect 150584 91740 150590 91752
rect 150710 91740 150716 91752
rect 150768 91740 150774 91792
rect 400766 91740 400772 91792
rect 400824 91780 400830 91792
rect 401042 91780 401048 91792
rect 400824 91752 401048 91780
rect 400824 91740 400830 91752
rect 401042 91740 401048 91752
rect 401100 91740 401106 91792
rect 185026 89808 185032 89820
rect 184952 89780 185032 89808
rect 184952 89684 184980 89780
rect 185026 89768 185032 89780
rect 185084 89768 185090 89820
rect 227806 89700 227812 89752
rect 227864 89700 227870 89752
rect 341334 89700 341340 89752
rect 341392 89740 341398 89752
rect 341518 89740 341524 89752
rect 341392 89712 341524 89740
rect 341392 89700 341398 89712
rect 341518 89700 341524 89712
rect 341576 89700 341582 89752
rect 409506 89700 409512 89752
rect 409564 89740 409570 89752
rect 409564 89712 409644 89740
rect 409564 89700 409570 89712
rect 180978 89632 180984 89684
rect 181036 89672 181042 89684
rect 181162 89672 181168 89684
rect 181036 89644 181168 89672
rect 181036 89632 181042 89644
rect 181162 89632 181168 89644
rect 181220 89632 181226 89684
rect 184934 89632 184940 89684
rect 184992 89632 184998 89684
rect 227824 89604 227852 89700
rect 409616 89684 409644 89712
rect 415118 89700 415124 89752
rect 415176 89700 415182 89752
rect 251266 89632 251272 89684
rect 251324 89632 251330 89684
rect 409598 89632 409604 89684
rect 409656 89632 409662 89684
rect 227898 89604 227904 89616
rect 227824 89576 227904 89604
rect 227898 89564 227904 89576
rect 227956 89564 227962 89616
rect 251284 89604 251312 89632
rect 415136 89616 415164 89700
rect 251358 89604 251364 89616
rect 251284 89576 251364 89604
rect 251358 89564 251364 89576
rect 251416 89564 251422 89616
rect 415118 89564 415124 89616
rect 415176 89564 415182 89616
rect 133506 88272 133512 88324
rect 133564 88312 133570 88324
rect 580166 88312 580172 88324
rect 133564 88284 580172 88312
rect 133564 88272 133570 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 140866 86980 140872 87032
rect 140924 87020 140930 87032
rect 140958 87020 140964 87032
rect 140924 86992 140964 87020
rect 140924 86980 140930 86992
rect 140958 86980 140964 86992
rect 141016 86980 141022 87032
rect 143626 86980 143632 87032
rect 143684 87020 143690 87032
rect 143902 87020 143908 87032
rect 143684 86992 143908 87020
rect 143684 86980 143690 86992
rect 143902 86980 143908 86992
rect 143960 86980 143966 87032
rect 147858 86980 147864 87032
rect 147916 87020 147922 87032
rect 148042 87020 148048 87032
rect 147916 86992 148048 87020
rect 147916 86980 147922 86992
rect 148042 86980 148048 86992
rect 148100 86980 148106 87032
rect 343910 86980 343916 87032
rect 343968 87020 343974 87032
rect 344094 87020 344100 87032
rect 343968 86992 344100 87020
rect 343968 86980 343974 86992
rect 344094 86980 344100 86992
rect 344152 86980 344158 87032
rect 382918 86980 382924 87032
rect 382976 87020 382982 87032
rect 383102 87020 383108 87032
rect 382976 86992 383108 87020
rect 382976 86980 382982 86992
rect 383102 86980 383108 86992
rect 383160 86980 383166 87032
rect 403710 86980 403716 87032
rect 403768 87020 403774 87032
rect 403894 87020 403900 87032
rect 403768 86992 403900 87020
rect 403768 86980 403774 86992
rect 403894 86980 403900 86992
rect 403952 86980 403958 87032
rect 151814 86912 151820 86964
rect 151872 86952 151878 86964
rect 151906 86952 151912 86964
rect 151872 86924 151912 86952
rect 151872 86912 151878 86924
rect 151906 86912 151912 86924
rect 151964 86912 151970 86964
rect 184750 86912 184756 86964
rect 184808 86952 184814 86964
rect 184934 86952 184940 86964
rect 184808 86924 184940 86952
rect 184808 86912 184814 86924
rect 184934 86912 184940 86924
rect 184992 86912 184998 86964
rect 203242 86912 203248 86964
rect 203300 86952 203306 86964
rect 203426 86952 203432 86964
rect 203300 86924 203432 86952
rect 203300 86912 203306 86924
rect 203426 86912 203432 86924
rect 203484 86912 203490 86964
rect 215478 86912 215484 86964
rect 215536 86952 215542 86964
rect 215570 86952 215576 86964
rect 215536 86924 215576 86952
rect 215536 86912 215542 86924
rect 215570 86912 215576 86924
rect 215628 86912 215634 86964
rect 216950 86912 216956 86964
rect 217008 86952 217014 86964
rect 217042 86952 217048 86964
rect 217008 86924 217048 86952
rect 217008 86912 217014 86924
rect 217042 86912 217048 86924
rect 217100 86912 217106 86964
rect 218238 86912 218244 86964
rect 218296 86952 218302 86964
rect 218330 86952 218336 86964
rect 218296 86924 218336 86952
rect 218296 86912 218302 86924
rect 218330 86912 218336 86924
rect 218388 86912 218394 86964
rect 219710 86912 219716 86964
rect 219768 86952 219774 86964
rect 219802 86952 219808 86964
rect 219768 86924 219808 86952
rect 219768 86912 219774 86924
rect 219802 86912 219808 86924
rect 219860 86912 219866 86964
rect 274634 86912 274640 86964
rect 274692 86952 274698 86964
rect 274818 86952 274824 86964
rect 274692 86924 274824 86952
rect 274692 86912 274698 86924
rect 274818 86912 274824 86924
rect 274876 86912 274882 86964
rect 316954 86912 316960 86964
rect 317012 86952 317018 86964
rect 317138 86952 317144 86964
rect 317012 86924 317144 86952
rect 317012 86912 317018 86924
rect 317138 86912 317144 86924
rect 317196 86912 317202 86964
rect 420546 86912 420552 86964
rect 420604 86952 420610 86964
rect 420638 86952 420644 86964
rect 420604 86924 420644 86952
rect 420604 86912 420610 86924
rect 420638 86912 420644 86924
rect 420696 86912 420702 86964
rect 403894 86844 403900 86896
rect 403952 86884 403958 86896
rect 403986 86884 403992 86896
rect 403952 86856 403992 86884
rect 403952 86844 403958 86856
rect 403986 86844 403992 86856
rect 404044 86844 404050 86896
rect 185946 85552 185952 85604
rect 186004 85592 186010 85604
rect 186222 85592 186228 85604
rect 186004 85564 186228 85592
rect 186004 85552 186010 85564
rect 186222 85552 186228 85564
rect 186280 85552 186286 85604
rect 189258 85552 189264 85604
rect 189316 85592 189322 85604
rect 189350 85592 189356 85604
rect 189316 85564 189356 85592
rect 189316 85552 189322 85564
rect 189350 85552 189356 85564
rect 189408 85552 189414 85604
rect 431494 85552 431500 85604
rect 431552 85592 431558 85604
rect 431586 85592 431592 85604
rect 431552 85564 431592 85592
rect 431552 85552 431558 85564
rect 431586 85552 431592 85564
rect 431644 85552 431650 85604
rect 143626 85484 143632 85536
rect 143684 85524 143690 85536
rect 143810 85524 143816 85536
rect 143684 85496 143816 85524
rect 143684 85484 143690 85496
rect 143810 85484 143816 85496
rect 143868 85484 143874 85536
rect 144822 85484 144828 85536
rect 144880 85524 144886 85536
rect 145098 85524 145104 85536
rect 144880 85496 145104 85524
rect 144880 85484 144886 85496
rect 145098 85484 145104 85496
rect 145156 85484 145162 85536
rect 218238 85484 218244 85536
rect 218296 85524 218302 85536
rect 218422 85524 218428 85536
rect 218296 85496 218428 85524
rect 218296 85484 218302 85496
rect 218422 85484 218428 85496
rect 218480 85484 218486 85536
rect 227530 85484 227536 85536
rect 227588 85524 227594 85536
rect 227898 85524 227904 85536
rect 227588 85496 227904 85524
rect 227588 85484 227594 85496
rect 227898 85484 227904 85496
rect 227956 85484 227962 85536
rect 253566 85484 253572 85536
rect 253624 85524 253630 85536
rect 253750 85524 253756 85536
rect 253624 85496 253756 85524
rect 253624 85484 253630 85496
rect 253750 85484 253756 85496
rect 253808 85484 253814 85536
rect 276106 85484 276112 85536
rect 276164 85524 276170 85536
rect 276198 85524 276204 85536
rect 276164 85496 276204 85524
rect 276164 85484 276170 85496
rect 276198 85484 276204 85496
rect 276256 85484 276262 85536
rect 313918 85484 313924 85536
rect 313976 85524 313982 85536
rect 314010 85524 314016 85536
rect 313976 85496 314016 85524
rect 313976 85484 313982 85496
rect 314010 85484 314016 85496
rect 314068 85484 314074 85536
rect 339126 85484 339132 85536
rect 339184 85524 339190 85536
rect 339218 85524 339224 85536
rect 339184 85496 339224 85524
rect 339184 85484 339190 85496
rect 339218 85484 339224 85496
rect 339276 85484 339282 85536
rect 400766 85484 400772 85536
rect 400824 85524 400830 85536
rect 400950 85524 400956 85536
rect 400824 85496 400956 85524
rect 400824 85484 400830 85496
rect 400950 85484 400956 85496
rect 401008 85484 401014 85536
rect 173802 84124 173808 84176
rect 173860 84164 173866 84176
rect 173986 84164 173992 84176
rect 173860 84136 173992 84164
rect 173860 84124 173866 84136
rect 173986 84124 173992 84136
rect 174044 84124 174050 84176
rect 276014 84124 276020 84176
rect 276072 84164 276078 84176
rect 276198 84164 276204 84176
rect 276072 84136 276204 84164
rect 276072 84124 276078 84136
rect 276198 84124 276204 84136
rect 276256 84124 276262 84176
rect 314010 84124 314016 84176
rect 314068 84164 314074 84176
rect 314194 84164 314200 84176
rect 314068 84136 314200 84164
rect 314068 84124 314074 84136
rect 314194 84124 314200 84136
rect 314252 84124 314258 84176
rect 338942 84124 338948 84176
rect 339000 84164 339006 84176
rect 339126 84164 339132 84176
rect 339000 84136 339132 84164
rect 339000 84124 339006 84136
rect 339126 84124 339132 84136
rect 339184 84124 339190 84176
rect 415026 84124 415032 84176
rect 415084 84164 415090 84176
rect 415118 84164 415124 84176
rect 415084 84136 415124 84164
rect 415084 84124 415090 84136
rect 415118 84124 415124 84136
rect 415176 84124 415182 84176
rect 164510 82084 164516 82136
rect 164568 82124 164574 82136
rect 164568 82096 164648 82124
rect 164568 82084 164574 82096
rect 164620 82068 164648 82096
rect 164602 82016 164608 82068
rect 164660 82016 164666 82068
rect 426066 80656 426072 80708
rect 426124 80696 426130 80708
rect 426158 80696 426164 80708
rect 426124 80668 426164 80696
rect 426124 80656 426130 80668
rect 426158 80656 426164 80668
rect 426216 80656 426222 80708
rect 196158 80180 196164 80232
rect 196216 80180 196222 80232
rect 196176 80096 196204 80180
rect 240318 80152 240324 80164
rect 240244 80124 240324 80152
rect 240244 80096 240272 80124
rect 240318 80112 240324 80124
rect 240376 80112 240382 80164
rect 249886 80152 249892 80164
rect 249812 80124 249892 80152
rect 249812 80096 249840 80124
rect 249886 80112 249892 80124
rect 249944 80112 249950 80164
rect 196158 80044 196164 80096
rect 196216 80044 196222 80096
rect 240226 80044 240232 80096
rect 240284 80044 240290 80096
rect 249794 80044 249800 80096
rect 249852 80044 249858 80096
rect 431586 80044 431592 80096
rect 431644 80084 431650 80096
rect 431770 80084 431776 80096
rect 431644 80056 431776 80084
rect 431644 80044 431650 80056
rect 431770 80044 431776 80056
rect 431828 80044 431834 80096
rect 3142 79976 3148 80028
rect 3200 80016 3206 80028
rect 436370 80016 436376 80028
rect 3200 79988 436376 80016
rect 3200 79976 3206 79988
rect 436370 79976 436376 79988
rect 436428 79976 436434 80028
rect 420546 77324 420552 77376
rect 420604 77364 420610 77376
rect 420730 77364 420736 77376
rect 420604 77336 420736 77364
rect 420604 77324 420610 77336
rect 420730 77324 420736 77336
rect 420788 77324 420794 77376
rect 183646 77256 183652 77308
rect 183704 77296 183710 77308
rect 183738 77296 183744 77308
rect 183704 77268 183744 77296
rect 183704 77256 183710 77268
rect 183738 77256 183744 77268
rect 183796 77256 183802 77308
rect 184750 77256 184756 77308
rect 184808 77296 184814 77308
rect 185026 77296 185032 77308
rect 184808 77268 185032 77296
rect 184808 77256 184814 77268
rect 185026 77256 185032 77268
rect 185084 77256 185090 77308
rect 189074 77256 189080 77308
rect 189132 77296 189138 77308
rect 189258 77296 189264 77308
rect 189132 77268 189264 77296
rect 189132 77256 189138 77268
rect 189258 77256 189264 77268
rect 189316 77256 189322 77308
rect 203058 77256 203064 77308
rect 203116 77296 203122 77308
rect 203426 77296 203432 77308
rect 203116 77268 203432 77296
rect 203116 77256 203122 77268
rect 203426 77256 203432 77268
rect 203484 77256 203490 77308
rect 204346 77256 204352 77308
rect 204404 77296 204410 77308
rect 204622 77296 204628 77308
rect 204404 77268 204628 77296
rect 204404 77256 204410 77268
rect 204622 77256 204628 77268
rect 204680 77256 204686 77308
rect 316954 77256 316960 77308
rect 317012 77296 317018 77308
rect 317230 77296 317236 77308
rect 317012 77268 317236 77296
rect 317012 77256 317018 77268
rect 317230 77256 317236 77268
rect 317288 77256 317294 77308
rect 128906 77188 128912 77240
rect 128964 77228 128970 77240
rect 128998 77228 129004 77240
rect 128964 77200 129004 77228
rect 128964 77188 128970 77200
rect 128998 77188 129004 77200
rect 129056 77188 129062 77240
rect 132310 77188 132316 77240
rect 132368 77228 132374 77240
rect 580166 77228 580172 77240
rect 132368 77200 580172 77228
rect 132368 77188 132374 77200
rect 580166 77188 580172 77200
rect 580224 77188 580230 77240
rect 186222 75964 186228 76016
rect 186280 75964 186286 76016
rect 186314 75964 186320 76016
rect 186372 75964 186378 76016
rect 186406 75964 186412 76016
rect 186464 75964 186470 76016
rect 186498 75964 186504 76016
rect 186556 75964 186562 76016
rect 143626 75896 143632 75948
rect 143684 75936 143690 75948
rect 143810 75936 143816 75948
rect 143684 75908 143816 75936
rect 143684 75896 143690 75908
rect 143810 75896 143816 75908
rect 143868 75896 143874 75948
rect 144822 75896 144828 75948
rect 144880 75936 144886 75948
rect 145006 75936 145012 75948
rect 144880 75908 145012 75936
rect 144880 75896 144886 75908
rect 145006 75896 145012 75908
rect 145064 75896 145070 75948
rect 186240 75880 186268 75964
rect 186332 75880 186360 75964
rect 186424 75880 186452 75964
rect 186516 75880 186544 75964
rect 218238 75896 218244 75948
rect 218296 75936 218302 75948
rect 218422 75936 218428 75948
rect 218296 75908 218428 75936
rect 218296 75896 218302 75908
rect 218422 75896 218428 75908
rect 218480 75896 218486 75948
rect 227530 75896 227536 75948
rect 227588 75936 227594 75948
rect 227714 75936 227720 75948
rect 227588 75908 227720 75936
rect 227588 75896 227594 75908
rect 227714 75896 227720 75908
rect 227772 75896 227778 75948
rect 244274 75896 244280 75948
rect 244332 75936 244338 75948
rect 244458 75936 244464 75948
rect 244332 75908 244464 75936
rect 244332 75896 244338 75908
rect 244458 75896 244464 75908
rect 244516 75896 244522 75948
rect 253566 75896 253572 75948
rect 253624 75936 253630 75948
rect 253750 75936 253756 75948
rect 253624 75908 253756 75936
rect 253624 75896 253630 75908
rect 253750 75896 253756 75908
rect 253808 75896 253814 75948
rect 341702 75896 341708 75948
rect 341760 75936 341766 75948
rect 341886 75936 341892 75948
rect 341760 75908 341892 75936
rect 341760 75896 341766 75908
rect 341886 75896 341892 75908
rect 341944 75896 341950 75948
rect 186222 75828 186228 75880
rect 186280 75828 186286 75880
rect 186314 75828 186320 75880
rect 186372 75828 186378 75880
rect 186406 75828 186412 75880
rect 186464 75828 186470 75880
rect 186498 75828 186504 75880
rect 186556 75828 186562 75880
rect 189074 75828 189080 75880
rect 189132 75868 189138 75880
rect 189166 75868 189172 75880
rect 189132 75840 189172 75868
rect 189132 75828 189138 75840
rect 189166 75828 189172 75840
rect 189224 75828 189230 75880
rect 220998 75828 221004 75880
rect 221056 75868 221062 75880
rect 221274 75868 221280 75880
rect 221056 75840 221280 75868
rect 221056 75828 221062 75840
rect 221274 75828 221280 75840
rect 221332 75828 221338 75880
rect 249794 75828 249800 75880
rect 249852 75868 249858 75880
rect 249886 75868 249892 75880
rect 249852 75840 249892 75868
rect 249852 75828 249858 75840
rect 249886 75828 249892 75840
rect 249944 75828 249950 75880
rect 431586 75828 431592 75880
rect 431644 75868 431650 75880
rect 431770 75868 431776 75880
rect 431644 75840 431776 75868
rect 431644 75828 431650 75840
rect 431770 75828 431776 75840
rect 431828 75828 431834 75880
rect 233234 74604 233240 74656
rect 233292 74644 233298 74656
rect 233694 74644 233700 74656
rect 233292 74616 233700 74644
rect 233292 74604 233298 74616
rect 233694 74604 233700 74616
rect 233752 74604 233758 74656
rect 173802 74536 173808 74588
rect 173860 74576 173866 74588
rect 173894 74576 173900 74588
rect 173860 74548 173900 74576
rect 173860 74536 173866 74548
rect 173894 74536 173900 74548
rect 173952 74536 173958 74588
rect 186222 74536 186228 74588
rect 186280 74576 186286 74588
rect 186590 74576 186596 74588
rect 186280 74548 186596 74576
rect 186280 74536 186286 74548
rect 186590 74536 186596 74548
rect 186648 74536 186654 74588
rect 275922 74536 275928 74588
rect 275980 74576 275986 74588
rect 276014 74576 276020 74588
rect 275980 74548 276020 74576
rect 275980 74536 275986 74548
rect 276014 74536 276020 74548
rect 276072 74536 276078 74588
rect 414934 74536 414940 74588
rect 414992 74576 414998 74588
rect 415026 74576 415032 74588
rect 414992 74548 415032 74576
rect 414992 74536 414998 74548
rect 415026 74536 415032 74548
rect 415084 74536 415090 74588
rect 426066 74468 426072 74520
rect 426124 74508 426130 74520
rect 426434 74508 426440 74520
rect 426124 74480 426440 74508
rect 426124 74468 426130 74480
rect 426434 74468 426440 74480
rect 426492 74468 426498 74520
rect 274726 72428 274732 72480
rect 274784 72468 274790 72480
rect 275094 72468 275100 72480
rect 274784 72440 275100 72468
rect 274784 72428 274790 72440
rect 275094 72428 275100 72440
rect 275152 72428 275158 72480
rect 138106 71068 138112 71120
rect 138164 71108 138170 71120
rect 138290 71108 138296 71120
rect 138164 71080 138296 71108
rect 138164 71068 138170 71080
rect 138290 71068 138296 71080
rect 138348 71068 138354 71120
rect 162946 71068 162952 71120
rect 163004 71108 163010 71120
rect 163130 71108 163136 71120
rect 163004 71080 163136 71108
rect 163004 71068 163010 71080
rect 163130 71068 163136 71080
rect 163188 71068 163194 71120
rect 184750 71068 184756 71120
rect 184808 71108 184814 71120
rect 185026 71108 185032 71120
rect 184808 71080 185032 71108
rect 184808 71068 184814 71080
rect 185026 71068 185032 71080
rect 185084 71068 185090 71120
rect 189166 70388 189172 70440
rect 189224 70388 189230 70440
rect 249886 70388 249892 70440
rect 249944 70388 249950 70440
rect 400950 70388 400956 70440
rect 401008 70428 401014 70440
rect 401008 70400 401088 70428
rect 401008 70388 401014 70400
rect 189184 70304 189212 70388
rect 203058 70320 203064 70372
rect 203116 70320 203122 70372
rect 249904 70360 249932 70388
rect 401060 70372 401088 70400
rect 249978 70360 249984 70372
rect 249904 70332 249984 70360
rect 249978 70320 249984 70332
rect 250036 70320 250042 70372
rect 401042 70320 401048 70372
rect 401100 70320 401106 70372
rect 189166 70252 189172 70304
rect 189224 70252 189230 70304
rect 203076 70292 203104 70320
rect 203150 70292 203156 70304
rect 203076 70264 203156 70292
rect 203150 70252 203156 70264
rect 203208 70252 203214 70304
rect 179598 67668 179604 67720
rect 179656 67668 179662 67720
rect 181070 67668 181076 67720
rect 181128 67668 181134 67720
rect 133138 67600 133144 67652
rect 133196 67640 133202 67652
rect 133230 67640 133236 67652
rect 133196 67612 133236 67640
rect 133196 67600 133202 67612
rect 133230 67600 133236 67612
rect 133288 67600 133294 67652
rect 161566 67600 161572 67652
rect 161624 67640 161630 67652
rect 161658 67640 161664 67652
rect 161624 67612 161664 67640
rect 161624 67600 161630 67612
rect 161658 67600 161664 67612
rect 161716 67600 161722 67652
rect 128814 67532 128820 67584
rect 128872 67572 128878 67584
rect 129090 67572 129096 67584
rect 128872 67544 129096 67572
rect 128872 67532 128878 67544
rect 129090 67532 129096 67544
rect 129148 67532 129154 67584
rect 179616 67504 179644 67668
rect 179690 67504 179696 67516
rect 179616 67476 179696 67504
rect 179690 67464 179696 67476
rect 179748 67464 179754 67516
rect 181088 67504 181116 67668
rect 209866 67600 209872 67652
rect 209924 67640 209930 67652
rect 209958 67640 209964 67652
rect 209924 67612 209964 67640
rect 209924 67600 209930 67612
rect 209958 67600 209964 67612
rect 210016 67600 210022 67652
rect 274910 67600 274916 67652
rect 274968 67640 274974 67652
rect 275094 67640 275100 67652
rect 274968 67612 275100 67640
rect 274968 67600 274974 67612
rect 275094 67600 275100 67612
rect 275152 67600 275158 67652
rect 341518 67600 341524 67652
rect 341576 67640 341582 67652
rect 341886 67640 341892 67652
rect 341576 67612 341892 67640
rect 341576 67600 341582 67612
rect 341886 67600 341892 67612
rect 341944 67600 341950 67652
rect 383286 67600 383292 67652
rect 383344 67640 383350 67652
rect 383654 67640 383660 67652
rect 383344 67612 383660 67640
rect 383344 67600 383350 67612
rect 383654 67600 383660 67612
rect 383712 67600 383718 67652
rect 400950 67600 400956 67652
rect 401008 67640 401014 67652
rect 401042 67640 401048 67652
rect 401008 67612 401048 67640
rect 401008 67600 401014 67612
rect 401042 67600 401048 67612
rect 401100 67600 401106 67652
rect 409506 67600 409512 67652
rect 409564 67640 409570 67652
rect 409598 67640 409604 67652
rect 409564 67612 409604 67640
rect 409564 67600 409570 67612
rect 409598 67600 409604 67612
rect 409656 67600 409662 67652
rect 420638 67600 420644 67652
rect 420696 67640 420702 67652
rect 421006 67640 421012 67652
rect 420696 67612 421012 67640
rect 420696 67600 420702 67612
rect 421006 67600 421012 67612
rect 421064 67600 421070 67652
rect 203058 67532 203064 67584
rect 203116 67572 203122 67584
rect 203150 67572 203156 67584
rect 203116 67544 203156 67572
rect 203116 67532 203122 67544
rect 203150 67532 203156 67544
rect 203208 67532 203214 67584
rect 238938 67532 238944 67584
rect 238996 67572 239002 67584
rect 239122 67572 239128 67584
rect 238996 67544 239128 67572
rect 238996 67532 239002 67544
rect 239122 67532 239128 67544
rect 239180 67532 239186 67584
rect 181162 67504 181168 67516
rect 181088 67476 181168 67504
rect 181162 67464 181168 67476
rect 181220 67464 181226 67516
rect 186222 66308 186228 66360
rect 186280 66348 186286 66360
rect 186590 66348 186596 66360
rect 186280 66320 186596 66348
rect 186280 66308 186286 66320
rect 186590 66308 186596 66320
rect 186648 66308 186654 66360
rect 339218 66308 339224 66360
rect 339276 66348 339282 66360
rect 339310 66348 339316 66360
rect 339276 66320 339316 66348
rect 339276 66308 339282 66320
rect 339310 66308 339316 66320
rect 339368 66308 339374 66360
rect 138106 66240 138112 66292
rect 138164 66280 138170 66292
rect 138290 66280 138296 66292
rect 138164 66252 138296 66280
rect 138164 66240 138170 66252
rect 138290 66240 138296 66252
rect 138348 66240 138354 66292
rect 144822 66240 144828 66292
rect 144880 66280 144886 66292
rect 145098 66280 145104 66292
rect 144880 66252 145104 66280
rect 144880 66240 144886 66252
rect 145098 66240 145104 66252
rect 145156 66240 145162 66292
rect 162946 66240 162952 66292
rect 163004 66280 163010 66292
rect 163130 66280 163136 66292
rect 163004 66252 163136 66280
rect 163004 66240 163010 66252
rect 163130 66240 163136 66252
rect 163188 66240 163194 66292
rect 219618 66240 219624 66292
rect 219676 66280 219682 66292
rect 219710 66280 219716 66292
rect 219676 66252 219716 66280
rect 219676 66240 219682 66252
rect 219710 66240 219716 66252
rect 219768 66240 219774 66292
rect 244366 66240 244372 66292
rect 244424 66280 244430 66292
rect 244642 66280 244648 66292
rect 244424 66252 244648 66280
rect 244424 66240 244430 66252
rect 244642 66240 244648 66252
rect 244700 66240 244706 66292
rect 251266 66240 251272 66292
rect 251324 66280 251330 66292
rect 251358 66280 251364 66292
rect 251324 66252 251364 66280
rect 251324 66240 251330 66252
rect 251358 66240 251364 66252
rect 251416 66240 251422 66292
rect 403802 66240 403808 66292
rect 403860 66280 403866 66292
rect 404078 66280 404084 66292
rect 403860 66252 404084 66280
rect 403860 66240 403866 66252
rect 404078 66240 404084 66252
rect 404136 66240 404142 66292
rect 143626 66172 143632 66224
rect 143684 66212 143690 66224
rect 143810 66212 143816 66224
rect 143684 66184 143816 66212
rect 143684 66172 143690 66184
rect 143810 66172 143816 66184
rect 143868 66172 143874 66224
rect 186130 66172 186136 66224
rect 186188 66212 186194 66224
rect 186222 66212 186228 66224
rect 186188 66184 186228 66212
rect 186188 66172 186194 66184
rect 186222 66172 186228 66184
rect 186280 66172 186286 66224
rect 220998 66172 221004 66224
rect 221056 66212 221062 66224
rect 221090 66212 221096 66224
rect 221056 66184 221096 66212
rect 221056 66172 221062 66184
rect 221090 66172 221096 66184
rect 221148 66172 221154 66224
rect 249886 66172 249892 66224
rect 249944 66172 249950 66224
rect 409414 66172 409420 66224
rect 409472 66212 409478 66224
rect 409506 66212 409512 66224
rect 409472 66184 409512 66212
rect 409472 66172 409478 66184
rect 409506 66172 409512 66184
rect 409564 66172 409570 66224
rect 414750 66172 414756 66224
rect 414808 66212 414814 66224
rect 414934 66212 414940 66224
rect 414808 66184 414940 66212
rect 414808 66172 414814 66184
rect 414934 66172 414940 66184
rect 414992 66172 414998 66224
rect 249904 66144 249932 66172
rect 250162 66144 250168 66156
rect 249904 66116 250168 66144
rect 250162 66104 250168 66116
rect 250220 66104 250226 66156
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 131574 64852 131580 64864
rect 3384 64824 131580 64852
rect 3384 64812 3390 64824
rect 131574 64812 131580 64824
rect 131632 64812 131638 64864
rect 164510 64812 164516 64864
rect 164568 64852 164574 64864
rect 164786 64852 164792 64864
rect 164568 64824 164792 64852
rect 164568 64812 164574 64824
rect 164786 64812 164792 64824
rect 164844 64812 164850 64864
rect 173802 64812 173808 64864
rect 173860 64852 173866 64864
rect 173986 64852 173992 64864
rect 173860 64824 173992 64852
rect 173860 64812 173866 64824
rect 173986 64812 173992 64824
rect 174044 64812 174050 64864
rect 220998 64812 221004 64864
rect 221056 64852 221062 64864
rect 221182 64852 221188 64864
rect 221056 64824 221188 64852
rect 221056 64812 221062 64824
rect 221182 64812 221188 64824
rect 221240 64812 221246 64864
rect 339126 64812 339132 64864
rect 339184 64852 339190 64864
rect 339494 64852 339500 64864
rect 339184 64824 339500 64852
rect 339184 64812 339190 64824
rect 339494 64812 339500 64824
rect 339552 64812 339558 64864
rect 425974 64812 425980 64864
rect 426032 64852 426038 64864
rect 426066 64852 426072 64864
rect 426032 64824 426072 64852
rect 426032 64812 426038 64824
rect 426066 64812 426072 64824
rect 426124 64812 426130 64864
rect 431402 64812 431408 64864
rect 431460 64852 431466 64864
rect 431586 64852 431592 64864
rect 431460 64824 431592 64852
rect 431460 64812 431466 64824
rect 431586 64812 431592 64824
rect 431644 64812 431650 64864
rect 436830 64812 436836 64864
rect 436888 64852 436894 64864
rect 579798 64852 579804 64864
rect 436888 64824 579804 64852
rect 436888 64812 436894 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 383286 60840 383292 60852
rect 383212 60812 383292 60840
rect 383212 60716 383240 60812
rect 383286 60800 383292 60812
rect 383344 60800 383350 60852
rect 420730 60772 420736 60784
rect 420656 60744 420736 60772
rect 420656 60716 420684 60744
rect 420730 60732 420736 60744
rect 420788 60732 420794 60784
rect 128814 60664 128820 60716
rect 128872 60704 128878 60716
rect 129090 60704 129096 60716
rect 128872 60676 129096 60704
rect 128872 60664 128878 60676
rect 129090 60664 129096 60676
rect 129148 60664 129154 60716
rect 189166 60664 189172 60716
rect 189224 60704 189230 60716
rect 189350 60704 189356 60716
rect 189224 60676 189356 60704
rect 189224 60664 189230 60676
rect 189350 60664 189356 60676
rect 189408 60664 189414 60716
rect 227806 60664 227812 60716
rect 227864 60704 227870 60716
rect 227990 60704 227996 60716
rect 227864 60676 227996 60704
rect 227864 60664 227870 60676
rect 227990 60664 227996 60676
rect 228048 60664 228054 60716
rect 383194 60664 383200 60716
rect 383252 60664 383258 60716
rect 420638 60664 420644 60716
rect 420696 60664 420702 60716
rect 203058 57944 203064 57996
rect 203116 57984 203122 57996
rect 203242 57984 203248 57996
rect 203116 57956 203248 57984
rect 203116 57944 203122 57956
rect 203242 57944 203248 57956
rect 203300 57944 203306 57996
rect 238938 57944 238944 57996
rect 238996 57984 239002 57996
rect 239122 57984 239128 57996
rect 238996 57956 239128 57984
rect 238996 57944 239002 57956
rect 239122 57944 239128 57956
rect 239180 57944 239186 57996
rect 314010 57944 314016 57996
rect 314068 57944 314074 57996
rect 132954 57876 132960 57928
rect 133012 57916 133018 57928
rect 133230 57916 133236 57928
rect 133012 57888 133236 57916
rect 133012 57876 133018 57888
rect 133230 57876 133236 57888
rect 133288 57876 133294 57928
rect 181070 57876 181076 57928
rect 181128 57916 181134 57928
rect 181162 57916 181168 57928
rect 181128 57888 181168 57916
rect 181128 57876 181134 57888
rect 181162 57876 181168 57888
rect 181220 57876 181226 57928
rect 209682 57876 209688 57928
rect 209740 57916 209746 57928
rect 209958 57916 209964 57928
rect 209740 57888 209964 57916
rect 209740 57876 209746 57888
rect 209958 57876 209964 57888
rect 210016 57876 210022 57928
rect 227714 57876 227720 57928
rect 227772 57916 227778 57928
rect 227990 57916 227996 57928
rect 227772 57888 227996 57916
rect 227772 57876 227778 57888
rect 227990 57876 227996 57888
rect 228048 57876 228054 57928
rect 233326 57876 233332 57928
rect 233384 57916 233390 57928
rect 233510 57916 233516 57928
rect 233384 57888 233516 57916
rect 233384 57876 233390 57888
rect 233510 57876 233516 57888
rect 233568 57876 233574 57928
rect 276106 57876 276112 57928
rect 276164 57916 276170 57928
rect 276198 57916 276204 57928
rect 276164 57888 276204 57916
rect 276164 57876 276170 57888
rect 276198 57876 276204 57888
rect 276256 57876 276262 57928
rect 314028 57860 314056 57944
rect 383010 57876 383016 57928
rect 383068 57916 383074 57928
rect 383194 57916 383200 57928
rect 383068 57888 383200 57916
rect 383068 57876 383074 57888
rect 383194 57876 383200 57888
rect 383252 57876 383258 57928
rect 420454 57876 420460 57928
rect 420512 57916 420518 57928
rect 420730 57916 420736 57928
rect 420512 57888 420736 57916
rect 420512 57876 420518 57888
rect 420730 57876 420736 57888
rect 420788 57876 420794 57928
rect 314010 57808 314016 57860
rect 314068 57808 314074 57860
rect 159082 56652 159088 56704
rect 159140 56652 159146 56704
rect 219618 56652 219624 56704
rect 219676 56692 219682 56704
rect 219802 56692 219808 56704
rect 219676 56664 219808 56692
rect 219676 56652 219682 56664
rect 219802 56652 219808 56664
rect 219860 56652 219866 56704
rect 143626 56584 143632 56636
rect 143684 56624 143690 56636
rect 143810 56624 143816 56636
rect 143684 56596 143816 56624
rect 143684 56584 143690 56596
rect 143810 56584 143816 56596
rect 143868 56584 143874 56636
rect 145098 56584 145104 56636
rect 145156 56624 145162 56636
rect 145190 56624 145196 56636
rect 145156 56596 145196 56624
rect 145156 56584 145162 56596
rect 145190 56584 145196 56596
rect 145248 56584 145254 56636
rect 159100 56624 159128 56652
rect 159174 56624 159180 56636
rect 159100 56596 159180 56624
rect 159174 56584 159180 56596
rect 159232 56584 159238 56636
rect 183738 56584 183744 56636
rect 183796 56624 183802 56636
rect 183830 56624 183836 56636
rect 183796 56596 183836 56624
rect 183796 56584 183802 56596
rect 183830 56584 183836 56596
rect 183888 56584 183894 56636
rect 184750 56584 184756 56636
rect 184808 56624 184814 56636
rect 184934 56624 184940 56636
rect 184808 56596 184940 56624
rect 184808 56584 184814 56596
rect 184934 56584 184940 56596
rect 184992 56584 184998 56636
rect 186130 56584 186136 56636
rect 186188 56624 186194 56636
rect 186222 56624 186228 56636
rect 186188 56596 186228 56624
rect 186188 56584 186194 56596
rect 186222 56584 186228 56596
rect 186280 56584 186286 56636
rect 244274 56584 244280 56636
rect 244332 56624 244338 56636
rect 244550 56624 244556 56636
rect 244332 56596 244556 56624
rect 244332 56584 244338 56596
rect 244550 56584 244556 56596
rect 244608 56584 244614 56636
rect 250070 56584 250076 56636
rect 250128 56624 250134 56636
rect 250162 56624 250168 56636
rect 250128 56596 250168 56624
rect 250128 56584 250134 56596
rect 250162 56584 250168 56596
rect 250220 56584 250226 56636
rect 253658 56584 253664 56636
rect 253716 56624 253722 56636
rect 253750 56624 253756 56636
rect 253716 56596 253756 56624
rect 253716 56584 253722 56596
rect 253750 56584 253756 56596
rect 253808 56584 253814 56636
rect 400766 56584 400772 56636
rect 400824 56624 400830 56636
rect 400950 56624 400956 56636
rect 400824 56596 400956 56624
rect 400824 56584 400830 56596
rect 400950 56584 400956 56596
rect 401008 56584 401014 56636
rect 409322 56584 409328 56636
rect 409380 56624 409386 56636
rect 409414 56624 409420 56636
rect 409380 56596 409420 56624
rect 409380 56584 409386 56596
rect 409414 56584 409420 56596
rect 409472 56584 409478 56636
rect 414750 56584 414756 56636
rect 414808 56624 414814 56636
rect 415210 56624 415216 56636
rect 414808 56596 415216 56624
rect 414808 56584 414814 56596
rect 415210 56584 415216 56596
rect 415268 56584 415274 56636
rect 162946 56516 162952 56568
rect 163004 56556 163010 56568
rect 163130 56556 163136 56568
rect 163004 56528 163136 56556
rect 163004 56516 163010 56528
rect 163130 56516 163136 56528
rect 163188 56516 163194 56568
rect 179506 56516 179512 56568
rect 179564 56556 179570 56568
rect 179598 56556 179604 56568
rect 179564 56528 179604 56556
rect 179564 56516 179570 56528
rect 179598 56516 179604 56528
rect 179656 56516 179662 56568
rect 180978 56516 180984 56568
rect 181036 56556 181042 56568
rect 181070 56556 181076 56568
rect 181036 56528 181076 56556
rect 181036 56516 181042 56528
rect 181070 56516 181076 56528
rect 181128 56516 181134 56568
rect 218146 56516 218152 56568
rect 218204 56556 218210 56568
rect 218238 56556 218244 56568
rect 218204 56528 218244 56556
rect 218204 56516 218210 56528
rect 218238 56516 218244 56528
rect 218296 56516 218302 56568
rect 403802 56516 403808 56568
rect 403860 56556 403866 56568
rect 403986 56556 403992 56568
rect 403860 56528 403992 56556
rect 403860 56516 403866 56528
rect 403986 56516 403992 56528
rect 404044 56516 404050 56568
rect 425974 55292 425980 55344
rect 426032 55332 426038 55344
rect 426066 55332 426072 55344
rect 426032 55304 426072 55332
rect 426032 55292 426038 55304
rect 426066 55292 426072 55304
rect 426124 55292 426130 55344
rect 173802 55224 173808 55276
rect 173860 55264 173866 55276
rect 174078 55264 174084 55276
rect 173860 55236 174084 55264
rect 173860 55224 173866 55236
rect 174078 55224 174084 55236
rect 174136 55224 174142 55276
rect 220998 55224 221004 55276
rect 221056 55264 221062 55276
rect 221182 55264 221188 55276
rect 221056 55236 221188 55264
rect 221056 55224 221062 55236
rect 221182 55224 221188 55236
rect 221240 55224 221246 55276
rect 431402 55224 431408 55276
rect 431460 55264 431466 55276
rect 431586 55264 431592 55276
rect 431460 55236 431592 55264
rect 431460 55224 431466 55236
rect 431586 55224 431592 55236
rect 431644 55224 431650 55276
rect 425790 55156 425796 55208
rect 425848 55196 425854 55208
rect 426066 55196 426072 55208
rect 425848 55168 426072 55196
rect 425848 55156 425854 55168
rect 426066 55156 426072 55168
rect 426124 55156 426130 55208
rect 274726 53116 274732 53168
rect 274784 53156 274790 53168
rect 275094 53156 275100 53168
rect 274784 53128 275100 53156
rect 274784 53116 274790 53128
rect 275094 53116 275100 53128
rect 275152 53116 275158 53168
rect 145190 51116 145196 51128
rect 145116 51088 145196 51116
rect 145116 51060 145144 51088
rect 145190 51076 145196 51088
rect 145248 51076 145254 51128
rect 189350 51076 189356 51128
rect 189408 51076 189414 51128
rect 314010 51076 314016 51128
rect 314068 51076 314074 51128
rect 145098 51008 145104 51060
rect 145156 51008 145162 51060
rect 189368 50992 189396 51076
rect 196066 51008 196072 51060
rect 196124 51008 196130 51060
rect 189350 50940 189356 50992
rect 189408 50940 189414 50992
rect 196084 50980 196112 51008
rect 314028 50992 314056 51076
rect 409322 51008 409328 51060
rect 409380 51048 409386 51060
rect 409506 51048 409512 51060
rect 409380 51020 409512 51048
rect 409380 51008 409386 51020
rect 409506 51008 409512 51020
rect 409564 51008 409570 51060
rect 196158 50980 196164 50992
rect 196084 50952 196164 50980
rect 196158 50940 196164 50952
rect 196216 50940 196222 50992
rect 314010 50940 314016 50992
rect 314068 50940 314074 50992
rect 253658 48356 253664 48408
rect 253716 48396 253722 48408
rect 253750 48396 253756 48408
rect 253716 48368 253756 48396
rect 253716 48356 253722 48368
rect 253750 48356 253756 48368
rect 253808 48356 253814 48408
rect 276106 48356 276112 48408
rect 276164 48396 276170 48408
rect 276198 48396 276204 48408
rect 276164 48368 276204 48396
rect 276164 48356 276170 48368
rect 276198 48356 276204 48368
rect 276256 48356 276262 48408
rect 129090 48328 129096 48340
rect 129016 48300 129096 48328
rect 129016 48272 129044 48300
rect 129090 48288 129096 48300
rect 129148 48288 129154 48340
rect 159082 48288 159088 48340
rect 159140 48288 159146 48340
rect 161566 48288 161572 48340
rect 161624 48328 161630 48340
rect 161750 48328 161756 48340
rect 161624 48300 161756 48328
rect 161624 48288 161630 48300
rect 161750 48288 161756 48300
rect 161808 48288 161814 48340
rect 227714 48288 227720 48340
rect 227772 48328 227778 48340
rect 227898 48328 227904 48340
rect 227772 48300 227904 48328
rect 227772 48288 227778 48300
rect 227898 48288 227904 48300
rect 227956 48288 227962 48340
rect 233326 48288 233332 48340
rect 233384 48328 233390 48340
rect 233602 48328 233608 48340
rect 233384 48300 233608 48328
rect 233384 48288 233390 48300
rect 233602 48288 233608 48300
rect 233660 48288 233666 48340
rect 274910 48288 274916 48340
rect 274968 48328 274974 48340
rect 275094 48328 275100 48340
rect 274968 48300 275100 48328
rect 274968 48288 274974 48300
rect 275094 48288 275100 48300
rect 275152 48288 275158 48340
rect 317138 48288 317144 48340
rect 317196 48328 317202 48340
rect 317230 48328 317236 48340
rect 317196 48300 317236 48328
rect 317196 48288 317202 48300
rect 317230 48288 317236 48300
rect 317288 48288 317294 48340
rect 383010 48288 383016 48340
rect 383068 48328 383074 48340
rect 383286 48328 383292 48340
rect 383068 48300 383292 48328
rect 383068 48288 383074 48300
rect 383286 48288 383292 48300
rect 383344 48288 383350 48340
rect 414934 48288 414940 48340
rect 414992 48328 414998 48340
rect 415210 48328 415216 48340
rect 414992 48300 415216 48328
rect 414992 48288 414998 48300
rect 415210 48288 415216 48300
rect 415268 48288 415274 48340
rect 128998 48220 129004 48272
rect 129056 48220 129062 48272
rect 159100 48260 159128 48288
rect 159174 48260 159180 48272
rect 159100 48232 159180 48260
rect 159174 48220 159180 48232
rect 159232 48220 159238 48272
rect 238754 48220 238760 48272
rect 238812 48260 238818 48272
rect 238938 48260 238944 48272
rect 238812 48232 238944 48260
rect 238812 48220 238818 48232
rect 238938 48220 238944 48232
rect 238996 48220 239002 48272
rect 420546 48220 420552 48272
rect 420604 48260 420610 48272
rect 420638 48260 420644 48272
rect 420604 48232 420644 48260
rect 420604 48220 420610 48232
rect 420638 48220 420644 48232
rect 420696 48220 420702 48272
rect 158990 46928 158996 46980
rect 159048 46968 159054 46980
rect 159174 46968 159180 46980
rect 159048 46940 159180 46968
rect 159048 46928 159054 46940
rect 159174 46928 159180 46940
rect 159232 46928 159238 46980
rect 162946 46928 162952 46980
rect 163004 46968 163010 46980
rect 163130 46968 163136 46980
rect 163004 46940 163136 46968
rect 163004 46928 163010 46940
rect 163130 46928 163136 46940
rect 163188 46928 163194 46980
rect 164602 46928 164608 46980
rect 164660 46968 164666 46980
rect 164786 46968 164792 46980
rect 164660 46940 164792 46968
rect 164660 46928 164666 46940
rect 164786 46928 164792 46940
rect 164844 46928 164850 46980
rect 168466 46928 168472 46980
rect 168524 46968 168530 46980
rect 168558 46968 168564 46980
rect 168524 46940 168564 46968
rect 168524 46928 168530 46940
rect 168558 46928 168564 46940
rect 168616 46928 168622 46980
rect 173894 46928 173900 46980
rect 173952 46968 173958 46980
rect 174078 46968 174084 46980
rect 173952 46940 174084 46968
rect 173952 46928 173958 46940
rect 174078 46928 174084 46940
rect 174136 46928 174142 46980
rect 179506 46928 179512 46980
rect 179564 46968 179570 46980
rect 179690 46968 179696 46980
rect 179564 46940 179696 46968
rect 179564 46928 179570 46940
rect 179690 46928 179696 46940
rect 179748 46928 179754 46980
rect 180978 46928 180984 46980
rect 181036 46968 181042 46980
rect 181162 46968 181168 46980
rect 181036 46940 181168 46968
rect 181036 46928 181042 46940
rect 181162 46928 181168 46940
rect 181220 46928 181226 46980
rect 218146 46928 218152 46980
rect 218204 46968 218210 46980
rect 218422 46968 218428 46980
rect 218204 46940 218428 46968
rect 218204 46928 218210 46940
rect 218422 46928 218428 46940
rect 218480 46928 218486 46980
rect 341242 46928 341248 46980
rect 341300 46968 341306 46980
rect 341334 46968 341340 46980
rect 341300 46940 341340 46968
rect 341300 46928 341306 46940
rect 341334 46928 341340 46940
rect 341392 46928 341398 46980
rect 403802 46928 403808 46980
rect 403860 46968 403866 46980
rect 404078 46968 404084 46980
rect 403860 46940 404084 46968
rect 403860 46928 403866 46940
rect 404078 46928 404084 46940
rect 404136 46928 404142 46980
rect 129090 46860 129096 46912
rect 129148 46860 129154 46912
rect 253474 46860 253480 46912
rect 253532 46900 253538 46912
rect 253750 46900 253756 46912
rect 253532 46872 253756 46900
rect 253532 46860 253538 46872
rect 253750 46860 253756 46872
rect 253808 46860 253814 46912
rect 276106 46860 276112 46912
rect 276164 46900 276170 46912
rect 276198 46900 276204 46912
rect 276164 46872 276204 46900
rect 276164 46860 276170 46872
rect 276198 46860 276204 46872
rect 276256 46860 276262 46912
rect 129108 46776 129136 46860
rect 341242 46792 341248 46844
rect 341300 46832 341306 46844
rect 341426 46832 341432 46844
rect 341300 46804 341432 46832
rect 341300 46792 341306 46804
rect 341426 46792 341432 46804
rect 341484 46792 341490 46844
rect 129090 46724 129096 46776
rect 129148 46724 129154 46776
rect 339218 45568 339224 45620
rect 339276 45608 339282 45620
rect 339494 45608 339500 45620
rect 339276 45580 339500 45608
rect 339276 45568 339282 45580
rect 339494 45568 339500 45580
rect 339552 45568 339558 45620
rect 425790 45568 425796 45620
rect 425848 45608 425854 45620
rect 425974 45608 425980 45620
rect 425848 45580 425980 45608
rect 425848 45568 425854 45580
rect 425974 45568 425980 45580
rect 426032 45568 426038 45620
rect 173710 45500 173716 45552
rect 173768 45540 173774 45552
rect 173894 45540 173900 45552
rect 173768 45512 173900 45540
rect 173768 45500 173774 45512
rect 173894 45500 173900 45512
rect 173952 45500 173958 45552
rect 179414 45500 179420 45552
rect 179472 45540 179478 45552
rect 179690 45540 179696 45552
rect 179472 45512 179696 45540
rect 179472 45500 179478 45512
rect 179690 45500 179696 45512
rect 179748 45500 179754 45552
rect 219710 45500 219716 45552
rect 219768 45540 219774 45552
rect 219894 45540 219900 45552
rect 219768 45512 219900 45540
rect 219768 45500 219774 45512
rect 219894 45500 219900 45512
rect 219952 45500 219958 45552
rect 220998 45500 221004 45552
rect 221056 45540 221062 45552
rect 221274 45540 221280 45552
rect 221056 45512 221280 45540
rect 221056 45500 221062 45512
rect 221274 45500 221280 45512
rect 221332 45500 221338 45552
rect 431494 45500 431500 45552
rect 431552 45540 431558 45552
rect 431586 45540 431592 45552
rect 431552 45512 431592 45540
rect 431552 45500 431558 45512
rect 431586 45500 431592 45512
rect 431644 45500 431650 45552
rect 425790 45432 425796 45484
rect 425848 45472 425854 45484
rect 425974 45472 425980 45484
rect 425848 45444 425980 45472
rect 425848 45432 425854 45444
rect 425974 45432 425980 45444
rect 426032 45432 426038 45484
rect 313734 43460 313740 43512
rect 313792 43500 313798 43512
rect 314010 43500 314016 43512
rect 313792 43472 314016 43500
rect 313792 43460 313798 43472
rect 314010 43460 314016 43472
rect 314068 43460 314074 43512
rect 227898 41556 227904 41608
rect 227956 41556 227962 41608
rect 227916 41472 227944 41556
rect 183572 41432 183876 41460
rect 132034 41352 132040 41404
rect 132092 41392 132098 41404
rect 183572 41392 183600 41432
rect 132092 41364 183600 41392
rect 183848 41392 183876 41432
rect 227898 41420 227904 41472
rect 227956 41420 227962 41472
rect 580166 41392 580172 41404
rect 183848 41364 580172 41392
rect 132092 41352 132098 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 157334 38632 157340 38684
rect 157392 38672 157398 38684
rect 157426 38672 157432 38684
rect 157392 38644 157432 38672
rect 157392 38632 157398 38644
rect 157426 38632 157432 38644
rect 157484 38632 157490 38684
rect 161566 38632 161572 38684
rect 161624 38672 161630 38684
rect 161658 38672 161664 38684
rect 161624 38644 161664 38672
rect 161624 38632 161630 38644
rect 161658 38632 161664 38644
rect 161716 38632 161722 38684
rect 189074 38632 189080 38684
rect 189132 38672 189138 38684
rect 189350 38672 189356 38684
rect 189132 38644 189356 38672
rect 189132 38632 189138 38644
rect 189350 38632 189356 38644
rect 189408 38632 189414 38684
rect 233234 38632 233240 38684
rect 233292 38672 233298 38684
rect 233602 38672 233608 38684
rect 233292 38644 233608 38672
rect 233292 38632 233298 38644
rect 233602 38632 233608 38644
rect 233660 38632 233666 38684
rect 244274 38632 244280 38684
rect 244332 38672 244338 38684
rect 244550 38672 244556 38684
rect 244332 38644 244556 38672
rect 244332 38632 244338 38644
rect 244550 38632 244556 38644
rect 244608 38632 244614 38684
rect 249794 38632 249800 38684
rect 249852 38672 249858 38684
rect 250070 38672 250076 38684
rect 249852 38644 250076 38672
rect 249852 38632 249858 38644
rect 250070 38632 250076 38644
rect 250128 38632 250134 38684
rect 313734 38632 313740 38684
rect 313792 38672 313798 38684
rect 313918 38672 313924 38684
rect 313792 38644 313924 38672
rect 313792 38632 313798 38644
rect 313918 38632 313924 38644
rect 313976 38632 313982 38684
rect 132954 38564 132960 38616
rect 133012 38604 133018 38616
rect 133230 38604 133236 38616
rect 133012 38576 133236 38604
rect 133012 38564 133018 38576
rect 133230 38564 133236 38576
rect 133288 38564 133294 38616
rect 168374 38564 168380 38616
rect 168432 38604 168438 38616
rect 168558 38604 168564 38616
rect 168432 38576 168564 38604
rect 168432 38564 168438 38576
rect 168558 38564 168564 38576
rect 168616 38564 168622 38616
rect 184934 38564 184940 38616
rect 184992 38604 184998 38616
rect 185026 38604 185032 38616
rect 184992 38576 185032 38604
rect 184992 38564 184998 38576
rect 185026 38564 185032 38576
rect 185084 38564 185090 38616
rect 251174 38564 251180 38616
rect 251232 38604 251238 38616
rect 251358 38604 251364 38616
rect 251232 38576 251364 38604
rect 251232 38564 251238 38576
rect 251358 38564 251364 38576
rect 251416 38564 251422 38616
rect 274726 38564 274732 38616
rect 274784 38604 274790 38616
rect 275094 38604 275100 38616
rect 274784 38576 275100 38604
rect 274784 38564 274790 38576
rect 275094 38564 275100 38576
rect 275152 38564 275158 38616
rect 383010 38564 383016 38616
rect 383068 38604 383074 38616
rect 383194 38604 383200 38616
rect 383068 38576 383200 38604
rect 383068 38564 383074 38576
rect 383194 38564 383200 38576
rect 383252 38564 383258 38616
rect 400582 38564 400588 38616
rect 400640 38604 400646 38616
rect 400766 38604 400772 38616
rect 400640 38576 400772 38604
rect 400640 38564 400646 38576
rect 400766 38564 400772 38576
rect 400824 38564 400830 38616
rect 409322 38564 409328 38616
rect 409380 38604 409386 38616
rect 409598 38604 409604 38616
rect 409380 38576 409604 38604
rect 409380 38564 409386 38576
rect 409598 38564 409604 38576
rect 409656 38564 409662 38616
rect 339218 37380 339224 37392
rect 339144 37352 339224 37380
rect 253474 37272 253480 37324
rect 253532 37312 253538 37324
rect 253566 37312 253572 37324
rect 253532 37284 253572 37312
rect 253532 37272 253538 37284
rect 253566 37272 253572 37284
rect 253624 37272 253630 37324
rect 339144 37256 339172 37352
rect 339218 37340 339224 37352
rect 339276 37340 339282 37392
rect 158714 37204 158720 37256
rect 158772 37244 158778 37256
rect 158990 37244 158996 37256
rect 158772 37216 158996 37244
rect 158772 37204 158778 37216
rect 158990 37204 158996 37216
rect 159048 37204 159054 37256
rect 244090 37204 244096 37256
rect 244148 37244 244154 37256
rect 244274 37244 244280 37256
rect 244148 37216 244280 37244
rect 244148 37204 244154 37216
rect 244274 37204 244280 37216
rect 244332 37204 244338 37256
rect 249794 37204 249800 37256
rect 249852 37244 249858 37256
rect 250162 37244 250168 37256
rect 249852 37216 250168 37244
rect 249852 37204 249858 37216
rect 250162 37204 250168 37216
rect 250220 37204 250226 37256
rect 339126 37204 339132 37256
rect 339184 37204 339190 37256
rect 173710 35912 173716 35964
rect 173768 35952 173774 35964
rect 173986 35952 173992 35964
rect 173768 35924 173992 35952
rect 173768 35912 173774 35924
rect 173986 35912 173992 35924
rect 174044 35912 174050 35964
rect 179414 35912 179420 35964
rect 179472 35952 179478 35964
rect 179598 35952 179604 35964
rect 179472 35924 179604 35952
rect 179472 35912 179478 35924
rect 179598 35912 179604 35924
rect 179656 35912 179662 35964
rect 219710 35912 219716 35964
rect 219768 35952 219774 35964
rect 219986 35952 219992 35964
rect 219768 35924 219992 35952
rect 219768 35912 219774 35924
rect 219986 35912 219992 35924
rect 220044 35912 220050 35964
rect 431402 35912 431408 35964
rect 431460 35952 431466 35964
rect 431494 35952 431500 35964
rect 431460 35924 431500 35952
rect 431460 35912 431466 35924
rect 431494 35912 431500 35924
rect 431552 35912 431558 35964
rect 3418 35844 3424 35896
rect 3476 35884 3482 35896
rect 436278 35884 436284 35896
rect 3476 35856 436284 35884
rect 3476 35844 3482 35856
rect 436278 35844 436284 35856
rect 436336 35844 436342 35896
rect 143810 34484 143816 34536
rect 143868 34524 143874 34536
rect 143994 34524 144000 34536
rect 143868 34496 144000 34524
rect 143868 34484 143874 34496
rect 143994 34484 144000 34496
rect 144052 34484 144058 34536
rect 425974 34484 425980 34536
rect 426032 34524 426038 34536
rect 426066 34524 426072 34536
rect 426032 34496 426072 34524
rect 426032 34484 426038 34496
rect 426066 34484 426072 34496
rect 426124 34484 426130 34536
rect 128814 33804 128820 33856
rect 128872 33844 128878 33856
rect 129090 33844 129096 33856
rect 128872 33816 129096 33844
rect 128872 33804 128878 33816
rect 129090 33804 129096 33816
rect 129148 33804 129154 33856
rect 420454 33804 420460 33856
rect 420512 33844 420518 33856
rect 420638 33844 420644 33856
rect 420512 33816 420644 33844
rect 420512 33804 420518 33816
rect 420638 33804 420644 33816
rect 420696 33804 420702 33856
rect 138106 31832 138112 31884
rect 138164 31872 138170 31884
rect 138290 31872 138296 31884
rect 138164 31844 138296 31872
rect 138164 31832 138170 31844
rect 138290 31832 138296 31844
rect 138348 31832 138354 31884
rect 227898 31764 227904 31816
rect 227956 31764 227962 31816
rect 251174 31764 251180 31816
rect 251232 31804 251238 31816
rect 251232 31776 251312 31804
rect 251232 31764 251238 31776
rect 190638 31696 190644 31748
rect 190696 31736 190702 31748
rect 190822 31736 190828 31748
rect 190696 31708 190828 31736
rect 190696 31696 190702 31708
rect 190822 31696 190828 31708
rect 190880 31696 190886 31748
rect 227916 31680 227944 31764
rect 251284 31748 251312 31776
rect 404078 31764 404084 31816
rect 404136 31764 404142 31816
rect 415118 31764 415124 31816
rect 415176 31764 415182 31816
rect 251266 31696 251272 31748
rect 251324 31696 251330 31748
rect 404096 31680 404124 31764
rect 415026 31696 415032 31748
rect 415084 31736 415090 31748
rect 415136 31736 415164 31764
rect 415084 31708 415164 31736
rect 415084 31696 415090 31708
rect 227898 31628 227904 31680
rect 227956 31628 227962 31680
rect 404078 31628 404084 31680
rect 404136 31628 404142 31680
rect 132126 30268 132132 30320
rect 132184 30308 132190 30320
rect 580166 30308 580172 30320
rect 132184 30280 580172 30308
rect 132184 30268 132190 30280
rect 580166 30268 580172 30280
rect 580224 30268 580230 30320
rect 161658 29084 161664 29096
rect 161584 29056 161664 29084
rect 161584 29028 161612 29056
rect 161658 29044 161664 29056
rect 161716 29044 161722 29096
rect 219986 29084 219992 29096
rect 219820 29056 219992 29084
rect 161566 28976 161572 29028
rect 161624 28976 161630 29028
rect 209590 28976 209596 29028
rect 209648 29016 209654 29028
rect 209958 29016 209964 29028
rect 209648 28988 209964 29016
rect 209648 28976 209654 28988
rect 209958 28976 209964 28988
rect 210016 28976 210022 29028
rect 218238 28976 218244 29028
rect 218296 29016 218302 29028
rect 218422 29016 218428 29028
rect 218296 28988 218428 29016
rect 218296 28976 218302 28988
rect 218422 28976 218428 28988
rect 218480 28976 218486 29028
rect 219820 28960 219848 29056
rect 219986 29044 219992 29056
rect 220044 29044 220050 29096
rect 253566 29044 253572 29096
rect 253624 29084 253630 29096
rect 253750 29084 253756 29096
rect 253624 29056 253756 29084
rect 253624 29044 253630 29056
rect 253750 29044 253756 29056
rect 253808 29044 253814 29096
rect 276106 29044 276112 29096
rect 276164 29084 276170 29096
rect 276198 29084 276204 29096
rect 276164 29056 276204 29084
rect 276164 29044 276170 29056
rect 276198 29044 276204 29056
rect 276256 29044 276262 29096
rect 227806 28976 227812 29028
rect 227864 29016 227870 29028
rect 227898 29016 227904 29028
rect 227864 28988 227904 29016
rect 227864 28976 227870 28988
rect 227898 28976 227904 28988
rect 227956 28976 227962 29028
rect 274910 28976 274916 29028
rect 274968 29016 274974 29028
rect 275094 29016 275100 29028
rect 274968 28988 275100 29016
rect 274968 28976 274974 28988
rect 275094 28976 275100 28988
rect 275152 28976 275158 29028
rect 317138 28976 317144 29028
rect 317196 29016 317202 29028
rect 317230 29016 317236 29028
rect 317196 28988 317236 29016
rect 317196 28976 317202 28988
rect 317230 28976 317236 28988
rect 317288 28976 317294 29028
rect 383010 28976 383016 29028
rect 383068 29016 383074 29028
rect 383286 29016 383292 29028
rect 383068 28988 383292 29016
rect 383068 28976 383074 28988
rect 383286 28976 383292 28988
rect 383344 28976 383350 29028
rect 400582 28976 400588 29028
rect 400640 29016 400646 29028
rect 400858 29016 400864 29028
rect 400640 28988 400864 29016
rect 400640 28976 400646 28988
rect 400858 28976 400864 28988
rect 400916 28976 400922 29028
rect 409322 28976 409328 29028
rect 409380 29016 409386 29028
rect 409414 29016 409420 29028
rect 409380 28988 409420 29016
rect 409380 28976 409386 28988
rect 409414 28976 409420 28988
rect 409472 28976 409478 29028
rect 415026 28976 415032 29028
rect 415084 29016 415090 29028
rect 415210 29016 415216 29028
rect 415084 28988 415216 29016
rect 415084 28976 415090 28988
rect 415210 28976 415216 28988
rect 415268 28976 415274 29028
rect 150526 28908 150532 28960
rect 150584 28948 150590 28960
rect 150618 28948 150624 28960
rect 150584 28920 150624 28948
rect 150584 28908 150590 28920
rect 150618 28908 150624 28920
rect 150676 28908 150682 28960
rect 151814 28908 151820 28960
rect 151872 28948 151878 28960
rect 151906 28948 151912 28960
rect 151872 28920 151912 28948
rect 151872 28908 151878 28920
rect 151906 28908 151912 28920
rect 151964 28908 151970 28960
rect 156046 28908 156052 28960
rect 156104 28948 156110 28960
rect 156138 28948 156144 28960
rect 156104 28920 156144 28948
rect 156104 28908 156110 28920
rect 156138 28908 156144 28920
rect 156196 28908 156202 28960
rect 157334 28908 157340 28960
rect 157392 28948 157398 28960
rect 157426 28948 157432 28960
rect 157392 28920 157432 28948
rect 157392 28908 157398 28920
rect 157426 28908 157432 28920
rect 157484 28908 157490 28960
rect 168466 28908 168472 28960
rect 168524 28948 168530 28960
rect 168650 28948 168656 28960
rect 168524 28920 168656 28948
rect 168524 28908 168530 28920
rect 168650 28908 168656 28920
rect 168708 28908 168714 28960
rect 173986 28908 173992 28960
rect 174044 28908 174050 28960
rect 179598 28908 179604 28960
rect 179656 28948 179662 28960
rect 179690 28948 179696 28960
rect 179656 28920 179696 28948
rect 179656 28908 179662 28920
rect 179690 28908 179696 28920
rect 179748 28908 179754 28960
rect 204346 28908 204352 28960
rect 204404 28948 204410 28960
rect 204530 28948 204536 28960
rect 204404 28920 204536 28948
rect 204404 28908 204410 28920
rect 204530 28908 204536 28920
rect 204588 28908 204594 28960
rect 219802 28908 219808 28960
rect 219860 28908 219866 28960
rect 420546 28908 420552 28960
rect 420604 28948 420610 28960
rect 420638 28948 420644 28960
rect 420604 28920 420644 28948
rect 420604 28908 420610 28920
rect 420638 28908 420644 28920
rect 420696 28908 420702 28960
rect 174004 28824 174032 28908
rect 233326 28840 233332 28892
rect 233384 28880 233390 28892
rect 233510 28880 233516 28892
rect 233384 28852 233516 28880
rect 233384 28840 233390 28852
rect 233510 28840 233516 28852
rect 233568 28840 233574 28892
rect 313642 28840 313648 28892
rect 313700 28880 313706 28892
rect 313918 28880 313924 28892
rect 313700 28852 313924 28880
rect 313700 28840 313706 28852
rect 313918 28840 313924 28852
rect 313976 28840 313982 28892
rect 173986 28772 173992 28824
rect 174044 28772 174050 28824
rect 158714 27616 158720 27668
rect 158772 27656 158778 27668
rect 158990 27656 158996 27668
rect 158772 27628 158996 27656
rect 158772 27616 158778 27628
rect 158990 27616 158996 27628
rect 159048 27616 159054 27668
rect 183370 27616 183376 27668
rect 183428 27656 183434 27668
rect 183830 27656 183836 27668
rect 183428 27628 183836 27656
rect 183428 27616 183434 27628
rect 183830 27616 183836 27628
rect 183888 27616 183894 27668
rect 221090 27616 221096 27668
rect 221148 27656 221154 27668
rect 221274 27656 221280 27668
rect 221148 27628 221280 27656
rect 221148 27616 221154 27628
rect 221274 27616 221280 27628
rect 221332 27616 221338 27668
rect 244090 27616 244096 27668
rect 244148 27656 244154 27668
rect 244366 27656 244372 27668
rect 244148 27628 244372 27656
rect 244148 27616 244154 27628
rect 244366 27616 244372 27628
rect 244424 27616 244430 27668
rect 249886 27616 249892 27668
rect 249944 27656 249950 27668
rect 250162 27656 250168 27668
rect 249944 27628 250168 27656
rect 249944 27616 249950 27628
rect 250162 27616 250168 27628
rect 250220 27616 250226 27668
rect 431402 27616 431408 27668
rect 431460 27656 431466 27668
rect 431678 27656 431684 27668
rect 431460 27628 431684 27656
rect 431460 27616 431466 27628
rect 431678 27616 431684 27628
rect 431736 27616 431742 27668
rect 180702 27548 180708 27600
rect 180760 27588 180766 27600
rect 181162 27588 181168 27600
rect 180760 27560 181168 27588
rect 180760 27548 180766 27560
rect 181162 27548 181168 27560
rect 181220 27548 181226 27600
rect 253566 27548 253572 27600
rect 253624 27588 253630 27600
rect 253750 27588 253756 27600
rect 253624 27560 253756 27588
rect 253624 27548 253630 27560
rect 253750 27548 253756 27560
rect 253808 27548 253814 27600
rect 275922 27548 275928 27600
rect 275980 27588 275986 27600
rect 276106 27588 276112 27600
rect 275980 27560 276112 27588
rect 275980 27548 275986 27560
rect 276106 27548 276112 27560
rect 276164 27548 276170 27600
rect 138106 26256 138112 26308
rect 138164 26296 138170 26308
rect 138290 26296 138296 26308
rect 138164 26268 138296 26296
rect 138164 26256 138170 26268
rect 138290 26256 138296 26268
rect 138348 26256 138354 26308
rect 426066 24760 426072 24812
rect 426124 24800 426130 24812
rect 426158 24800 426164 24812
rect 426124 24772 426164 24800
rect 426124 24760 426130 24772
rect 426158 24760 426164 24772
rect 426216 24760 426222 24812
rect 238938 24148 238944 24200
rect 238996 24188 239002 24200
rect 239122 24188 239128 24200
rect 238996 24160 239128 24188
rect 238996 24148 239002 24160
rect 239122 24148 239128 24160
rect 239180 24148 239186 24200
rect 238018 22040 238024 22092
rect 238076 22040 238082 22092
rect 244366 22040 244372 22092
rect 244424 22080 244430 22092
rect 244550 22080 244556 22092
rect 244424 22052 244556 22080
rect 244424 22040 244430 22052
rect 244550 22040 244556 22052
rect 244608 22040 244614 22092
rect 249886 22040 249892 22092
rect 249944 22080 249950 22092
rect 250070 22080 250076 22092
rect 249944 22052 250076 22080
rect 249944 22040 249950 22052
rect 250070 22040 250076 22052
rect 250128 22040 250134 22092
rect 341518 22040 341524 22092
rect 341576 22080 341582 22092
rect 341702 22080 341708 22092
rect 341576 22052 341708 22080
rect 341576 22040 341582 22052
rect 341702 22040 341708 22052
rect 341760 22040 341766 22092
rect 238036 22012 238064 22040
rect 238110 22012 238116 22024
rect 238036 21984 238116 22012
rect 238110 21972 238116 21984
rect 238168 21972 238174 22024
rect 2774 21428 2780 21480
rect 2832 21468 2838 21480
rect 4798 21468 4804 21480
rect 2832 21440 4804 21468
rect 2832 21428 2838 21440
rect 4798 21428 4804 21440
rect 4856 21428 4862 21480
rect 143718 19320 143724 19372
rect 143776 19360 143782 19372
rect 143810 19360 143816 19372
rect 143776 19332 143816 19360
rect 143776 19320 143782 19332
rect 143810 19320 143816 19332
rect 143868 19320 143874 19372
rect 157334 19320 157340 19372
rect 157392 19360 157398 19372
rect 157426 19360 157432 19372
rect 157392 19332 157432 19360
rect 157392 19320 157398 19332
rect 157426 19320 157432 19332
rect 157484 19320 157490 19372
rect 161566 19320 161572 19372
rect 161624 19360 161630 19372
rect 161658 19360 161664 19372
rect 161624 19332 161664 19360
rect 161624 19320 161630 19332
rect 161658 19320 161664 19332
rect 161716 19320 161722 19372
rect 162946 19320 162952 19372
rect 163004 19360 163010 19372
rect 163004 19332 163084 19360
rect 163004 19320 163010 19332
rect 163056 19304 163084 19332
rect 204346 19320 204352 19372
rect 204404 19360 204410 19372
rect 204438 19360 204444 19372
rect 204404 19332 204444 19360
rect 204404 19320 204410 19332
rect 204438 19320 204444 19332
rect 204496 19320 204502 19372
rect 209590 19320 209596 19372
rect 209648 19360 209654 19372
rect 209774 19360 209780 19372
rect 209648 19332 209780 19360
rect 209648 19320 209654 19332
rect 209774 19320 209780 19332
rect 209832 19320 209838 19372
rect 238938 19320 238944 19372
rect 238996 19360 239002 19372
rect 239122 19360 239128 19372
rect 238996 19332 239128 19360
rect 238996 19320 239002 19332
rect 239122 19320 239128 19332
rect 239180 19320 239186 19372
rect 313642 19320 313648 19372
rect 313700 19360 313706 19372
rect 313918 19360 313924 19372
rect 313700 19332 313924 19360
rect 313700 19320 313706 19332
rect 313918 19320 313924 19332
rect 313976 19320 313982 19372
rect 409414 19320 409420 19372
rect 409472 19360 409478 19372
rect 409598 19360 409604 19372
rect 409472 19332 409604 19360
rect 409472 19320 409478 19332
rect 409598 19320 409604 19332
rect 409656 19320 409662 19372
rect 128722 19252 128728 19304
rect 128780 19292 128786 19304
rect 129090 19292 129096 19304
rect 128780 19264 129096 19292
rect 128780 19252 128786 19264
rect 129090 19252 129096 19264
rect 129148 19252 129154 19304
rect 140866 19252 140872 19304
rect 140924 19252 140930 19304
rect 145006 19252 145012 19304
rect 145064 19292 145070 19304
rect 145190 19292 145196 19304
rect 145064 19264 145196 19292
rect 145064 19252 145070 19264
rect 145190 19252 145196 19264
rect 145248 19252 145254 19304
rect 163038 19252 163044 19304
rect 163096 19252 163102 19304
rect 168190 19252 168196 19304
rect 168248 19292 168254 19304
rect 168374 19292 168380 19304
rect 168248 19264 168380 19292
rect 168248 19252 168254 19264
rect 168374 19252 168380 19264
rect 168432 19252 168438 19304
rect 173986 19252 173992 19304
rect 174044 19292 174050 19304
rect 174170 19292 174176 19304
rect 174044 19264 174176 19292
rect 174044 19252 174050 19264
rect 174170 19252 174176 19264
rect 174228 19252 174234 19304
rect 183738 19252 183744 19304
rect 183796 19292 183802 19304
rect 183922 19292 183928 19304
rect 183796 19264 183928 19292
rect 183796 19252 183802 19264
rect 183922 19252 183928 19264
rect 183980 19252 183986 19304
rect 400766 19252 400772 19304
rect 400824 19292 400830 19304
rect 401042 19292 401048 19304
rect 400824 19264 401048 19292
rect 400824 19252 400830 19264
rect 401042 19252 401048 19264
rect 401100 19252 401106 19304
rect 140884 19224 140912 19252
rect 140958 19224 140964 19236
rect 140884 19196 140964 19224
rect 140958 19184 140964 19196
rect 141016 19184 141022 19236
rect 163038 17960 163044 18012
rect 163096 18000 163102 18012
rect 163130 18000 163136 18012
rect 163096 17972 163136 18000
rect 163096 17960 163102 17972
rect 163130 17960 163136 17972
rect 163188 17960 163194 18012
rect 180702 17960 180708 18012
rect 180760 18000 180766 18012
rect 181070 18000 181076 18012
rect 180760 17972 181076 18000
rect 180760 17960 180766 17972
rect 181070 17960 181076 17972
rect 181128 17960 181134 18012
rect 219710 17960 219716 18012
rect 219768 18000 219774 18012
rect 219802 18000 219808 18012
rect 219768 17972 219808 18000
rect 219768 17960 219774 17972
rect 219802 17960 219808 17972
rect 219860 17960 219866 18012
rect 220998 17960 221004 18012
rect 221056 18000 221062 18012
rect 221090 18000 221096 18012
rect 221056 17972 221096 18000
rect 221056 17960 221062 17972
rect 221090 17960 221096 17972
rect 221148 17960 221154 18012
rect 247954 17960 247960 18012
rect 248012 18000 248018 18012
rect 248322 18000 248328 18012
rect 248012 17972 248328 18000
rect 248012 17960 248018 17972
rect 248322 17960 248328 17972
rect 248380 17960 248386 18012
rect 253474 17960 253480 18012
rect 253532 18000 253538 18012
rect 253566 18000 253572 18012
rect 253532 17972 253572 18000
rect 253532 17960 253538 17972
rect 253566 17960 253572 17972
rect 253624 17960 253630 18012
rect 275922 17960 275928 18012
rect 275980 18000 275986 18012
rect 276106 18000 276112 18012
rect 275980 17972 276112 18000
rect 275980 17960 275986 17972
rect 276106 17960 276112 17972
rect 276164 17960 276170 18012
rect 339310 17960 339316 18012
rect 339368 18000 339374 18012
rect 339402 18000 339408 18012
rect 339368 17972 339408 18000
rect 339368 17960 339374 17972
rect 339402 17960 339408 17972
rect 339460 17960 339466 18012
rect 154850 17892 154856 17944
rect 154908 17932 154914 17944
rect 161658 17932 161664 17944
rect 154908 17904 161664 17932
rect 154908 17892 154914 17904
rect 161658 17892 161664 17904
rect 161716 17892 161722 17944
rect 436738 17892 436744 17944
rect 436796 17932 436802 17944
rect 579798 17932 579804 17944
rect 436796 17904 579804 17932
rect 436796 17892 436802 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 158714 17824 158720 17876
rect 158772 17864 158778 17876
rect 158990 17864 158996 17876
rect 158772 17836 158996 17864
rect 158772 17824 158778 17836
rect 158990 17824 158996 17836
rect 159048 17824 159054 17876
rect 420454 14492 420460 14544
rect 420512 14532 420518 14544
rect 420638 14532 420644 14544
rect 420512 14504 420644 14532
rect 420512 14492 420518 14504
rect 420638 14492 420644 14504
rect 420696 14492 420702 14544
rect 204438 12492 204444 12504
rect 204364 12464 204444 12492
rect 204364 12436 204392 12464
rect 204438 12452 204444 12464
rect 204496 12452 204502 12504
rect 276106 12452 276112 12504
rect 276164 12452 276170 12504
rect 204346 12384 204352 12436
rect 204404 12384 204410 12436
rect 276124 12356 276152 12452
rect 314654 12384 314660 12436
rect 314712 12424 314718 12436
rect 315758 12424 315764 12436
rect 314712 12396 315764 12424
rect 314712 12384 314718 12396
rect 315758 12384 315764 12396
rect 315816 12384 315822 12436
rect 276474 12356 276480 12368
rect 276124 12328 276480 12356
rect 276474 12316 276480 12328
rect 276532 12316 276538 12368
rect 386230 12180 386236 12232
rect 386288 12220 386294 12232
rect 488534 12220 488540 12232
rect 386288 12192 488540 12220
rect 386288 12180 386294 12192
rect 488534 12180 488540 12192
rect 488592 12180 488598 12232
rect 388898 12112 388904 12164
rect 388956 12152 388962 12164
rect 492674 12152 492680 12164
rect 388956 12124 492680 12152
rect 388956 12112 388962 12124
rect 492674 12112 492680 12124
rect 492732 12112 492738 12164
rect 390370 12044 390376 12096
rect 390428 12084 390434 12096
rect 495434 12084 495440 12096
rect 390428 12056 495440 12084
rect 390428 12044 390434 12056
rect 495434 12044 495440 12056
rect 495492 12044 495498 12096
rect 391750 11976 391756 12028
rect 391808 12016 391814 12028
rect 499574 12016 499580 12028
rect 391808 11988 499580 12016
rect 391808 11976 391814 11988
rect 499574 11976 499580 11988
rect 499632 11976 499638 12028
rect 394418 11908 394424 11960
rect 394476 11948 394482 11960
rect 502334 11948 502340 11960
rect 394476 11920 502340 11948
rect 394476 11908 394482 11920
rect 502334 11908 502340 11920
rect 502392 11908 502398 11960
rect 395890 11840 395896 11892
rect 395948 11880 395954 11892
rect 506474 11880 506480 11892
rect 395948 11852 506480 11880
rect 395948 11840 395954 11852
rect 506474 11840 506480 11852
rect 506532 11840 506538 11892
rect 397270 11772 397276 11824
rect 397328 11812 397334 11824
rect 510614 11812 510620 11824
rect 397328 11784 510620 11812
rect 397328 11772 397334 11784
rect 510614 11772 510620 11784
rect 510672 11772 510678 11824
rect 399938 11704 399944 11756
rect 399996 11744 400002 11756
rect 513374 11744 513380 11756
rect 399996 11716 513380 11744
rect 399996 11704 400002 11716
rect 513374 11704 513380 11716
rect 513432 11704 513438 11756
rect 366910 10956 366916 11008
rect 366968 10996 366974 11008
rect 451274 10996 451280 11008
rect 366968 10968 451280 10996
rect 366968 10956 366974 10968
rect 451274 10956 451280 10968
rect 451332 10956 451338 11008
rect 369762 10888 369768 10940
rect 369820 10928 369826 10940
rect 455414 10928 455420 10940
rect 369820 10900 455420 10928
rect 369820 10888 369826 10900
rect 455414 10888 455420 10900
rect 455472 10888 455478 10940
rect 371050 10820 371056 10872
rect 371108 10860 371114 10872
rect 459646 10860 459652 10872
rect 371108 10832 459652 10860
rect 371108 10820 371114 10832
rect 459646 10820 459652 10832
rect 459704 10820 459710 10872
rect 372430 10752 372436 10804
rect 372488 10792 372494 10804
rect 462314 10792 462320 10804
rect 372488 10764 462320 10792
rect 372488 10752 372494 10764
rect 462314 10752 462320 10764
rect 462372 10752 462378 10804
rect 114462 10684 114468 10736
rect 114520 10724 114526 10736
rect 190546 10724 190552 10736
rect 114520 10696 190552 10724
rect 114520 10684 114526 10696
rect 190546 10684 190552 10696
rect 190604 10684 190610 10736
rect 375190 10684 375196 10736
rect 375248 10724 375254 10736
rect 466454 10724 466460 10736
rect 375248 10696 466460 10724
rect 375248 10684 375254 10696
rect 466454 10684 466460 10696
rect 466512 10684 466518 10736
rect 86862 10616 86868 10668
rect 86920 10656 86926 10668
rect 178126 10656 178132 10668
rect 86920 10628 178132 10656
rect 86920 10616 86926 10628
rect 178126 10616 178132 10628
rect 178184 10616 178190 10668
rect 376570 10616 376576 10668
rect 376628 10656 376634 10668
rect 469214 10656 469220 10668
rect 376628 10628 469220 10656
rect 376628 10616 376634 10628
rect 469214 10616 469220 10628
rect 469272 10616 469278 10668
rect 79962 10548 79968 10600
rect 80020 10588 80026 10600
rect 174170 10588 174176 10600
rect 80020 10560 174176 10588
rect 80020 10548 80026 10560
rect 174170 10548 174176 10560
rect 174228 10548 174234 10600
rect 377950 10548 377956 10600
rect 378008 10588 378014 10600
rect 473354 10588 473360 10600
rect 378008 10560 473360 10588
rect 378008 10548 378014 10560
rect 473354 10548 473360 10560
rect 473412 10548 473418 10600
rect 72970 10480 72976 10532
rect 73028 10520 73034 10532
rect 169846 10520 169852 10532
rect 73028 10492 169852 10520
rect 73028 10480 73034 10492
rect 169846 10480 169852 10492
rect 169904 10480 169910 10532
rect 380802 10480 380808 10532
rect 380860 10520 380866 10532
rect 477586 10520 477592 10532
rect 380860 10492 477592 10520
rect 380860 10480 380866 10492
rect 477586 10480 477592 10492
rect 477644 10480 477650 10532
rect 64782 10412 64788 10464
rect 64840 10452 64846 10464
rect 167086 10452 167092 10464
rect 64840 10424 167092 10452
rect 64840 10412 64846 10424
rect 167086 10412 167092 10424
rect 167144 10412 167150 10464
rect 382090 10412 382096 10464
rect 382148 10452 382154 10464
rect 480254 10452 480260 10464
rect 382148 10424 480260 10452
rect 382148 10412 382154 10424
rect 480254 10412 480260 10424
rect 480312 10412 480318 10464
rect 38562 10344 38568 10396
rect 38620 10384 38626 10396
rect 146478 10384 146484 10396
rect 38620 10356 146484 10384
rect 38620 10344 38626 10356
rect 146478 10344 146484 10356
rect 146536 10344 146542 10396
rect 384850 10344 384856 10396
rect 384908 10384 384914 10396
rect 485774 10384 485780 10396
rect 384908 10356 485780 10384
rect 384908 10344 384914 10356
rect 485774 10344 485780 10356
rect 485832 10344 485838 10396
rect 42702 10276 42708 10328
rect 42760 10316 42766 10328
rect 154666 10316 154672 10328
rect 42760 10288 154672 10316
rect 42760 10276 42766 10288
rect 154666 10276 154672 10288
rect 154724 10276 154730 10328
rect 433150 10276 433156 10328
rect 433208 10316 433214 10328
rect 581086 10316 581092 10328
rect 433208 10288 581092 10316
rect 433208 10276 433214 10288
rect 581086 10276 581092 10288
rect 581144 10276 581150 10328
rect 365530 10208 365536 10260
rect 365588 10248 365594 10260
rect 448514 10248 448520 10260
rect 365588 10220 448520 10248
rect 365588 10208 365594 10220
rect 448514 10208 448520 10220
rect 448572 10208 448578 10260
rect 361390 10140 361396 10192
rect 361448 10180 361454 10192
rect 441614 10180 441620 10192
rect 361448 10152 441620 10180
rect 361448 10140 361454 10152
rect 441614 10140 441620 10152
rect 441672 10140 441678 10192
rect 364242 10072 364248 10124
rect 364300 10112 364306 10124
rect 444374 10112 444380 10124
rect 364300 10084 444380 10112
rect 364300 10072 364306 10084
rect 444374 10072 444380 10084
rect 444432 10072 444438 10124
rect 360010 10004 360016 10056
rect 360068 10044 360074 10056
rect 437474 10044 437480 10056
rect 360068 10016 437480 10044
rect 360068 10004 360074 10016
rect 437474 10004 437480 10016
rect 437532 10004 437538 10056
rect 358630 9936 358636 9988
rect 358688 9976 358694 9988
rect 434622 9976 434628 9988
rect 358688 9948 434628 9976
rect 358688 9936 358694 9948
rect 434622 9936 434628 9948
rect 434680 9936 434686 9988
rect 128722 9664 128728 9716
rect 128780 9704 128786 9716
rect 128906 9704 128912 9716
rect 128780 9676 128912 9704
rect 128780 9664 128786 9676
rect 128906 9664 128912 9676
rect 128964 9664 128970 9716
rect 162854 9664 162860 9716
rect 162912 9704 162918 9716
rect 163130 9704 163136 9716
rect 162912 9676 163136 9704
rect 162912 9664 162918 9676
rect 163130 9664 163136 9676
rect 163188 9664 163194 9716
rect 168190 9664 168196 9716
rect 168248 9704 168254 9716
rect 168466 9704 168472 9716
rect 168248 9676 168472 9704
rect 168248 9664 168254 9676
rect 168466 9664 168472 9676
rect 168524 9664 168530 9716
rect 185854 9664 185860 9716
rect 185912 9704 185918 9716
rect 186038 9704 186044 9716
rect 185912 9676 186044 9704
rect 185912 9664 185918 9676
rect 186038 9664 186044 9676
rect 186096 9664 186102 9716
rect 253474 9664 253480 9716
rect 253532 9704 253538 9716
rect 253658 9704 253664 9716
rect 253532 9676 253664 9704
rect 253532 9664 253538 9676
rect 253658 9664 253664 9676
rect 253716 9664 253722 9716
rect 275002 9664 275008 9716
rect 275060 9704 275066 9716
rect 275278 9704 275284 9716
rect 275060 9676 275284 9704
rect 275060 9664 275066 9676
rect 275278 9664 275284 9676
rect 275336 9664 275342 9716
rect 339126 9664 339132 9716
rect 339184 9704 339190 9716
rect 339402 9704 339408 9716
rect 339184 9676 339408 9704
rect 339184 9664 339190 9676
rect 339402 9664 339408 9676
rect 339460 9664 339466 9716
rect 400766 9664 400772 9716
rect 400824 9704 400830 9716
rect 400950 9704 400956 9716
rect 400824 9676 400956 9704
rect 400824 9664 400830 9676
rect 400950 9664 400956 9676
rect 401008 9664 401014 9716
rect 420454 9664 420460 9716
rect 420512 9704 420518 9716
rect 420638 9704 420644 9716
rect 420512 9676 420644 9704
rect 420512 9664 420518 9676
rect 420638 9664 420644 9676
rect 420696 9664 420702 9716
rect 94498 9596 94504 9648
rect 94556 9636 94562 9648
rect 182266 9636 182272 9648
rect 94556 9608 182272 9636
rect 94556 9596 94562 9608
rect 182266 9596 182272 9608
rect 182324 9596 182330 9648
rect 183646 9596 183652 9648
rect 183704 9636 183710 9648
rect 183830 9636 183836 9648
rect 183704 9608 183836 9636
rect 183704 9596 183710 9608
rect 183830 9596 183836 9608
rect 183888 9596 183894 9648
rect 184290 9596 184296 9648
rect 184348 9636 184354 9648
rect 185026 9636 185032 9648
rect 184348 9608 185032 9636
rect 184348 9596 184354 9608
rect 185026 9596 185032 9608
rect 185084 9596 185090 9648
rect 232866 9596 232872 9648
rect 232924 9636 232930 9648
rect 238938 9636 238944 9648
rect 232924 9608 238944 9636
rect 232924 9596 232930 9608
rect 238938 9596 238944 9608
rect 238996 9596 239002 9648
rect 245378 9596 245384 9648
rect 245436 9596 245442 9648
rect 246758 9596 246764 9648
rect 246816 9596 246822 9648
rect 247954 9596 247960 9648
rect 248012 9596 248018 9648
rect 368382 9596 368388 9648
rect 368440 9636 368446 9648
rect 454862 9636 454868 9648
rect 368440 9608 454868 9636
rect 368440 9596 368446 9608
rect 454862 9596 454868 9608
rect 454920 9596 454926 9648
rect 45738 9528 45744 9580
rect 45796 9568 45802 9580
rect 138658 9568 138664 9580
rect 45796 9540 138664 9568
rect 45796 9528 45802 9540
rect 138658 9528 138664 9540
rect 138716 9528 138722 9580
rect 143258 9528 143264 9580
rect 143316 9568 143322 9580
rect 207106 9568 207112 9580
rect 143316 9540 207112 9568
rect 143316 9528 143322 9540
rect 207106 9528 207112 9540
rect 207164 9528 207170 9580
rect 245396 9568 245424 9596
rect 245470 9568 245476 9580
rect 245396 9540 245476 9568
rect 245470 9528 245476 9540
rect 245528 9528 245534 9580
rect 246776 9512 246804 9596
rect 247972 9512 248000 9596
rect 339126 9528 339132 9580
rect 339184 9568 339190 9580
rect 343082 9568 343088 9580
rect 339184 9540 343088 9568
rect 339184 9528 339190 9540
rect 343082 9528 343088 9540
rect 343140 9528 343146 9580
rect 371142 9528 371148 9580
rect 371200 9568 371206 9580
rect 458450 9568 458456 9580
rect 371200 9540 458456 9568
rect 371200 9528 371206 9540
rect 458450 9528 458456 9540
rect 458508 9528 458514 9580
rect 62390 9460 62396 9512
rect 62448 9500 62454 9512
rect 165706 9500 165712 9512
rect 62448 9472 165712 9500
rect 62448 9460 62454 9472
rect 165706 9460 165712 9472
rect 165764 9460 165770 9512
rect 246758 9460 246764 9512
rect 246816 9460 246822 9512
rect 247954 9460 247960 9512
rect 248012 9460 248018 9512
rect 372522 9460 372528 9512
rect 372580 9500 372586 9512
rect 462038 9500 462044 9512
rect 372580 9472 462044 9500
rect 372580 9460 372586 9472
rect 462038 9460 462044 9472
rect 462096 9460 462102 9512
rect 58802 9392 58808 9444
rect 58860 9432 58866 9444
rect 164326 9432 164332 9444
rect 58860 9404 164332 9432
rect 58860 9392 58866 9404
rect 164326 9392 164332 9404
rect 164384 9392 164390 9444
rect 393130 9392 393136 9444
rect 393188 9432 393194 9444
rect 501230 9432 501236 9444
rect 393188 9404 501236 9432
rect 393188 9392 393194 9404
rect 501230 9392 501236 9404
rect 501288 9392 501294 9444
rect 55214 9324 55220 9376
rect 55272 9364 55278 9376
rect 154850 9364 154856 9376
rect 55272 9336 154856 9364
rect 55272 9324 55278 9336
rect 154850 9324 154856 9336
rect 154908 9324 154914 9376
rect 394510 9324 394516 9376
rect 394568 9364 394574 9376
rect 504818 9364 504824 9376
rect 394568 9336 504824 9364
rect 394568 9324 394574 9336
rect 504818 9324 504824 9336
rect 504876 9324 504882 9376
rect 51626 9256 51632 9308
rect 51684 9296 51690 9308
rect 160186 9296 160192 9308
rect 51684 9268 160192 9296
rect 51684 9256 51690 9268
rect 160186 9256 160192 9268
rect 160244 9256 160250 9308
rect 395982 9256 395988 9308
rect 396040 9296 396046 9308
rect 508406 9296 508412 9308
rect 396040 9268 508412 9296
rect 396040 9256 396046 9268
rect 508406 9256 508412 9268
rect 508464 9256 508470 9308
rect 40954 9188 40960 9240
rect 41012 9228 41018 9240
rect 154574 9228 154580 9240
rect 41012 9200 154580 9228
rect 41012 9188 41018 9200
rect 154574 9188 154580 9200
rect 154632 9188 154638 9240
rect 398650 9188 398656 9240
rect 398708 9228 398714 9240
rect 511994 9228 512000 9240
rect 398708 9200 512000 9228
rect 398708 9188 398714 9200
rect 511994 9188 512000 9200
rect 512052 9188 512058 9240
rect 33870 9120 33876 9172
rect 33928 9160 33934 9172
rect 150618 9160 150624 9172
rect 33928 9132 150624 9160
rect 33928 9120 33934 9132
rect 150618 9120 150624 9132
rect 150676 9120 150682 9172
rect 426158 9120 426164 9172
rect 426216 9160 426222 9172
rect 566734 9160 566740 9172
rect 426216 9132 566740 9160
rect 426216 9120 426222 9132
rect 566734 9120 566740 9132
rect 566792 9120 566798 9172
rect 13630 9052 13636 9104
rect 13688 9092 13694 9104
rect 133046 9092 133052 9104
rect 13688 9064 133052 9092
rect 13688 9052 13694 9064
rect 133046 9052 133052 9064
rect 133104 9052 133110 9104
rect 134886 9052 134892 9104
rect 134944 9092 134950 9104
rect 202966 9092 202972 9104
rect 134944 9064 202972 9092
rect 134944 9052 134950 9064
rect 202966 9052 202972 9064
rect 203024 9052 203030 9104
rect 409506 9052 409512 9104
rect 409564 9092 409570 9104
rect 409782 9092 409788 9104
rect 409564 9064 409788 9092
rect 409564 9052 409570 9064
rect 409782 9052 409788 9064
rect 409840 9052 409846 9104
rect 430482 9052 430488 9104
rect 430540 9092 430546 9104
rect 573818 9092 573824 9104
rect 430540 9064 573824 9092
rect 430540 9052 430546 9064
rect 573818 9052 573824 9064
rect 573876 9052 573882 9104
rect 6454 8984 6460 9036
rect 6512 9024 6518 9036
rect 136726 9024 136732 9036
rect 6512 8996 136732 9024
rect 6512 8984 6518 8996
rect 136726 8984 136732 8996
rect 136784 8984 136790 9036
rect 139670 8984 139676 9036
rect 139728 9024 139734 9036
rect 205726 9024 205732 9036
rect 139728 8996 205732 9024
rect 139728 8984 139734 8996
rect 205726 8984 205732 8996
rect 205784 8984 205790 9036
rect 354490 8984 354496 9036
rect 354548 9024 354554 9036
rect 427538 9024 427544 9036
rect 354548 8996 427544 9024
rect 354548 8984 354554 8996
rect 427538 8984 427544 8996
rect 427596 8984 427602 9036
rect 427630 8984 427636 9036
rect 427688 9024 427694 9036
rect 570230 9024 570236 9036
rect 427688 8996 570236 9024
rect 427688 8984 427694 8996
rect 570230 8984 570236 8996
rect 570288 8984 570294 9036
rect 5258 8916 5264 8968
rect 5316 8956 5322 8968
rect 136818 8956 136824 8968
rect 5316 8928 136824 8956
rect 5316 8916 5322 8928
rect 136818 8916 136824 8928
rect 136876 8916 136882 8968
rect 138474 8916 138480 8968
rect 138532 8956 138538 8968
rect 204346 8956 204352 8968
rect 138532 8928 204352 8956
rect 138532 8916 138538 8928
rect 204346 8916 204352 8928
rect 204404 8916 204410 8968
rect 355870 8916 355876 8968
rect 355928 8956 355934 8968
rect 431126 8956 431132 8968
rect 355928 8928 431132 8956
rect 355928 8916 355934 8928
rect 431126 8916 431132 8928
rect 431184 8916 431190 8968
rect 431678 8916 431684 8968
rect 431736 8956 431742 8968
rect 577406 8956 577412 8968
rect 431736 8928 577412 8956
rect 431736 8916 431742 8928
rect 577406 8916 577412 8928
rect 577464 8916 577470 8968
rect 98086 8848 98092 8900
rect 98144 8888 98150 8900
rect 183830 8888 183836 8900
rect 98144 8860 183836 8888
rect 98144 8848 98150 8860
rect 183830 8848 183836 8860
rect 183888 8848 183894 8900
rect 367002 8848 367008 8900
rect 367060 8888 367066 8900
rect 451366 8888 451372 8900
rect 367060 8860 451372 8888
rect 367060 8848 367066 8860
rect 451366 8848 451372 8860
rect 451424 8848 451430 8900
rect 77846 8780 77852 8832
rect 77904 8820 77910 8832
rect 77904 8792 126008 8820
rect 77904 8780 77910 8792
rect 84930 8712 84936 8764
rect 84988 8752 84994 8764
rect 125980 8752 126008 8792
rect 128998 8780 129004 8832
rect 129056 8820 129062 8832
rect 200206 8820 200212 8832
rect 129056 8792 200212 8820
rect 129056 8780 129062 8792
rect 200206 8780 200212 8792
rect 200264 8780 200270 8832
rect 365622 8780 365628 8832
rect 365680 8820 365686 8832
rect 447778 8820 447784 8832
rect 365680 8792 447784 8820
rect 365680 8780 365686 8792
rect 447778 8780 447784 8792
rect 447836 8780 447842 8832
rect 129182 8752 129188 8764
rect 84988 8724 125916 8752
rect 125980 8724 129188 8752
rect 84988 8712 84994 8724
rect 95694 8644 95700 8696
rect 95752 8684 95758 8696
rect 125888 8684 125916 8724
rect 129182 8712 129188 8724
rect 129240 8712 129246 8764
rect 131390 8712 131396 8764
rect 131448 8752 131454 8764
rect 201586 8752 201592 8764
rect 131448 8724 201592 8752
rect 131448 8712 131454 8724
rect 201586 8712 201592 8724
rect 201644 8712 201650 8764
rect 362862 8712 362868 8764
rect 362920 8752 362926 8764
rect 444190 8752 444196 8764
rect 362920 8724 444196 8752
rect 362920 8712 362926 8724
rect 444190 8712 444196 8724
rect 444248 8712 444254 8764
rect 129274 8684 129280 8696
rect 95752 8656 125732 8684
rect 125888 8656 129280 8684
rect 95752 8644 95758 8656
rect 120626 8576 120632 8628
rect 120684 8616 120690 8628
rect 120684 8588 122880 8616
rect 120684 8576 120690 8588
rect 122852 8480 122880 8588
rect 125704 8548 125732 8656
rect 129274 8644 129280 8656
rect 129332 8644 129338 8696
rect 132586 8644 132592 8696
rect 132644 8684 132650 8696
rect 201494 8684 201500 8696
rect 132644 8656 201500 8684
rect 132644 8644 132650 8656
rect 201494 8644 201500 8656
rect 201552 8644 201558 8696
rect 361482 8644 361488 8696
rect 361540 8684 361546 8696
rect 440602 8684 440608 8696
rect 361540 8656 440608 8684
rect 361540 8644 361546 8656
rect 440602 8644 440608 8656
rect 440660 8644 440666 8696
rect 136082 8576 136088 8628
rect 136140 8616 136146 8628
rect 203150 8616 203156 8628
rect 136140 8588 203156 8616
rect 136140 8576 136146 8588
rect 203150 8576 203156 8588
rect 203208 8576 203214 8628
rect 360102 8576 360108 8628
rect 360160 8616 360166 8628
rect 437014 8616 437020 8628
rect 360160 8588 437020 8616
rect 360160 8576 360166 8588
rect 437014 8576 437020 8588
rect 437072 8576 437078 8628
rect 129366 8548 129372 8560
rect 125704 8520 129372 8548
rect 129366 8508 129372 8520
rect 129424 8508 129430 8560
rect 126238 8480 126244 8492
rect 122852 8452 126244 8480
rect 126238 8440 126244 8452
rect 126296 8440 126302 8492
rect 34974 8236 34980 8288
rect 35032 8276 35038 8288
rect 115198 8276 115204 8288
rect 35032 8248 115204 8276
rect 35032 8236 35038 8248
rect 115198 8236 115204 8248
rect 115256 8236 115262 8288
rect 118234 8236 118240 8288
rect 118292 8276 118298 8288
rect 194686 8276 194692 8288
rect 118292 8248 194692 8276
rect 118292 8236 118298 8248
rect 194686 8236 194692 8248
rect 194744 8236 194750 8288
rect 388990 8236 388996 8288
rect 389048 8276 389054 8288
rect 494146 8276 494152 8288
rect 389048 8248 494152 8276
rect 389048 8236 389054 8248
rect 494146 8236 494152 8248
rect 494204 8236 494210 8288
rect 96890 8168 96896 8220
rect 96948 8208 96954 8220
rect 183554 8208 183560 8220
rect 96948 8180 183560 8208
rect 96948 8168 96954 8180
rect 183554 8168 183560 8180
rect 183612 8168 183618 8220
rect 390462 8168 390468 8220
rect 390520 8208 390526 8220
rect 497734 8208 497740 8220
rect 390520 8180 497740 8208
rect 390520 8168 390526 8180
rect 497734 8168 497740 8180
rect 497792 8168 497798 8220
rect 89714 8100 89720 8152
rect 89772 8140 89778 8152
rect 179598 8140 179604 8152
rect 89772 8112 179604 8140
rect 89772 8100 89778 8112
rect 179598 8100 179604 8112
rect 179656 8100 179662 8152
rect 409598 8100 409604 8152
rect 409656 8140 409662 8152
rect 534534 8140 534540 8152
rect 409656 8112 534540 8140
rect 409656 8100 409662 8112
rect 534534 8100 534540 8112
rect 534592 8100 534598 8152
rect 82630 8032 82636 8084
rect 82688 8072 82694 8084
rect 175366 8072 175372 8084
rect 82688 8044 175372 8072
rect 82688 8032 82694 8044
rect 175366 8032 175372 8044
rect 175424 8032 175430 8084
rect 411070 8032 411076 8084
rect 411128 8072 411134 8084
rect 538122 8072 538128 8084
rect 411128 8044 538128 8072
rect 411128 8032 411134 8044
rect 538122 8032 538128 8044
rect 538180 8032 538186 8084
rect 75454 7964 75460 8016
rect 75512 8004 75518 8016
rect 172606 8004 172612 8016
rect 75512 7976 172612 8004
rect 75512 7964 75518 7976
rect 172606 7964 172612 7976
rect 172664 7964 172670 8016
rect 342162 7964 342168 8016
rect 342220 8004 342226 8016
rect 402514 8004 402520 8016
rect 342220 7976 402520 8004
rect 342220 7964 342226 7976
rect 402514 7964 402520 7976
rect 402572 7964 402578 8016
rect 413922 7964 413928 8016
rect 413980 8004 413986 8016
rect 541710 8004 541716 8016
rect 413980 7976 541716 8004
rect 413980 7964 413986 7976
rect 541710 7964 541716 7976
rect 541768 7964 541774 8016
rect 68278 7896 68284 7948
rect 68336 7936 68342 7948
rect 168466 7936 168472 7948
rect 68336 7908 168472 7936
rect 68336 7896 68342 7908
rect 168466 7896 168472 7908
rect 168524 7896 168530 7948
rect 343450 7896 343456 7948
rect 343508 7936 343514 7948
rect 406102 7936 406108 7948
rect 343508 7908 406108 7936
rect 343508 7896 343514 7908
rect 406102 7896 406108 7908
rect 406160 7896 406166 7948
rect 415118 7896 415124 7948
rect 415176 7936 415182 7948
rect 545298 7936 545304 7948
rect 415176 7908 545304 7936
rect 415176 7896 415182 7908
rect 545298 7896 545304 7908
rect 545356 7896 545362 7948
rect 48130 7828 48136 7880
rect 48188 7868 48194 7880
rect 158806 7868 158812 7880
rect 48188 7840 158812 7868
rect 48188 7828 48194 7840
rect 158806 7828 158812 7840
rect 158864 7828 158870 7880
rect 344830 7828 344836 7880
rect 344888 7868 344894 7880
rect 409690 7868 409696 7880
rect 344888 7840 409696 7868
rect 344888 7828 344894 7840
rect 409690 7828 409696 7840
rect 409748 7828 409754 7880
rect 416590 7828 416596 7880
rect 416648 7868 416654 7880
rect 548886 7868 548892 7880
rect 416648 7840 548892 7868
rect 416648 7828 416654 7840
rect 548886 7828 548892 7840
rect 548944 7828 548950 7880
rect 7650 7760 7656 7812
rect 7708 7800 7714 7812
rect 136634 7800 136640 7812
rect 7708 7772 136640 7800
rect 7708 7760 7714 7772
rect 136634 7760 136640 7772
rect 136692 7760 136698 7812
rect 171778 7760 171784 7812
rect 171836 7800 171842 7812
rect 222286 7800 222292 7812
rect 171836 7772 222292 7800
rect 171836 7760 171842 7772
rect 222286 7760 222292 7772
rect 222344 7760 222350 7812
rect 347682 7760 347688 7812
rect 347740 7800 347746 7812
rect 413278 7800 413284 7812
rect 347740 7772 413284 7800
rect 347740 7760 347746 7772
rect 413278 7760 413284 7772
rect 413336 7760 413342 7812
rect 419442 7760 419448 7812
rect 419500 7800 419506 7812
rect 552382 7800 552388 7812
rect 419500 7772 552388 7800
rect 419500 7760 419506 7772
rect 552382 7760 552388 7772
rect 552440 7760 552446 7812
rect 1670 7692 1676 7744
rect 1728 7732 1734 7744
rect 133874 7732 133880 7744
rect 1728 7704 133880 7732
rect 1728 7692 1734 7704
rect 133874 7692 133880 7704
rect 133932 7692 133938 7744
rect 140866 7692 140872 7744
rect 140924 7732 140930 7744
rect 205634 7732 205640 7744
rect 140924 7704 205640 7732
rect 140924 7692 140930 7704
rect 205634 7692 205640 7704
rect 205692 7692 205698 7744
rect 348970 7692 348976 7744
rect 349028 7732 349034 7744
rect 416866 7732 416872 7744
rect 349028 7704 416872 7732
rect 349028 7692 349034 7704
rect 416866 7692 416872 7704
rect 416924 7692 416930 7744
rect 420638 7692 420644 7744
rect 420696 7732 420702 7744
rect 555970 7732 555976 7744
rect 420696 7704 555976 7732
rect 420696 7692 420702 7704
rect 555970 7692 555976 7704
rect 556028 7692 556034 7744
rect 2866 7624 2872 7676
rect 2924 7664 2930 7676
rect 135346 7664 135352 7676
rect 2924 7636 135352 7664
rect 2924 7624 2930 7636
rect 135346 7624 135352 7636
rect 135404 7624 135410 7676
rect 144454 7624 144460 7676
rect 144512 7664 144518 7676
rect 208578 7664 208584 7676
rect 144512 7636 208584 7664
rect 144512 7624 144518 7636
rect 208578 7624 208584 7636
rect 208636 7624 208642 7676
rect 350350 7624 350356 7676
rect 350408 7664 350414 7676
rect 420362 7664 420368 7676
rect 350408 7636 420368 7664
rect 350408 7624 350414 7636
rect 420362 7624 420368 7636
rect 420420 7624 420426 7676
rect 422110 7624 422116 7676
rect 422168 7664 422174 7676
rect 559558 7664 559564 7676
rect 422168 7636 559564 7664
rect 422168 7624 422174 7636
rect 559558 7624 559564 7636
rect 559616 7624 559622 7676
rect 566 7556 572 7608
rect 624 7596 630 7608
rect 133966 7596 133972 7608
rect 624 7568 133972 7596
rect 624 7556 630 7568
rect 133966 7556 133972 7568
rect 134024 7556 134030 7608
rect 137278 7556 137284 7608
rect 137336 7596 137342 7608
rect 204254 7596 204260 7608
rect 137336 7568 204260 7596
rect 137336 7556 137342 7568
rect 204254 7556 204260 7568
rect 204312 7556 204318 7608
rect 353202 7556 353208 7608
rect 353260 7596 353266 7608
rect 423950 7596 423956 7608
rect 353260 7568 423956 7596
rect 353260 7556 353266 7568
rect 423950 7556 423956 7568
rect 424008 7556 424014 7608
rect 424962 7556 424968 7608
rect 425020 7596 425026 7608
rect 563146 7596 563152 7608
rect 425020 7568 563152 7596
rect 425020 7556 425026 7568
rect 563146 7556 563152 7568
rect 563204 7556 563210 7608
rect 97994 7488 98000 7540
rect 98052 7528 98058 7540
rect 99282 7528 99288 7540
rect 98052 7500 99288 7528
rect 98052 7488 98058 7500
rect 99282 7488 99288 7500
rect 99340 7488 99346 7540
rect 111150 7488 111156 7540
rect 111208 7528 111214 7540
rect 190638 7528 190644 7540
rect 111208 7500 190644 7528
rect 111208 7488 111214 7500
rect 190638 7488 190644 7500
rect 190696 7488 190702 7540
rect 376386 7488 376392 7540
rect 376444 7528 376450 7540
rect 376662 7528 376668 7540
rect 376444 7500 376668 7528
rect 376444 7488 376450 7500
rect 376662 7488 376668 7500
rect 376720 7488 376726 7540
rect 387610 7488 387616 7540
rect 387668 7528 387674 7540
rect 490558 7528 490564 7540
rect 387668 7500 490564 7528
rect 387668 7488 387674 7500
rect 490558 7488 490564 7500
rect 490616 7488 490622 7540
rect 121822 7420 121828 7472
rect 121880 7460 121886 7472
rect 195974 7460 195980 7472
rect 121880 7432 195980 7460
rect 121880 7420 121886 7432
rect 195974 7420 195980 7432
rect 196032 7420 196038 7472
rect 384942 7420 384948 7472
rect 385000 7460 385006 7472
rect 486970 7460 486976 7472
rect 385000 7432 486976 7460
rect 385000 7420 385006 7432
rect 486970 7420 486976 7432
rect 487028 7420 487034 7472
rect 126606 7352 126612 7404
rect 126664 7392 126670 7404
rect 198826 7392 198832 7404
rect 126664 7364 198832 7392
rect 126664 7352 126670 7364
rect 198826 7352 198832 7364
rect 198884 7352 198890 7404
rect 383378 7352 383384 7404
rect 383436 7392 383442 7404
rect 483474 7392 483480 7404
rect 383436 7364 483480 7392
rect 383436 7352 383442 7364
rect 483474 7352 483480 7364
rect 483532 7352 483538 7404
rect 109954 7284 109960 7336
rect 110012 7324 110018 7336
rect 127618 7324 127624 7336
rect 110012 7296 127624 7324
rect 110012 7284 110018 7296
rect 127618 7284 127624 7296
rect 127676 7284 127682 7336
rect 127802 7284 127808 7336
rect 127860 7324 127866 7336
rect 198734 7324 198740 7336
rect 127860 7296 198740 7324
rect 127860 7284 127866 7296
rect 198734 7284 198740 7296
rect 198792 7284 198798 7336
rect 357342 7284 357348 7336
rect 357400 7324 357406 7336
rect 433518 7324 433524 7336
rect 357400 7296 433524 7324
rect 357400 7284 357406 7296
rect 433518 7284 433524 7296
rect 433576 7284 433582 7336
rect 63586 7216 63592 7268
rect 63644 7256 63650 7268
rect 128906 7256 128912 7268
rect 63644 7228 128912 7256
rect 63644 7216 63650 7228
rect 128906 7216 128912 7228
rect 128964 7216 128970 7268
rect 133782 7216 133788 7268
rect 133840 7256 133846 7268
rect 202874 7256 202880 7268
rect 133840 7228 202880 7256
rect 133840 7216 133846 7228
rect 202874 7216 202880 7228
rect 202932 7216 202938 7268
rect 358722 7216 358728 7268
rect 358780 7256 358786 7268
rect 435818 7256 435824 7268
rect 358780 7228 435824 7256
rect 358780 7216 358786 7228
rect 435818 7216 435824 7228
rect 435876 7216 435882 7268
rect 130194 7148 130200 7200
rect 130252 7188 130258 7200
rect 200114 7188 200120 7200
rect 130252 7160 200120 7188
rect 130252 7148 130258 7160
rect 200114 7148 200120 7160
rect 200172 7148 200178 7200
rect 138014 6876 138020 6928
rect 138072 6916 138078 6928
rect 138198 6916 138204 6928
rect 138072 6888 138204 6916
rect 138072 6876 138078 6888
rect 138198 6876 138204 6888
rect 138256 6876 138262 6928
rect 360194 6876 360200 6928
rect 360252 6916 360258 6928
rect 360252 6888 362264 6916
rect 360252 6876 360258 6888
rect 101582 6808 101588 6860
rect 101640 6848 101646 6860
rect 186406 6848 186412 6860
rect 101640 6820 186412 6848
rect 101640 6808 101646 6820
rect 186406 6808 186412 6820
rect 186464 6808 186470 6860
rect 321370 6808 321376 6860
rect 321428 6848 321434 6860
rect 362126 6848 362132 6860
rect 321428 6820 362132 6848
rect 321428 6808 321434 6820
rect 362126 6808 362132 6820
rect 362184 6808 362190 6860
rect 362236 6848 362264 6888
rect 371896 6888 376708 6916
rect 371896 6848 371924 6888
rect 362236 6820 371924 6848
rect 376680 6848 376708 6888
rect 376754 6876 376760 6928
rect 376812 6876 376818 6928
rect 376772 6848 376800 6876
rect 376680 6820 376800 6848
rect 389082 6808 389088 6860
rect 389140 6848 389146 6860
rect 495342 6848 495348 6860
rect 389140 6820 495348 6848
rect 389140 6808 389146 6820
rect 495342 6808 495348 6820
rect 495400 6808 495406 6860
rect 61194 6740 61200 6792
rect 61252 6780 61258 6792
rect 164510 6780 164516 6792
rect 61252 6752 164516 6780
rect 61252 6740 61258 6752
rect 164510 6740 164516 6752
rect 164568 6740 164574 6792
rect 321462 6740 321468 6792
rect 321520 6780 321526 6792
rect 363322 6780 363328 6792
rect 321520 6752 363328 6780
rect 321520 6740 321526 6752
rect 363322 6740 363328 6752
rect 363380 6740 363386 6792
rect 379606 6740 379612 6792
rect 379664 6780 379670 6792
rect 387242 6780 387248 6792
rect 379664 6752 387248 6780
rect 379664 6740 379670 6752
rect 387242 6740 387248 6752
rect 387300 6740 387306 6792
rect 498930 6780 498936 6792
rect 391952 6752 498936 6780
rect 57606 6672 57612 6724
rect 57664 6712 57670 6724
rect 162854 6712 162860 6724
rect 57664 6684 162860 6712
rect 57664 6672 57670 6684
rect 162854 6672 162860 6684
rect 162912 6672 162918 6724
rect 197170 6672 197176 6724
rect 197228 6712 197234 6724
rect 212626 6712 212632 6724
rect 197228 6684 212632 6712
rect 197228 6672 197234 6684
rect 212626 6672 212632 6684
rect 212684 6672 212690 6724
rect 354490 6672 354496 6724
rect 354548 6712 354554 6724
rect 360194 6712 360200 6724
rect 354548 6684 360200 6712
rect 354548 6672 354554 6684
rect 360194 6672 360200 6684
rect 360252 6672 360258 6724
rect 391750 6672 391756 6724
rect 391808 6712 391814 6724
rect 391952 6712 391980 6752
rect 498930 6740 498936 6752
rect 498988 6740 498994 6792
rect 391808 6684 391980 6712
rect 391808 6672 391814 6684
rect 393222 6672 393228 6724
rect 393280 6712 393286 6724
rect 502426 6712 502432 6724
rect 393280 6684 502432 6712
rect 393280 6672 393286 6684
rect 502426 6672 502432 6684
rect 502484 6672 502490 6724
rect 54018 6604 54024 6656
rect 54076 6644 54082 6656
rect 161474 6644 161480 6656
rect 54076 6616 161480 6644
rect 54076 6604 54082 6616
rect 161474 6604 161480 6616
rect 161532 6604 161538 6656
rect 194594 6604 194600 6656
rect 194652 6644 194658 6656
rect 214098 6644 214104 6656
rect 194652 6616 214104 6644
rect 194652 6604 194658 6616
rect 214098 6604 214104 6616
rect 214156 6604 214162 6656
rect 322750 6604 322756 6656
rect 322808 6644 322814 6656
rect 366910 6644 366916 6656
rect 322808 6616 366916 6644
rect 322808 6604 322814 6616
rect 366910 6604 366916 6616
rect 366968 6604 366974 6656
rect 394602 6604 394608 6656
rect 394660 6644 394666 6656
rect 506014 6644 506020 6656
rect 394660 6616 506020 6644
rect 394660 6604 394666 6616
rect 506014 6604 506020 6616
rect 506072 6604 506078 6656
rect 50522 6536 50528 6588
rect 50580 6576 50586 6588
rect 158714 6576 158720 6588
rect 50580 6548 158720 6576
rect 50580 6536 50586 6548
rect 158714 6536 158720 6548
rect 158772 6536 158778 6588
rect 193306 6536 193312 6588
rect 193364 6576 193370 6588
rect 215478 6576 215484 6588
rect 193364 6548 215484 6576
rect 193364 6536 193370 6548
rect 215478 6536 215484 6548
rect 215536 6536 215542 6588
rect 315942 6536 315948 6588
rect 316000 6576 316006 6588
rect 351086 6576 351092 6588
rect 316000 6548 351092 6576
rect 316000 6536 316006 6548
rect 351086 6536 351092 6548
rect 351144 6536 351150 6588
rect 351178 6536 351184 6588
rect 351236 6576 351242 6588
rect 395430 6576 395436 6588
rect 351236 6548 395436 6576
rect 351236 6536 351242 6548
rect 395430 6536 395436 6548
rect 395488 6536 395494 6588
rect 397362 6536 397368 6588
rect 397420 6576 397426 6588
rect 509602 6576 509608 6588
rect 397420 6548 509608 6576
rect 397420 6536 397426 6548
rect 509602 6536 509608 6548
rect 509660 6536 509666 6588
rect 46934 6468 46940 6520
rect 46992 6508 46998 6520
rect 157334 6508 157340 6520
rect 46992 6480 157340 6508
rect 46992 6468 46998 6480
rect 157334 6468 157340 6480
rect 157392 6468 157398 6520
rect 188614 6468 188620 6520
rect 188672 6508 188678 6520
rect 218238 6508 218244 6520
rect 188672 6480 218244 6508
rect 188672 6468 188678 6480
rect 218238 6468 218244 6480
rect 218296 6468 218302 6520
rect 325510 6468 325516 6520
rect 325568 6508 325574 6520
rect 370406 6508 370412 6520
rect 325568 6480 370412 6508
rect 325568 6468 325574 6480
rect 370406 6468 370412 6480
rect 370464 6468 370470 6520
rect 387242 6468 387248 6520
rect 387300 6508 387306 6520
rect 391842 6508 391848 6520
rect 387300 6480 391848 6508
rect 387300 6468 387306 6480
rect 391842 6468 391848 6480
rect 391900 6468 391906 6520
rect 398742 6468 398748 6520
rect 398800 6508 398806 6520
rect 513190 6508 513196 6520
rect 398800 6480 513196 6508
rect 398800 6468 398806 6480
rect 513190 6468 513196 6480
rect 513248 6468 513254 6520
rect 44542 6400 44548 6452
rect 44600 6440 44606 6452
rect 156138 6440 156144 6452
rect 44600 6412 156144 6440
rect 44600 6400 44606 6412
rect 156138 6400 156144 6412
rect 156196 6400 156202 6452
rect 188062 6400 188068 6452
rect 188120 6440 188126 6452
rect 219710 6440 219716 6452
rect 188120 6412 219716 6440
rect 188120 6400 188126 6412
rect 219710 6400 219716 6412
rect 219768 6400 219774 6452
rect 326890 6400 326896 6452
rect 326948 6440 326954 6452
rect 373994 6440 374000 6452
rect 326948 6412 374000 6440
rect 326948 6400 326954 6412
rect 373994 6400 374000 6412
rect 374052 6400 374058 6452
rect 400030 6400 400036 6452
rect 400088 6440 400094 6452
rect 516778 6440 516784 6452
rect 400088 6412 516784 6440
rect 400088 6400 400094 6412
rect 516778 6400 516784 6412
rect 516836 6400 516842 6452
rect 39758 6332 39764 6384
rect 39816 6372 39822 6384
rect 153286 6372 153292 6384
rect 39816 6344 153292 6372
rect 39816 6332 39822 6344
rect 153286 6332 153292 6344
rect 153344 6332 153350 6384
rect 157518 6332 157524 6384
rect 157576 6372 157582 6384
rect 214006 6372 214012 6384
rect 157576 6344 214012 6372
rect 157576 6332 157582 6344
rect 214006 6332 214012 6344
rect 214064 6332 214070 6384
rect 328270 6332 328276 6384
rect 328328 6372 328334 6384
rect 377582 6372 377588 6384
rect 328328 6344 377588 6372
rect 328328 6332 328334 6344
rect 377582 6332 377588 6344
rect 377640 6332 377646 6384
rect 402790 6332 402796 6384
rect 402848 6372 402854 6384
rect 520274 6372 520280 6384
rect 402848 6344 520280 6372
rect 402848 6332 402854 6344
rect 520274 6332 520280 6344
rect 520332 6332 520338 6384
rect 18322 6264 18328 6316
rect 18380 6304 18386 6316
rect 135438 6304 135444 6316
rect 18380 6276 135444 6304
rect 18380 6264 18386 6276
rect 135438 6264 135444 6276
rect 135496 6264 135502 6316
rect 161106 6264 161112 6316
rect 161164 6304 161170 6316
rect 216766 6304 216772 6316
rect 161164 6276 216772 6304
rect 161164 6264 161170 6276
rect 216766 6264 216772 6276
rect 216824 6264 216830 6316
rect 331122 6264 331128 6316
rect 331180 6304 331186 6316
rect 381170 6304 381176 6316
rect 331180 6276 381176 6304
rect 331180 6264 331186 6276
rect 381170 6264 381176 6276
rect 381228 6264 381234 6316
rect 404170 6264 404176 6316
rect 404228 6304 404234 6316
rect 523862 6304 523868 6316
rect 404228 6276 523868 6304
rect 404228 6264 404234 6276
rect 523862 6264 523868 6276
rect 523920 6264 523926 6316
rect 32674 6196 32680 6248
rect 32732 6236 32738 6248
rect 84194 6236 84200 6248
rect 32732 6208 84200 6236
rect 32732 6196 32738 6208
rect 84194 6196 84200 6208
rect 84252 6196 84258 6248
rect 103422 6196 103428 6248
rect 103480 6236 103486 6248
rect 113174 6236 113180 6248
rect 103480 6208 113180 6236
rect 103480 6196 103486 6208
rect 113174 6196 113180 6208
rect 113232 6196 113238 6248
rect 122742 6196 122748 6248
rect 122800 6236 122806 6248
rect 128354 6236 128360 6248
rect 122800 6208 128360 6236
rect 122800 6196 122806 6208
rect 128354 6196 128360 6208
rect 128412 6196 128418 6248
rect 153930 6196 153936 6248
rect 153988 6236 153994 6248
rect 212534 6236 212540 6248
rect 153988 6208 212540 6236
rect 153988 6196 153994 6208
rect 212534 6196 212540 6208
rect 212592 6196 212598 6248
rect 332410 6196 332416 6248
rect 332468 6236 332474 6248
rect 384666 6236 384672 6248
rect 332468 6208 384672 6236
rect 332468 6196 332474 6208
rect 384666 6196 384672 6208
rect 384724 6196 384730 6248
rect 408402 6196 408408 6248
rect 408460 6236 408466 6248
rect 531038 6236 531044 6248
rect 408460 6208 531044 6236
rect 408460 6196 408466 6208
rect 531038 6196 531044 6208
rect 531096 6196 531102 6248
rect 4062 6128 4068 6180
rect 4120 6168 4126 6180
rect 135254 6168 135260 6180
rect 4120 6140 135260 6168
rect 4120 6128 4126 6140
rect 135254 6128 135260 6140
rect 135312 6128 135318 6180
rect 135346 6128 135352 6180
rect 135404 6168 135410 6180
rect 150342 6168 150348 6180
rect 135404 6140 150348 6168
rect 135404 6128 135410 6140
rect 150342 6128 150348 6140
rect 150400 6128 150406 6180
rect 150434 6128 150440 6180
rect 150492 6168 150498 6180
rect 211246 6168 211252 6180
rect 150492 6140 211252 6168
rect 150492 6128 150498 6140
rect 211246 6128 211252 6140
rect 211304 6128 211310 6180
rect 333698 6128 333704 6180
rect 333756 6168 333762 6180
rect 388254 6168 388260 6180
rect 333756 6140 388260 6168
rect 333756 6128 333762 6140
rect 388254 6128 388260 6140
rect 388312 6128 388318 6180
rect 405550 6128 405556 6180
rect 405608 6168 405614 6180
rect 527450 6168 527456 6180
rect 405608 6140 527456 6168
rect 405608 6128 405614 6140
rect 527450 6128 527456 6140
rect 527508 6128 527514 6180
rect 102778 6060 102784 6112
rect 102836 6100 102842 6112
rect 186498 6100 186504 6112
rect 102836 6072 186504 6100
rect 102836 6060 102842 6072
rect 186498 6060 186504 6072
rect 186556 6060 186562 6112
rect 318610 6060 318616 6112
rect 318668 6100 318674 6112
rect 358538 6100 358544 6112
rect 318668 6072 358544 6100
rect 318668 6060 318674 6072
rect 358538 6060 358544 6072
rect 358596 6060 358602 6112
rect 387702 6060 387708 6112
rect 387760 6100 387766 6112
rect 491754 6100 491760 6112
rect 387760 6072 491760 6100
rect 387760 6060 387766 6072
rect 491754 6060 491760 6072
rect 491812 6060 491818 6112
rect 84194 5992 84200 6044
rect 84252 6032 84258 6044
rect 103422 6032 103428 6044
rect 84252 6004 103428 6032
rect 84252 5992 84258 6004
rect 103422 5992 103428 6004
rect 103480 5992 103486 6044
rect 105170 5992 105176 6044
rect 105228 6032 105234 6044
rect 187694 6032 187700 6044
rect 105228 6004 187700 6032
rect 105228 5992 105234 6004
rect 187694 5992 187700 6004
rect 187752 5992 187758 6044
rect 317322 5992 317328 6044
rect 317380 6032 317386 6044
rect 356146 6032 356152 6044
rect 317380 6004 356152 6032
rect 317380 5992 317386 6004
rect 356146 5992 356152 6004
rect 356204 5992 356210 6044
rect 383470 5992 383476 6044
rect 383528 6032 383534 6044
rect 484578 6032 484584 6044
rect 383528 6004 484584 6032
rect 383528 5992 383534 6004
rect 484578 5992 484584 6004
rect 484636 5992 484642 6044
rect 106366 5924 106372 5976
rect 106424 5964 106430 5976
rect 187786 5964 187792 5976
rect 106424 5936 187792 5964
rect 106424 5924 106430 5936
rect 187786 5924 187792 5936
rect 187844 5924 187850 5976
rect 320082 5924 320088 5976
rect 320140 5964 320146 5976
rect 359734 5964 359740 5976
rect 320140 5936 359740 5964
rect 320140 5924 320146 5936
rect 359734 5924 359740 5936
rect 359792 5924 359798 5976
rect 386322 5924 386328 5976
rect 386380 5964 386386 5976
rect 488166 5964 488172 5976
rect 386380 5936 488172 5964
rect 386380 5924 386386 5936
rect 488166 5924 488172 5936
rect 488224 5924 488230 5976
rect 108758 5856 108764 5908
rect 108816 5896 108822 5908
rect 189350 5896 189356 5908
rect 108816 5868 189356 5896
rect 108816 5856 108822 5868
rect 189350 5856 189356 5868
rect 189408 5856 189414 5908
rect 317046 5856 317052 5908
rect 317104 5896 317110 5908
rect 354950 5896 354956 5908
rect 317104 5868 354956 5896
rect 317104 5856 317110 5868
rect 354950 5856 354956 5868
rect 355008 5856 355014 5908
rect 379330 5856 379336 5908
rect 379388 5896 379394 5908
rect 476298 5896 476304 5908
rect 379388 5868 476304 5896
rect 379388 5856 379394 5868
rect 476298 5856 476304 5868
rect 476356 5856 476362 5908
rect 81434 5788 81440 5840
rect 81492 5828 81498 5840
rect 109678 5828 109684 5840
rect 81492 5800 109684 5828
rect 81492 5788 81498 5800
rect 109678 5788 109684 5800
rect 109736 5788 109742 5840
rect 112346 5788 112352 5840
rect 112404 5828 112410 5840
rect 191926 5828 191932 5840
rect 112404 5800 191932 5828
rect 112404 5788 112410 5800
rect 191926 5788 191932 5800
rect 191984 5788 191990 5840
rect 315850 5788 315856 5840
rect 315908 5828 315914 5840
rect 352558 5828 352564 5840
rect 315908 5800 352564 5828
rect 315908 5788 315914 5800
rect 352558 5788 352564 5800
rect 352616 5788 352622 5840
rect 382182 5788 382188 5840
rect 382240 5828 382246 5840
rect 479886 5828 479892 5840
rect 382240 5800 479892 5828
rect 382240 5788 382246 5800
rect 479886 5788 479892 5800
rect 479944 5788 479950 5840
rect 116026 5720 116032 5772
rect 116084 5760 116090 5772
rect 193214 5760 193220 5772
rect 116084 5732 193220 5760
rect 116084 5720 116090 5732
rect 193214 5720 193220 5732
rect 193272 5720 193278 5772
rect 348418 5720 348424 5772
rect 348476 5760 348482 5772
rect 354490 5760 354496 5772
rect 348476 5732 354496 5760
rect 348476 5720 348482 5732
rect 354490 5720 354496 5732
rect 354548 5720 354554 5772
rect 378042 5720 378048 5772
rect 378100 5760 378106 5772
rect 472710 5760 472716 5772
rect 378100 5732 472716 5760
rect 378100 5720 378106 5732
rect 472710 5720 472716 5732
rect 472768 5720 472774 5772
rect 119430 5652 119436 5704
rect 119488 5692 119494 5704
rect 194686 5692 194692 5704
rect 119488 5664 194692 5692
rect 119488 5652 119494 5664
rect 194686 5652 194692 5664
rect 194744 5652 194750 5704
rect 373902 5652 373908 5704
rect 373960 5692 373966 5704
rect 465626 5692 465632 5704
rect 373960 5664 465632 5692
rect 373960 5652 373966 5664
rect 465626 5652 465632 5664
rect 465684 5652 465690 5704
rect 113174 5584 113180 5636
rect 113232 5624 113238 5636
rect 122742 5624 122748 5636
rect 113232 5596 122748 5624
rect 113232 5584 113238 5596
rect 122742 5584 122748 5596
rect 122800 5584 122806 5636
rect 123018 5584 123024 5636
rect 123076 5624 123082 5636
rect 197538 5624 197544 5636
rect 123076 5596 197544 5624
rect 123076 5584 123082 5596
rect 197538 5584 197544 5596
rect 197596 5584 197602 5636
rect 376386 5584 376392 5636
rect 376444 5624 376450 5636
rect 469122 5624 469128 5636
rect 376444 5596 469128 5624
rect 376444 5584 376450 5596
rect 469122 5584 469128 5596
rect 469180 5584 469186 5636
rect 128354 5516 128360 5568
rect 128412 5556 128418 5568
rect 135346 5556 135352 5568
rect 128412 5528 135352 5556
rect 128412 5516 128418 5528
rect 135346 5516 135352 5528
rect 135404 5516 135410 5568
rect 353938 5516 353944 5568
rect 353996 5556 354002 5568
rect 399018 5556 399024 5568
rect 353996 5528 399024 5556
rect 353996 5516 354002 5528
rect 399018 5516 399024 5528
rect 399076 5516 399082 5568
rect 80238 5448 80244 5500
rect 80296 5488 80302 5500
rect 175458 5488 175464 5500
rect 80296 5460 175464 5488
rect 80296 5448 80302 5460
rect 175458 5448 175464 5460
rect 175516 5448 175522 5500
rect 209222 5448 209228 5500
rect 209280 5488 209286 5500
rect 232866 5488 232872 5500
rect 209280 5460 232872 5488
rect 209280 5448 209286 5460
rect 232866 5448 232872 5460
rect 232924 5448 232930 5500
rect 335262 5448 335268 5500
rect 335320 5488 335326 5500
rect 390646 5488 390652 5500
rect 335320 5460 390652 5488
rect 335320 5448 335326 5460
rect 390646 5448 390652 5460
rect 390704 5448 390710 5500
rect 415302 5448 415308 5500
rect 415360 5488 415366 5500
rect 544102 5488 544108 5500
rect 415360 5460 544108 5488
rect 415360 5448 415366 5460
rect 544102 5448 544108 5460
rect 544160 5448 544166 5500
rect 76650 5380 76656 5432
rect 76708 5420 76714 5432
rect 172514 5420 172520 5432
rect 76708 5392 172520 5420
rect 76708 5380 76714 5392
rect 172514 5380 172520 5392
rect 172572 5380 172578 5432
rect 208302 5380 208308 5432
rect 208360 5420 208366 5432
rect 237466 5420 237472 5432
rect 208360 5392 237472 5420
rect 208360 5380 208366 5392
rect 237466 5380 237472 5392
rect 237524 5380 237530 5432
rect 343082 5380 343088 5432
rect 343140 5420 343146 5432
rect 397822 5420 397828 5432
rect 343140 5392 397828 5420
rect 343140 5380 343146 5392
rect 397822 5380 397828 5392
rect 397880 5380 397886 5432
rect 416682 5380 416688 5432
rect 416740 5420 416746 5432
rect 547690 5420 547696 5432
rect 416740 5392 547696 5420
rect 416740 5380 416746 5392
rect 547690 5380 547696 5392
rect 547748 5380 547754 5432
rect 73062 5312 73068 5364
rect 73120 5352 73126 5364
rect 171226 5352 171232 5364
rect 73120 5324 171232 5352
rect 73120 5312 73126 5324
rect 171226 5312 171232 5324
rect 171284 5312 171290 5364
rect 173894 5312 173900 5364
rect 173952 5352 173958 5364
rect 213914 5352 213920 5364
rect 173952 5324 213920 5352
rect 173952 5312 173958 5324
rect 213914 5312 213920 5324
rect 213972 5312 213978 5364
rect 340782 5312 340788 5364
rect 340840 5352 340846 5364
rect 401318 5352 401324 5364
rect 340840 5324 401324 5352
rect 340840 5312 340846 5324
rect 401318 5312 401324 5324
rect 401376 5312 401382 5364
rect 418062 5312 418068 5364
rect 418120 5352 418126 5364
rect 551186 5352 551192 5364
rect 418120 5324 551192 5352
rect 418120 5312 418126 5324
rect 551186 5312 551192 5324
rect 551244 5312 551250 5364
rect 69474 5244 69480 5296
rect 69532 5284 69538 5296
rect 169938 5284 169944 5296
rect 69532 5256 169944 5284
rect 69532 5244 69538 5256
rect 169938 5244 169944 5256
rect 169996 5244 170002 5296
rect 174170 5244 174176 5296
rect 174228 5284 174234 5296
rect 223666 5284 223672 5296
rect 174228 5256 223672 5284
rect 174228 5244 174234 5256
rect 223666 5244 223672 5256
rect 223724 5244 223730 5296
rect 343542 5244 343548 5296
rect 343600 5284 343606 5296
rect 404906 5284 404912 5296
rect 343600 5256 404912 5284
rect 343600 5244 343606 5256
rect 404906 5244 404912 5256
rect 404964 5244 404970 5296
rect 420822 5244 420828 5296
rect 420880 5284 420886 5296
rect 554774 5284 554780 5296
rect 420880 5256 554780 5284
rect 420880 5244 420886 5256
rect 554774 5244 554780 5256
rect 554832 5244 554838 5296
rect 65978 5176 65984 5228
rect 66036 5216 66042 5228
rect 166994 5216 167000 5228
rect 66036 5188 167000 5216
rect 66036 5176 66042 5188
rect 166994 5176 167000 5188
rect 167052 5176 167058 5228
rect 170582 5176 170588 5228
rect 170640 5216 170646 5228
rect 220998 5216 221004 5228
rect 170640 5188 221004 5216
rect 170640 5176 170646 5188
rect 220998 5176 221004 5188
rect 221056 5176 221062 5228
rect 303522 5176 303528 5228
rect 303580 5216 303586 5228
rect 327626 5216 327632 5228
rect 303580 5188 327632 5216
rect 303580 5176 303586 5188
rect 327626 5176 327632 5188
rect 327684 5176 327690 5228
rect 344922 5176 344928 5228
rect 344980 5216 344986 5228
rect 408494 5216 408500 5228
rect 344980 5188 408500 5216
rect 344980 5176 344986 5188
rect 408494 5176 408500 5188
rect 408552 5176 408558 5228
rect 422202 5176 422208 5228
rect 422260 5216 422266 5228
rect 558362 5216 558368 5228
rect 422260 5188 558368 5216
rect 422260 5176 422266 5188
rect 558362 5176 558368 5188
rect 558420 5176 558426 5228
rect 37366 5108 37372 5160
rect 37424 5148 37430 5160
rect 153378 5148 153384 5160
rect 37424 5120 153384 5148
rect 37424 5108 37430 5120
rect 153378 5108 153384 5120
rect 153436 5108 153442 5160
rect 160002 5108 160008 5160
rect 160060 5148 160066 5160
rect 209866 5148 209872 5160
rect 160060 5120 209872 5148
rect 160060 5108 160066 5120
rect 209866 5108 209872 5120
rect 209924 5108 209930 5160
rect 307662 5108 307668 5160
rect 307720 5148 307726 5160
rect 334710 5148 334716 5160
rect 307720 5120 334716 5148
rect 307720 5108 307726 5120
rect 334710 5108 334716 5120
rect 334768 5108 334774 5160
rect 346302 5108 346308 5160
rect 346360 5148 346366 5160
rect 412082 5148 412088 5160
rect 346360 5120 412088 5148
rect 346360 5108 346366 5120
rect 412082 5108 412088 5120
rect 412140 5108 412146 5160
rect 426342 5108 426348 5160
rect 426400 5148 426406 5160
rect 565538 5148 565544 5160
rect 426400 5120 565544 5148
rect 426400 5108 426406 5120
rect 565538 5108 565544 5120
rect 565596 5108 565602 5160
rect 30282 5040 30288 5092
rect 30340 5080 30346 5092
rect 149054 5080 149060 5092
rect 30340 5052 149060 5080
rect 30340 5040 30346 5052
rect 149054 5040 149060 5052
rect 149112 5040 149118 5092
rect 167086 5040 167092 5092
rect 167144 5080 167150 5092
rect 219526 5080 219532 5092
rect 167144 5052 219532 5080
rect 167144 5040 167150 5052
rect 219526 5040 219532 5052
rect 219584 5040 219590 5092
rect 304902 5040 304908 5092
rect 304960 5080 304966 5092
rect 331214 5080 331220 5092
rect 304960 5052 331220 5080
rect 304960 5040 304966 5052
rect 331214 5040 331220 5052
rect 331272 5040 331278 5092
rect 349062 5040 349068 5092
rect 349120 5080 349126 5092
rect 415670 5080 415676 5092
rect 349120 5052 415676 5080
rect 349120 5040 349126 5052
rect 415670 5040 415676 5052
rect 415728 5040 415734 5092
rect 423490 5040 423496 5092
rect 423548 5080 423554 5092
rect 561950 5080 561956 5092
rect 423548 5052 561956 5080
rect 423548 5040 423554 5052
rect 561950 5040 561956 5052
rect 562008 5040 562014 5092
rect 26694 4972 26700 5024
rect 26752 5012 26758 5024
rect 147766 5012 147772 5024
rect 26752 4984 147772 5012
rect 26752 4972 26758 4984
rect 147766 4972 147772 4984
rect 147824 4972 147830 5024
rect 163498 4972 163504 5024
rect 163556 5012 163562 5024
rect 218054 5012 218060 5024
rect 163556 4984 218060 5012
rect 163556 4972 163562 4984
rect 218054 4972 218060 4984
rect 218112 4972 218118 5024
rect 219342 4972 219348 5024
rect 219400 5012 219406 5024
rect 245746 5012 245752 5024
rect 219400 4984 245752 5012
rect 219400 4972 219406 4984
rect 245746 4972 245752 4984
rect 245804 4972 245810 5024
rect 308950 4972 308956 5024
rect 309008 5012 309014 5024
rect 338298 5012 338304 5024
rect 309008 4984 338304 5012
rect 309008 4972 309014 4984
rect 338298 4972 338304 4984
rect 338356 4972 338362 5024
rect 350442 4972 350448 5024
rect 350500 5012 350506 5024
rect 419166 5012 419172 5024
rect 350500 4984 419172 5012
rect 350500 4972 350506 4984
rect 419166 4972 419172 4984
rect 419224 4972 419230 5024
rect 427722 4972 427728 5024
rect 427780 5012 427786 5024
rect 569034 5012 569040 5024
rect 427780 4984 569040 5012
rect 427780 4972 427786 4984
rect 569034 4972 569040 4984
rect 569092 4972 569098 5024
rect 21910 4904 21916 4956
rect 21968 4944 21974 4956
rect 145006 4944 145012 4956
rect 21968 4916 145012 4944
rect 21968 4904 21974 4916
rect 145006 4904 145012 4916
rect 145064 4904 145070 4956
rect 158714 4904 158720 4956
rect 158772 4944 158778 4956
rect 215294 4944 215300 4956
rect 158772 4916 215300 4944
rect 158772 4904 158778 4916
rect 215294 4904 215300 4916
rect 215352 4904 215358 4956
rect 215846 4904 215852 4956
rect 215904 4944 215910 4956
rect 244550 4944 244556 4956
rect 215904 4916 244556 4944
rect 215904 4904 215910 4916
rect 244550 4904 244556 4916
rect 244608 4904 244614 4956
rect 310422 4904 310428 4956
rect 310480 4944 310486 4956
rect 341886 4944 341892 4956
rect 310480 4916 341892 4944
rect 310480 4904 310486 4916
rect 341886 4904 341892 4916
rect 341944 4904 341950 4956
rect 351822 4904 351828 4956
rect 351880 4944 351886 4956
rect 422754 4944 422760 4956
rect 351880 4916 422760 4944
rect 351880 4904 351886 4916
rect 422754 4904 422760 4916
rect 422812 4904 422818 4956
rect 429102 4904 429108 4956
rect 429160 4944 429166 4956
rect 572622 4944 572628 4956
rect 429160 4916 572628 4944
rect 429160 4904 429166 4916
rect 572622 4904 572628 4916
rect 572680 4904 572686 4956
rect 17218 4836 17224 4888
rect 17276 4876 17282 4888
rect 142246 4876 142252 4888
rect 17276 4848 142252 4876
rect 17276 4836 17282 4848
rect 142246 4836 142252 4848
rect 142304 4836 142310 4888
rect 145650 4836 145656 4888
rect 145708 4876 145714 4888
rect 208394 4876 208400 4888
rect 145708 4848 208400 4876
rect 145708 4836 145714 4848
rect 208394 4836 208400 4848
rect 208452 4836 208458 4888
rect 208670 4836 208676 4888
rect 208728 4876 208734 4888
rect 240134 4876 240140 4888
rect 208728 4848 240140 4876
rect 208728 4836 208734 4848
rect 240134 4836 240140 4848
rect 240192 4836 240198 4888
rect 311802 4836 311808 4888
rect 311860 4876 311866 4888
rect 345474 4876 345480 4888
rect 311860 4848 345480 4876
rect 311860 4836 311866 4848
rect 345474 4836 345480 4848
rect 345532 4836 345538 4888
rect 354582 4836 354588 4888
rect 354640 4876 354646 4888
rect 426342 4876 426348 4888
rect 354640 4848 426348 4876
rect 354640 4836 354646 4848
rect 426342 4836 426348 4848
rect 426400 4836 426406 4888
rect 431862 4836 431868 4888
rect 431920 4876 431926 4888
rect 576210 4876 576216 4888
rect 431920 4848 576216 4876
rect 431920 4836 431926 4848
rect 576210 4836 576216 4848
rect 576268 4836 576274 4888
rect 12434 4768 12440 4820
rect 12492 4808 12498 4820
rect 139486 4808 139492 4820
rect 12492 4780 139492 4808
rect 12492 4768 12498 4780
rect 139486 4768 139492 4780
rect 139544 4768 139550 4820
rect 142062 4768 142068 4820
rect 142120 4808 142126 4820
rect 207014 4808 207020 4820
rect 142120 4780 207020 4808
rect 142120 4768 142126 4780
rect 207014 4768 207020 4780
rect 207072 4768 207078 4820
rect 212258 4768 212264 4820
rect 212316 4808 212322 4820
rect 242986 4808 242992 4820
rect 212316 4780 242992 4808
rect 212316 4768 212322 4780
rect 242986 4768 242992 4780
rect 243044 4768 243050 4820
rect 314562 4768 314568 4820
rect 314620 4808 314626 4820
rect 349062 4808 349068 4820
rect 314620 4780 349068 4808
rect 314620 4768 314626 4780
rect 349062 4768 349068 4780
rect 349120 4768 349126 4820
rect 355962 4768 355968 4820
rect 356020 4808 356026 4820
rect 429930 4808 429936 4820
rect 356020 4780 429936 4808
rect 356020 4768 356026 4780
rect 429930 4768 429936 4780
rect 429988 4768 429994 4820
rect 433242 4768 433248 4820
rect 433300 4808 433306 4820
rect 579798 4808 579804 4820
rect 433300 4780 579804 4808
rect 433300 4768 433306 4780
rect 579798 4768 579804 4780
rect 579856 4768 579862 4820
rect 83826 4700 83832 4752
rect 83884 4740 83890 4752
rect 176746 4740 176752 4752
rect 83884 4712 176752 4740
rect 83884 4700 83890 4712
rect 176746 4700 176752 4712
rect 176804 4700 176810 4752
rect 206922 4700 206928 4752
rect 206980 4740 206986 4752
rect 234706 4740 234712 4752
rect 206980 4712 234712 4740
rect 206980 4700 206986 4712
rect 234706 4700 234712 4712
rect 234764 4700 234770 4752
rect 338022 4700 338028 4752
rect 338080 4740 338086 4752
rect 394234 4740 394240 4752
rect 338080 4712 394240 4740
rect 338080 4700 338086 4712
rect 394234 4700 394240 4712
rect 394292 4700 394298 4752
rect 412542 4700 412548 4752
rect 412600 4740 412606 4752
rect 540514 4740 540520 4752
rect 412600 4712 540520 4740
rect 412600 4700 412606 4712
rect 540514 4700 540520 4712
rect 540572 4700 540578 4752
rect 90910 4632 90916 4684
rect 90968 4672 90974 4684
rect 180886 4672 180892 4684
rect 90968 4644 180892 4672
rect 90968 4632 90974 4644
rect 180886 4632 180892 4644
rect 180944 4632 180950 4684
rect 204346 4632 204352 4684
rect 204404 4672 204410 4684
rect 233510 4672 233516 4684
rect 204404 4644 233516 4672
rect 204404 4632 204410 4644
rect 233510 4632 233516 4644
rect 233568 4632 233574 4684
rect 333790 4632 333796 4684
rect 333848 4672 333854 4684
rect 387058 4672 387064 4684
rect 333848 4644 387064 4672
rect 333848 4632 333854 4644
rect 387058 4632 387064 4644
rect 387116 4632 387122 4684
rect 411162 4632 411168 4684
rect 411220 4672 411226 4684
rect 536926 4672 536932 4684
rect 411220 4644 536932 4672
rect 411220 4632 411226 4644
rect 536926 4632 536932 4644
rect 536984 4632 536990 4684
rect 87322 4564 87328 4616
rect 87380 4604 87386 4616
rect 178034 4604 178040 4616
rect 87380 4576 178040 4604
rect 87380 4564 87386 4576
rect 178034 4564 178040 4576
rect 178092 4564 178098 4616
rect 204254 4564 204260 4616
rect 204312 4604 204318 4616
rect 231946 4604 231952 4616
rect 204312 4576 231952 4604
rect 204312 4564 204318 4576
rect 231946 4564 231952 4576
rect 232004 4564 232010 4616
rect 329650 4564 329656 4616
rect 329708 4604 329714 4616
rect 379974 4604 379980 4616
rect 329708 4576 379980 4604
rect 329708 4564 329714 4576
rect 379974 4564 379980 4576
rect 380032 4564 380038 4616
rect 409782 4564 409788 4616
rect 409840 4604 409846 4616
rect 533430 4604 533436 4616
rect 409840 4576 533436 4604
rect 409840 4564 409846 4576
rect 533430 4564 533436 4576
rect 533488 4564 533494 4616
rect 49326 4496 49332 4548
rect 49384 4536 49390 4548
rect 130470 4536 130476 4548
rect 49384 4508 130476 4536
rect 49384 4496 49390 4508
rect 130470 4496 130476 4508
rect 130528 4496 130534 4548
rect 162118 4496 162124 4548
rect 162176 4536 162182 4548
rect 208486 4536 208492 4548
rect 162176 4508 208492 4536
rect 162176 4496 162182 4508
rect 208486 4496 208492 4508
rect 208544 4496 208550 4548
rect 332502 4496 332508 4548
rect 332560 4536 332566 4548
rect 383562 4536 383568 4548
rect 332560 4508 383568 4536
rect 332560 4496 332566 4508
rect 383562 4496 383568 4508
rect 383620 4496 383626 4548
rect 406930 4496 406936 4548
rect 406988 4536 406994 4548
rect 529842 4536 529848 4548
rect 406988 4508 529848 4536
rect 406988 4496 406994 4508
rect 529842 4496 529848 4508
rect 529900 4496 529906 4548
rect 52822 4428 52828 4480
rect 52880 4468 52886 4480
rect 122098 4468 122104 4480
rect 52880 4440 122104 4468
rect 52880 4428 52886 4440
rect 122098 4428 122104 4440
rect 122156 4428 122162 4480
rect 202966 4428 202972 4480
rect 203024 4468 203030 4480
rect 229186 4468 229192 4480
rect 203024 4440 229192 4468
rect 203024 4428 203030 4440
rect 229186 4428 229192 4440
rect 229244 4428 229250 4480
rect 328362 4428 328368 4480
rect 328420 4468 328426 4480
rect 376386 4468 376392 4480
rect 328420 4440 376392 4468
rect 328420 4428 328426 4440
rect 376386 4428 376392 4440
rect 376444 4428 376450 4480
rect 405642 4428 405648 4480
rect 405700 4468 405706 4480
rect 526254 4468 526260 4480
rect 405700 4440 526260 4468
rect 405700 4428 405706 4440
rect 526254 4428 526260 4440
rect 526312 4428 526318 4480
rect 70670 4360 70676 4412
rect 70728 4400 70734 4412
rect 120718 4400 120724 4412
rect 70728 4372 120724 4400
rect 70728 4360 70734 4372
rect 120718 4360 120724 4372
rect 120776 4360 120782 4412
rect 120810 4360 120816 4412
rect 120868 4400 120874 4412
rect 146386 4400 146392 4412
rect 120868 4372 146392 4400
rect 120868 4360 120874 4372
rect 146386 4360 146392 4372
rect 146444 4360 146450 4412
rect 202874 4360 202880 4412
rect 202932 4400 202938 4412
rect 227990 4400 227996 4412
rect 202932 4372 227996 4400
rect 202932 4360 202938 4372
rect 227990 4360 227996 4372
rect 228048 4360 228054 4412
rect 326982 4360 326988 4412
rect 327040 4400 327046 4412
rect 372798 4400 372804 4412
rect 327040 4372 372804 4400
rect 327040 4360 327046 4372
rect 372798 4360 372804 4372
rect 372856 4360 372862 4412
rect 404262 4360 404268 4412
rect 404320 4400 404326 4412
rect 522666 4400 522672 4412
rect 404320 4372 522672 4400
rect 404320 4360 404326 4372
rect 522666 4360 522672 4372
rect 522724 4360 522730 4412
rect 324130 4292 324136 4344
rect 324188 4332 324194 4344
rect 369210 4332 369216 4344
rect 324188 4304 369216 4332
rect 324188 4292 324194 4304
rect 369210 4292 369216 4304
rect 369268 4292 369274 4344
rect 401502 4292 401508 4344
rect 401560 4332 401566 4344
rect 519078 4332 519084 4344
rect 401560 4304 519084 4332
rect 401560 4292 401566 4304
rect 519078 4292 519084 4304
rect 519136 4292 519142 4344
rect 322842 4224 322848 4276
rect 322900 4264 322906 4276
rect 365714 4264 365720 4276
rect 322900 4236 365720 4264
rect 322900 4224 322906 4236
rect 365714 4224 365720 4236
rect 365772 4224 365778 4276
rect 400122 4224 400128 4276
rect 400180 4264 400186 4276
rect 515582 4264 515588 4276
rect 400180 4236 515588 4264
rect 400180 4224 400186 4236
rect 515582 4224 515588 4236
rect 515640 4224 515646 4276
rect 25498 4088 25504 4140
rect 25556 4128 25562 4140
rect 120810 4128 120816 4140
rect 25556 4100 120816 4128
rect 25556 4088 25562 4100
rect 120810 4088 120816 4100
rect 120868 4088 120874 4140
rect 125410 4088 125416 4140
rect 125468 4128 125474 4140
rect 170398 4128 170404 4140
rect 125468 4100 170404 4128
rect 125468 4088 125474 4100
rect 170398 4088 170404 4100
rect 170456 4088 170462 4140
rect 175366 4088 175372 4140
rect 175424 4128 175430 4140
rect 176562 4128 176568 4140
rect 175424 4100 176568 4128
rect 175424 4088 175430 4100
rect 176562 4088 176568 4100
rect 176620 4088 176626 4140
rect 181346 4088 181352 4140
rect 181404 4128 181410 4140
rect 182082 4128 182088 4140
rect 181404 4100 182088 4128
rect 181404 4088 181410 4100
rect 182082 4088 182088 4100
rect 182140 4088 182146 4140
rect 182542 4088 182548 4140
rect 182600 4128 182606 4140
rect 183462 4128 183468 4140
rect 182600 4100 183468 4128
rect 182600 4088 182606 4100
rect 183462 4088 183468 4100
rect 183520 4088 183526 4140
rect 188430 4088 188436 4140
rect 188488 4128 188494 4140
rect 188982 4128 188988 4140
rect 188488 4100 188988 4128
rect 188488 4088 188494 4100
rect 188982 4088 188988 4100
rect 189040 4088 189046 4140
rect 196802 4088 196808 4140
rect 196860 4128 196866 4140
rect 197262 4128 197268 4140
rect 196860 4100 197268 4128
rect 196860 4088 196866 4100
rect 197262 4088 197268 4100
rect 197320 4088 197326 4140
rect 199194 4088 199200 4140
rect 199252 4128 199258 4140
rect 200022 4128 200028 4140
rect 199252 4100 200028 4128
rect 199252 4088 199258 4100
rect 200022 4088 200028 4100
rect 200080 4088 200086 4140
rect 203886 4088 203892 4140
rect 203944 4128 203950 4140
rect 229738 4128 229744 4140
rect 203944 4100 229744 4128
rect 203944 4088 203950 4100
rect 229738 4088 229744 4100
rect 229796 4088 229802 4140
rect 231302 4088 231308 4140
rect 231360 4128 231366 4140
rect 231762 4128 231768 4140
rect 231360 4100 231768 4128
rect 231360 4088 231366 4100
rect 231762 4088 231768 4100
rect 231820 4088 231826 4140
rect 232498 4088 232504 4140
rect 232556 4128 232562 4140
rect 233142 4128 233148 4140
rect 232556 4100 233148 4128
rect 232556 4088 232562 4100
rect 233142 4088 233148 4100
rect 233200 4088 233206 4140
rect 233694 4088 233700 4140
rect 233752 4128 233758 4140
rect 234522 4128 234528 4140
rect 233752 4100 234528 4128
rect 233752 4088 233758 4100
rect 234522 4088 234528 4100
rect 234580 4088 234586 4140
rect 234798 4088 234804 4140
rect 234856 4128 234862 4140
rect 235902 4128 235908 4140
rect 234856 4100 235908 4128
rect 234856 4088 234862 4100
rect 235902 4088 235908 4100
rect 235960 4088 235966 4140
rect 235994 4088 236000 4140
rect 236052 4128 236058 4140
rect 237282 4128 237288 4140
rect 236052 4100 237288 4128
rect 236052 4088 236058 4100
rect 237282 4088 237288 4100
rect 237340 4088 237346 4140
rect 239582 4088 239588 4140
rect 239640 4128 239646 4140
rect 240042 4128 240048 4140
rect 239640 4100 240048 4128
rect 239640 4088 239646 4100
rect 240042 4088 240048 4100
rect 240100 4088 240106 4140
rect 240778 4088 240784 4140
rect 240836 4128 240842 4140
rect 241422 4128 241428 4140
rect 240836 4100 241428 4128
rect 240836 4088 240842 4100
rect 241422 4088 241428 4100
rect 241480 4088 241486 4140
rect 243170 4088 243176 4140
rect 243228 4128 243234 4140
rect 244182 4128 244188 4140
rect 243228 4100 244188 4128
rect 243228 4088 243234 4100
rect 244182 4088 244188 4100
rect 244240 4088 244246 4140
rect 244366 4088 244372 4140
rect 244424 4128 244430 4140
rect 245562 4128 245568 4140
rect 244424 4100 245568 4128
rect 244424 4088 244430 4100
rect 245562 4088 245568 4100
rect 245620 4088 245626 4140
rect 249150 4088 249156 4140
rect 249208 4128 249214 4140
rect 249702 4128 249708 4140
rect 249208 4100 249708 4128
rect 249208 4088 249214 4100
rect 249702 4088 249708 4100
rect 249760 4088 249766 4140
rect 251450 4088 251456 4140
rect 251508 4128 251514 4140
rect 252462 4128 252468 4140
rect 251508 4100 252468 4128
rect 251508 4088 251514 4100
rect 252462 4088 252468 4100
rect 252520 4088 252526 4140
rect 252646 4088 252652 4140
rect 252704 4128 252710 4140
rect 253842 4128 253848 4140
rect 252704 4100 253848 4128
rect 252704 4088 252710 4100
rect 253842 4088 253848 4100
rect 253900 4088 253906 4140
rect 274082 4088 274088 4140
rect 274140 4128 274146 4140
rect 274542 4128 274548 4140
rect 274140 4100 274548 4128
rect 274140 4088 274146 4100
rect 274542 4088 274548 4100
rect 274600 4088 274606 4140
rect 277302 4088 277308 4140
rect 277360 4128 277366 4140
rect 277670 4128 277676 4140
rect 277360 4100 277676 4128
rect 277360 4088 277366 4100
rect 277670 4088 277676 4100
rect 277728 4088 277734 4140
rect 278590 4088 278596 4140
rect 278648 4128 278654 4140
rect 280062 4128 280068 4140
rect 278648 4100 280068 4128
rect 278648 4088 278654 4100
rect 280062 4088 280068 4100
rect 280120 4088 280126 4140
rect 284110 4088 284116 4140
rect 284168 4128 284174 4140
rect 289538 4128 289544 4140
rect 284168 4100 289544 4128
rect 284168 4088 284174 4100
rect 289538 4088 289544 4100
rect 289596 4088 289602 4140
rect 289722 4088 289728 4140
rect 289780 4128 289786 4140
rect 301406 4128 301412 4140
rect 289780 4100 301412 4128
rect 289780 4088 289786 4100
rect 301406 4088 301412 4100
rect 301464 4088 301470 4140
rect 312538 4088 312544 4140
rect 312596 4128 312602 4140
rect 314562 4128 314568 4140
rect 312596 4100 314568 4128
rect 312596 4088 312602 4100
rect 314562 4088 314568 4100
rect 314620 4088 314626 4140
rect 324222 4088 324228 4140
rect 324280 4128 324286 4140
rect 368014 4128 368020 4140
rect 324280 4100 368020 4128
rect 324280 4088 324286 4100
rect 368014 4088 368020 4100
rect 368072 4088 368078 4140
rect 379422 4088 379428 4140
rect 379480 4128 379486 4140
rect 475102 4128 475108 4140
rect 379480 4100 475108 4128
rect 379480 4088 379486 4100
rect 475102 4088 475108 4100
rect 475160 4088 475166 4140
rect 477494 4088 477500 4140
rect 477552 4128 477558 4140
rect 478690 4128 478696 4140
rect 477552 4100 478696 4128
rect 477552 4088 477558 4100
rect 478690 4088 478696 4100
rect 478748 4088 478754 4140
rect 480898 4088 480904 4140
rect 480956 4128 480962 4140
rect 481266 4128 481272 4140
rect 480956 4100 481272 4128
rect 480956 4088 480962 4100
rect 481266 4088 481272 4100
rect 481324 4088 481330 4140
rect 489178 4088 489184 4140
rect 489236 4128 489242 4140
rect 489546 4128 489552 4140
rect 489236 4100 489552 4128
rect 489236 4088 489242 4100
rect 489546 4088 489552 4100
rect 489604 4088 489610 4140
rect 496078 4088 496084 4140
rect 496136 4128 496142 4140
rect 503530 4128 503536 4140
rect 496136 4100 503536 4128
rect 496136 4088 496142 4100
rect 503530 4088 503536 4100
rect 503588 4088 503594 4140
rect 503806 4088 503812 4140
rect 503864 4128 503870 4140
rect 571426 4128 571432 4140
rect 503864 4100 571432 4128
rect 503864 4088 503870 4100
rect 571426 4088 571432 4100
rect 571484 4088 571490 4140
rect 42150 4020 42156 4072
rect 42208 4060 42214 4072
rect 42702 4060 42708 4072
rect 42208 4032 42708 4060
rect 42208 4020 42214 4032
rect 42702 4020 42708 4032
rect 42760 4020 42766 4072
rect 43346 4020 43352 4072
rect 43404 4060 43410 4072
rect 155954 4060 155960 4072
rect 43404 4032 155960 4060
rect 43404 4020 43410 4032
rect 155954 4020 155960 4032
rect 156012 4020 156018 4072
rect 164694 4020 164700 4072
rect 164752 4060 164758 4072
rect 188614 4060 188620 4072
rect 164752 4032 188620 4060
rect 164752 4020 164758 4032
rect 188614 4020 188620 4032
rect 188672 4020 188678 4072
rect 189626 4020 189632 4072
rect 189684 4060 189690 4072
rect 225598 4060 225604 4072
rect 189684 4032 225604 4060
rect 189684 4020 189690 4032
rect 225598 4020 225604 4032
rect 225656 4020 225662 4072
rect 253658 4020 253664 4072
rect 253716 4060 253722 4072
rect 253716 4032 253888 4060
rect 253716 4020 253722 4032
rect 253860 4004 253888 4032
rect 279970 4020 279976 4072
rect 280028 4060 280034 4072
rect 282454 4060 282460 4072
rect 280028 4032 282460 4060
rect 280028 4020 280034 4032
rect 282454 4020 282460 4032
rect 282512 4020 282518 4072
rect 291102 4020 291108 4072
rect 291160 4060 291166 4072
rect 303798 4060 303804 4072
rect 291160 4032 303804 4060
rect 291160 4020 291166 4032
rect 303798 4020 303804 4032
rect 303856 4020 303862 4072
rect 325602 4020 325608 4072
rect 325660 4060 325666 4072
rect 371602 4060 371608 4072
rect 325660 4032 371608 4060
rect 325660 4020 325666 4032
rect 371602 4020 371608 4032
rect 371660 4020 371666 4072
rect 383470 4020 383476 4072
rect 383528 4060 383534 4072
rect 482278 4060 482284 4072
rect 383528 4032 482284 4060
rect 383528 4020 383534 4032
rect 482278 4020 482284 4032
rect 482336 4020 482342 4072
rect 500218 4020 500224 4072
rect 500276 4060 500282 4072
rect 578602 4060 578608 4072
rect 500276 4032 578608 4060
rect 500276 4020 500282 4032
rect 578602 4020 578608 4032
rect 578660 4020 578666 4072
rect 36170 3952 36176 4004
rect 36228 3992 36234 4004
rect 151906 3992 151912 4004
rect 36228 3964 151912 3992
rect 36228 3952 36234 3964
rect 151906 3952 151912 3964
rect 151964 3952 151970 4004
rect 156322 3952 156328 4004
rect 156380 3992 156386 4004
rect 194594 3992 194600 4004
rect 156380 3964 194600 3992
rect 156380 3952 156386 3964
rect 194594 3952 194600 3964
rect 194652 3952 194658 4004
rect 209866 3952 209872 4004
rect 209924 3992 209930 4004
rect 238110 3992 238116 4004
rect 209924 3964 238116 3992
rect 209924 3952 209930 3964
rect 238110 3952 238116 3964
rect 238168 3952 238174 4004
rect 253842 3952 253848 4004
rect 253900 3952 253906 4004
rect 286962 3952 286968 4004
rect 287020 3992 287026 4004
rect 295518 3992 295524 4004
rect 287020 3964 295524 3992
rect 287020 3952 287026 3964
rect 295518 3952 295524 3964
rect 295576 3952 295582 4004
rect 297910 3952 297916 4004
rect 297968 3992 297974 4004
rect 316954 3992 316960 4004
rect 297968 3964 316960 3992
rect 297968 3952 297974 3964
rect 316954 3952 316960 3964
rect 317012 3952 317018 4004
rect 329742 3952 329748 4004
rect 329800 3992 329806 4004
rect 378778 3992 378784 4004
rect 329800 3964 378784 3992
rect 329800 3952 329806 3964
rect 378778 3952 378784 3964
rect 378836 3952 378842 4004
rect 521470 3992 521476 4004
rect 403912 3964 521476 3992
rect 29086 3884 29092 3936
rect 29144 3924 29150 3936
rect 147950 3924 147956 3936
rect 29144 3896 147956 3924
rect 29144 3884 29150 3896
rect 147950 3884 147956 3896
rect 148008 3884 148014 3936
rect 152734 3884 152740 3936
rect 152792 3924 152798 3936
rect 197170 3924 197176 3936
rect 152792 3896 197176 3924
rect 152792 3884 152798 3896
rect 197170 3884 197176 3896
rect 197228 3884 197234 3936
rect 202690 3884 202696 3936
rect 202748 3924 202754 3936
rect 231118 3924 231124 3936
rect 202748 3896 231124 3924
rect 202748 3884 202754 3896
rect 231118 3884 231124 3896
rect 231176 3884 231182 3936
rect 293862 3884 293868 3936
rect 293920 3924 293926 3936
rect 309778 3924 309784 3936
rect 293920 3896 309784 3924
rect 293920 3884 293926 3896
rect 309778 3884 309784 3896
rect 309836 3884 309842 3936
rect 312630 3884 312636 3936
rect 312688 3924 312694 3936
rect 332410 3924 332416 3936
rect 312688 3896 332416 3924
rect 312688 3884 312694 3896
rect 332410 3884 332416 3896
rect 332468 3884 332474 3936
rect 338758 3884 338764 3936
rect 338816 3924 338822 3936
rect 389450 3924 389456 3936
rect 338816 3896 389456 3924
rect 338816 3884 338822 3896
rect 389450 3884 389456 3896
rect 389508 3884 389514 3936
rect 402882 3884 402888 3936
rect 402940 3924 402946 3936
rect 403912 3924 403940 3964
rect 521470 3952 521476 3964
rect 521528 3952 521534 4004
rect 402940 3896 403940 3924
rect 402940 3884 402946 3896
rect 407022 3884 407028 3936
rect 407080 3924 407086 3936
rect 528646 3924 528652 3936
rect 407080 3896 528652 3924
rect 407080 3884 407086 3896
rect 528646 3884 528652 3896
rect 528704 3884 528710 3936
rect 24302 3816 24308 3868
rect 24360 3856 24366 3868
rect 146294 3856 146300 3868
rect 24360 3828 146300 3856
rect 24360 3816 24366 3828
rect 146294 3816 146300 3828
rect 146352 3816 146358 3868
rect 151538 3816 151544 3868
rect 151596 3856 151602 3868
rect 196618 3856 196624 3868
rect 151596 3828 196624 3856
rect 151596 3816 151602 3828
rect 196618 3816 196624 3828
rect 196676 3816 196682 3868
rect 197998 3816 198004 3868
rect 198056 3856 198062 3868
rect 206922 3856 206928 3868
rect 198056 3828 206928 3856
rect 198056 3816 198062 3828
rect 206922 3816 206928 3828
rect 206980 3816 206986 3868
rect 211062 3816 211068 3868
rect 211120 3856 211126 3868
rect 239398 3856 239404 3868
rect 211120 3828 239404 3856
rect 211120 3816 211126 3828
rect 239398 3816 239404 3828
rect 239456 3816 239462 3868
rect 285582 3816 285588 3868
rect 285640 3856 285646 3868
rect 293126 3856 293132 3868
rect 285640 3828 293132 3856
rect 285640 3816 285646 3828
rect 293126 3816 293132 3828
rect 293184 3816 293190 3868
rect 295242 3816 295248 3868
rect 295300 3856 295306 3868
rect 310974 3856 310980 3868
rect 295300 3828 310980 3856
rect 295300 3816 295306 3828
rect 310974 3816 310980 3828
rect 311032 3816 311038 3868
rect 313918 3816 313924 3868
rect 313976 3856 313982 3868
rect 335906 3856 335912 3868
rect 313976 3828 335912 3856
rect 313976 3816 313982 3828
rect 335906 3816 335912 3828
rect 335964 3816 335970 3868
rect 341702 3816 341708 3868
rect 341760 3856 341766 3868
rect 393038 3856 393044 3868
rect 341760 3828 393044 3856
rect 341760 3816 341766 3828
rect 393038 3816 393044 3828
rect 393096 3816 393102 3868
rect 409506 3816 409512 3868
rect 409564 3856 409570 3868
rect 535730 3856 535736 3868
rect 409564 3828 535736 3856
rect 409564 3816 409570 3828
rect 535730 3816 535736 3828
rect 535788 3816 535794 3868
rect 20714 3748 20720 3800
rect 20772 3788 20778 3800
rect 143718 3788 143724 3800
rect 20772 3760 143724 3788
rect 20772 3748 20778 3760
rect 143718 3748 143724 3760
rect 143776 3748 143782 3800
rect 172974 3748 172980 3800
rect 173032 3788 173038 3800
rect 180058 3788 180064 3800
rect 173032 3760 180064 3788
rect 173032 3748 173038 3760
rect 180058 3748 180064 3760
rect 180116 3748 180122 3800
rect 180150 3748 180156 3800
rect 180208 3788 180214 3800
rect 222102 3788 222108 3800
rect 180208 3760 222108 3788
rect 180208 3748 180214 3760
rect 222102 3748 222108 3760
rect 222160 3748 222166 3800
rect 222838 3748 222844 3800
rect 222896 3788 222902 3800
rect 226426 3788 226432 3800
rect 222896 3760 226432 3788
rect 222896 3748 222902 3760
rect 226426 3748 226432 3760
rect 226484 3748 226490 3800
rect 228910 3748 228916 3800
rect 228968 3788 228974 3800
rect 228968 3760 229324 3788
rect 228968 3748 228974 3760
rect 19518 3680 19524 3732
rect 19576 3720 19582 3732
rect 143534 3720 143540 3732
rect 19576 3692 143540 3720
rect 19576 3680 19582 3692
rect 143534 3680 143540 3692
rect 143592 3680 143598 3732
rect 155126 3680 155132 3732
rect 155184 3720 155190 3732
rect 173894 3720 173900 3732
rect 155184 3692 173900 3720
rect 155184 3680 155190 3692
rect 173894 3680 173900 3692
rect 173952 3680 173958 3732
rect 176746 3680 176752 3732
rect 176804 3720 176810 3732
rect 223758 3720 223764 3732
rect 176804 3692 223764 3720
rect 176804 3680 176810 3692
rect 223758 3680 223764 3692
rect 223816 3680 223822 3732
rect 226518 3680 226524 3732
rect 226576 3720 226582 3732
rect 226576 3692 229232 3720
rect 226576 3680 226582 3692
rect 14826 3612 14832 3664
rect 14884 3652 14890 3664
rect 140958 3652 140964 3664
rect 14884 3624 140964 3652
rect 14884 3612 14890 3624
rect 140958 3612 140964 3624
rect 141016 3612 141022 3664
rect 186222 3612 186228 3664
rect 186280 3652 186286 3664
rect 222194 3652 222200 3664
rect 186280 3624 222200 3652
rect 186280 3612 186286 3624
rect 222194 3612 222200 3624
rect 222252 3612 222258 3664
rect 227714 3612 227720 3664
rect 227772 3652 227778 3664
rect 229002 3652 229008 3664
rect 227772 3624 229008 3652
rect 227772 3612 227778 3624
rect 229002 3612 229008 3624
rect 229060 3612 229066 3664
rect 16022 3544 16028 3596
rect 16080 3584 16086 3596
rect 142338 3584 142344 3596
rect 16080 3556 142344 3584
rect 16080 3544 16086 3556
rect 142338 3544 142344 3556
rect 142396 3544 142402 3596
rect 169386 3544 169392 3596
rect 169444 3584 169450 3596
rect 220814 3584 220820 3596
rect 169444 3556 220820 3584
rect 169444 3544 169450 3556
rect 220814 3544 220820 3556
rect 220872 3544 220878 3596
rect 229204 3584 229232 3692
rect 229296 3652 229324 3760
rect 288250 3748 288256 3800
rect 288308 3788 288314 3800
rect 299106 3788 299112 3800
rect 288308 3760 299112 3788
rect 288308 3748 288314 3760
rect 299106 3748 299112 3760
rect 299164 3748 299170 3800
rect 302878 3748 302884 3800
rect 302936 3788 302942 3800
rect 302936 3760 308168 3788
rect 302936 3748 302942 3760
rect 230106 3680 230112 3732
rect 230164 3720 230170 3732
rect 251174 3720 251180 3732
rect 230164 3692 251180 3720
rect 230164 3680 230170 3692
rect 251174 3680 251180 3692
rect 251232 3680 251238 3732
rect 291010 3680 291016 3732
rect 291068 3720 291074 3732
rect 302602 3720 302608 3732
rect 291068 3692 302608 3720
rect 291068 3680 291074 3692
rect 302602 3680 302608 3692
rect 302660 3680 302666 3732
rect 306190 3720 306196 3732
rect 302712 3692 306196 3720
rect 250438 3652 250444 3664
rect 229296 3624 250444 3652
rect 250438 3612 250444 3624
rect 250496 3612 250502 3664
rect 284202 3612 284208 3664
rect 284260 3652 284266 3664
rect 290734 3652 290740 3664
rect 284260 3624 290740 3652
rect 284260 3612 284266 3624
rect 290734 3612 290740 3624
rect 290792 3612 290798 3664
rect 292390 3612 292396 3664
rect 292448 3652 292454 3664
rect 302712 3652 302740 3692
rect 306190 3680 306196 3692
rect 306248 3680 306254 3732
rect 308140 3720 308168 3760
rect 309594 3748 309600 3800
rect 309652 3788 309658 3800
rect 321646 3788 321652 3800
rect 309652 3760 321652 3788
rect 309652 3748 309658 3760
rect 321646 3748 321652 3760
rect 321704 3748 321710 3800
rect 333882 3748 333888 3800
rect 333940 3788 333946 3800
rect 385862 3788 385868 3800
rect 333940 3760 385868 3788
rect 333940 3748 333946 3760
rect 385862 3748 385868 3760
rect 385920 3748 385926 3800
rect 414658 3748 414664 3800
rect 414716 3788 414722 3800
rect 542906 3788 542912 3800
rect 414716 3760 542912 3788
rect 414716 3748 414722 3760
rect 542906 3748 542912 3760
rect 542964 3748 542970 3800
rect 325234 3720 325240 3732
rect 308140 3692 325240 3720
rect 325234 3680 325240 3692
rect 325292 3680 325298 3732
rect 342898 3680 342904 3732
rect 342956 3720 342962 3732
rect 400214 3720 400220 3732
rect 342956 3692 400220 3720
rect 342956 3680 342962 3692
rect 400214 3680 400220 3692
rect 400272 3680 400278 3732
rect 420178 3680 420184 3732
rect 420236 3720 420242 3732
rect 553578 3720 553584 3732
rect 420236 3692 553584 3720
rect 420236 3680 420242 3692
rect 553578 3680 553584 3692
rect 553636 3680 553642 3732
rect 292448 3624 302740 3652
rect 292448 3612 292454 3624
rect 305638 3612 305644 3664
rect 305696 3652 305702 3664
rect 328822 3652 328828 3664
rect 305696 3624 328828 3652
rect 305696 3612 305702 3624
rect 328822 3612 328828 3624
rect 328880 3612 328886 3664
rect 345658 3612 345664 3664
rect 345716 3652 345722 3664
rect 407298 3652 407304 3664
rect 345716 3624 407304 3652
rect 345716 3612 345722 3624
rect 407298 3612 407304 3624
rect 407356 3612 407362 3664
rect 407758 3612 407764 3664
rect 407816 3652 407822 3664
rect 410886 3652 410892 3664
rect 407816 3624 410892 3652
rect 407816 3612 407822 3624
rect 410886 3612 410892 3624
rect 410944 3612 410950 3664
rect 423582 3612 423588 3664
rect 423640 3652 423646 3664
rect 560754 3652 560760 3664
rect 423640 3624 560760 3652
rect 423640 3612 423646 3624
rect 560754 3612 560760 3624
rect 560812 3612 560818 3664
rect 250070 3584 250076 3596
rect 229204 3556 250076 3584
rect 250070 3544 250076 3556
rect 250128 3544 250134 3596
rect 279786 3544 279792 3596
rect 279844 3584 279850 3596
rect 283650 3584 283656 3596
rect 279844 3556 283656 3584
rect 279844 3544 279850 3556
rect 283650 3544 283656 3556
rect 283708 3544 283714 3596
rect 286870 3544 286876 3596
rect 286928 3584 286934 3596
rect 296714 3584 296720 3596
rect 286928 3556 296720 3584
rect 286928 3544 286934 3556
rect 296714 3544 296720 3556
rect 296772 3544 296778 3596
rect 298002 3544 298008 3596
rect 298060 3584 298066 3596
rect 318058 3584 318064 3596
rect 298060 3556 318064 3584
rect 298060 3544 298066 3556
rect 318058 3544 318064 3556
rect 318116 3544 318122 3596
rect 318702 3544 318708 3596
rect 318760 3584 318766 3596
rect 357342 3584 357348 3596
rect 318760 3556 357348 3584
rect 318760 3544 318766 3556
rect 357342 3544 357348 3556
rect 357400 3544 357406 3596
rect 358078 3544 358084 3596
rect 358136 3584 358142 3596
rect 364518 3584 364524 3596
rect 358136 3556 364524 3584
rect 358136 3544 358142 3556
rect 364518 3544 364524 3556
rect 364576 3544 364582 3596
rect 364978 3544 364984 3596
rect 365036 3584 365042 3596
rect 428734 3584 428740 3596
rect 365036 3556 428740 3584
rect 365036 3544 365042 3556
rect 428734 3544 428740 3556
rect 428792 3544 428798 3596
rect 429838 3544 429844 3596
rect 429896 3584 429902 3596
rect 567838 3584 567844 3596
rect 429896 3556 567844 3584
rect 429896 3544 429902 3556
rect 567838 3544 567844 3556
rect 567896 3544 567902 3596
rect 8846 3476 8852 3528
rect 8904 3516 8910 3528
rect 9582 3516 9588 3528
rect 8904 3488 9588 3516
rect 8904 3476 8910 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 138014 3516 138020 3528
rect 10100 3488 138020 3516
rect 10100 3476 10106 3488
rect 138014 3476 138020 3488
rect 138072 3476 138078 3528
rect 146846 3476 146852 3528
rect 146904 3516 146910 3528
rect 162118 3516 162124 3528
rect 146904 3488 162124 3516
rect 146904 3476 146910 3488
rect 162118 3476 162124 3488
rect 162176 3476 162182 3528
rect 165890 3476 165896 3528
rect 165948 3516 165954 3528
rect 219434 3516 219440 3528
rect 165948 3488 219440 3516
rect 165948 3476 165954 3488
rect 219434 3476 219440 3488
rect 219492 3476 219498 3528
rect 222102 3476 222108 3528
rect 222160 3516 222166 3528
rect 222838 3516 222844 3528
rect 222160 3488 222844 3516
rect 222160 3476 222166 3488
rect 222838 3476 222844 3488
rect 222896 3476 222902 3528
rect 222930 3476 222936 3528
rect 222988 3516 222994 3528
rect 248506 3516 248512 3528
rect 222988 3488 248512 3516
rect 222988 3476 222994 3488
rect 248506 3476 248512 3488
rect 248564 3476 248570 3528
rect 257430 3476 257436 3528
rect 257488 3516 257494 3528
rect 257982 3516 257988 3528
rect 257488 3488 257988 3516
rect 257488 3476 257494 3488
rect 257982 3476 257988 3488
rect 258040 3476 258046 3528
rect 259822 3476 259828 3528
rect 259880 3516 259886 3528
rect 260742 3516 260748 3528
rect 259880 3488 260748 3516
rect 259880 3476 259886 3488
rect 260742 3476 260748 3488
rect 260800 3476 260806 3528
rect 262214 3476 262220 3528
rect 262272 3516 262278 3528
rect 263502 3516 263508 3528
rect 262272 3488 263508 3516
rect 262272 3476 262278 3488
rect 263502 3476 263508 3488
rect 263560 3476 263566 3528
rect 265802 3476 265808 3528
rect 265860 3516 265866 3528
rect 266262 3516 266268 3528
rect 265860 3488 266268 3516
rect 265860 3476 265866 3488
rect 266262 3476 266268 3488
rect 266320 3476 266326 3528
rect 268102 3476 268108 3528
rect 268160 3516 268166 3528
rect 269022 3516 269028 3528
rect 268160 3488 269028 3516
rect 268160 3476 268166 3488
rect 269022 3476 269028 3488
rect 269080 3476 269086 3528
rect 271690 3476 271696 3528
rect 271748 3516 271754 3528
rect 272518 3516 272524 3528
rect 271748 3488 272524 3516
rect 271748 3476 271754 3488
rect 272518 3476 272524 3488
rect 272576 3476 272582 3528
rect 281442 3476 281448 3528
rect 281500 3516 281506 3528
rect 284754 3516 284760 3528
rect 281500 3488 284760 3516
rect 281500 3476 281506 3488
rect 284754 3476 284760 3488
rect 284812 3476 284818 3528
rect 285398 3476 285404 3528
rect 285456 3516 285462 3528
rect 294322 3516 294328 3528
rect 285456 3488 294328 3516
rect 285456 3476 285462 3488
rect 294322 3476 294328 3488
rect 294380 3476 294386 3528
rect 296622 3476 296628 3528
rect 296680 3516 296686 3528
rect 296680 3488 308628 3516
rect 296680 3476 296686 3488
rect 11238 3408 11244 3460
rect 11296 3448 11302 3460
rect 139578 3448 139584 3460
rect 11296 3420 139584 3448
rect 11296 3408 11302 3420
rect 139578 3408 139584 3420
rect 139636 3408 139642 3460
rect 149238 3408 149244 3460
rect 149296 3448 149302 3460
rect 160002 3448 160008 3460
rect 149296 3420 160008 3448
rect 149296 3408 149302 3420
rect 160002 3408 160008 3420
rect 160060 3408 160066 3460
rect 162302 3408 162308 3460
rect 162360 3448 162366 3460
rect 216950 3448 216956 3460
rect 162360 3420 216956 3448
rect 162360 3408 162366 3420
rect 216950 3408 216956 3420
rect 217008 3408 217014 3460
rect 218146 3408 218152 3460
rect 218204 3448 218210 3460
rect 245838 3448 245844 3460
rect 218204 3420 245844 3448
rect 218204 3408 218210 3420
rect 245838 3408 245844 3420
rect 245896 3408 245902 3460
rect 266998 3408 267004 3460
rect 267056 3448 267062 3460
rect 267642 3448 267648 3460
rect 267056 3420 267648 3448
rect 267056 3408 267062 3420
rect 267642 3408 267648 3420
rect 267700 3408 267706 3460
rect 270494 3408 270500 3460
rect 270552 3448 270558 3460
rect 271782 3448 271788 3460
rect 270552 3420 271788 3448
rect 270552 3408 270558 3420
rect 271782 3408 271788 3420
rect 271840 3408 271846 3460
rect 285490 3408 285496 3460
rect 285548 3448 285554 3460
rect 291930 3448 291936 3460
rect 285548 3420 291936 3448
rect 285548 3408 285554 3420
rect 291930 3408 291936 3420
rect 291988 3408 291994 3460
rect 292482 3408 292488 3460
rect 292540 3448 292546 3460
rect 307386 3448 307392 3460
rect 292540 3420 307392 3448
rect 292540 3408 292546 3420
rect 307386 3408 307392 3420
rect 307444 3408 307450 3460
rect 308600 3448 308628 3488
rect 315298 3476 315304 3528
rect 315356 3516 315362 3528
rect 343082 3516 343088 3528
rect 315356 3488 343088 3516
rect 315356 3476 315362 3488
rect 343082 3476 343088 3488
rect 343140 3476 343146 3528
rect 349798 3476 349804 3528
rect 349856 3516 349862 3528
rect 414474 3516 414480 3528
rect 349856 3488 414480 3516
rect 349856 3476 349862 3488
rect 414474 3476 414480 3488
rect 414532 3476 414538 3528
rect 439498 3476 439504 3528
rect 439556 3516 439562 3528
rect 582190 3516 582196 3528
rect 439556 3488 582196 3516
rect 439556 3476 439562 3488
rect 582190 3476 582196 3488
rect 582248 3476 582254 3528
rect 313366 3448 313372 3460
rect 308600 3420 313372 3448
rect 313366 3408 313372 3420
rect 313424 3408 313430 3460
rect 339494 3448 339500 3460
rect 316696 3420 339500 3448
rect 27890 3340 27896 3392
rect 27948 3380 27954 3392
rect 28902 3380 28908 3392
rect 27948 3352 28908 3380
rect 27948 3340 27954 3352
rect 28902 3340 28908 3352
rect 28960 3340 28966 3392
rect 59998 3340 60004 3392
rect 60056 3380 60062 3392
rect 60642 3380 60648 3392
rect 60056 3352 60648 3380
rect 60056 3340 60062 3352
rect 60642 3340 60648 3352
rect 60700 3340 60706 3392
rect 71866 3340 71872 3392
rect 71924 3380 71930 3392
rect 72970 3380 72976 3392
rect 71924 3352 72976 3380
rect 71924 3340 71930 3352
rect 72970 3340 72976 3352
rect 73028 3340 73034 3392
rect 73798 3340 73804 3392
rect 73856 3380 73862 3392
rect 74258 3380 74264 3392
rect 73856 3352 74264 3380
rect 73856 3340 73862 3352
rect 74258 3340 74264 3352
rect 74316 3340 74322 3392
rect 86126 3340 86132 3392
rect 86184 3380 86190 3392
rect 86862 3380 86868 3392
rect 86184 3352 86868 3380
rect 86184 3340 86190 3352
rect 86862 3340 86868 3352
rect 86920 3340 86926 3392
rect 93302 3340 93308 3392
rect 93360 3380 93366 3392
rect 174262 3380 174268 3392
rect 93360 3352 174268 3380
rect 93360 3340 93366 3352
rect 174262 3340 174268 3352
rect 174320 3340 174326 3392
rect 183738 3340 183744 3392
rect 183796 3380 183802 3392
rect 202874 3380 202880 3392
rect 183796 3352 202880 3380
rect 183796 3340 183802 3352
rect 202874 3340 202880 3352
rect 202932 3340 202938 3392
rect 206278 3340 206284 3392
rect 206336 3380 206342 3392
rect 232314 3380 232320 3392
rect 206336 3352 232320 3380
rect 206336 3340 206342 3352
rect 232314 3340 232320 3352
rect 232372 3340 232378 3392
rect 250346 3340 250352 3392
rect 250404 3380 250410 3392
rect 251082 3380 251088 3392
rect 250404 3352 251088 3380
rect 250404 3340 250410 3352
rect 251082 3340 251088 3352
rect 251140 3340 251146 3392
rect 282822 3340 282828 3392
rect 282880 3380 282886 3392
rect 287146 3380 287152 3392
rect 282880 3352 287152 3380
rect 282880 3340 282886 3352
rect 287146 3340 287152 3352
rect 287204 3340 287210 3392
rect 289630 3340 289636 3392
rect 289688 3380 289694 3392
rect 300302 3380 300308 3392
rect 289688 3352 300308 3380
rect 289688 3340 289694 3352
rect 300302 3340 300308 3352
rect 300360 3340 300366 3392
rect 300762 3340 300768 3392
rect 300820 3380 300826 3392
rect 309594 3380 309600 3392
rect 300820 3352 309600 3380
rect 300820 3340 300826 3352
rect 309594 3340 309600 3352
rect 309652 3340 309658 3392
rect 100478 3272 100484 3324
rect 100536 3312 100542 3324
rect 184290 3312 184296 3324
rect 100536 3284 184296 3312
rect 100536 3272 100542 3284
rect 184290 3272 184296 3284
rect 184348 3272 184354 3324
rect 193214 3272 193220 3324
rect 193272 3312 193278 3324
rect 194502 3312 194508 3324
rect 193272 3284 194508 3312
rect 193272 3272 193278 3284
rect 194502 3272 194508 3284
rect 194560 3272 194566 3324
rect 194594 3272 194600 3324
rect 194652 3312 194658 3324
rect 202966 3312 202972 3324
rect 194652 3284 202972 3312
rect 194652 3272 194658 3284
rect 202966 3272 202972 3284
rect 203024 3272 203030 3324
rect 207474 3272 207480 3324
rect 207532 3312 207538 3324
rect 225230 3312 225236 3324
rect 207532 3284 225236 3312
rect 207532 3272 207538 3284
rect 225230 3272 225236 3284
rect 225288 3272 225294 3324
rect 225322 3272 225328 3324
rect 225380 3312 225386 3324
rect 226242 3312 226248 3324
rect 225380 3284 226248 3312
rect 225380 3272 225386 3284
rect 226242 3272 226248 3284
rect 226300 3272 226306 3324
rect 282730 3272 282736 3324
rect 282788 3312 282794 3324
rect 282788 3284 286088 3312
rect 282788 3272 282794 3284
rect 103974 3204 103980 3256
rect 104032 3244 104038 3256
rect 186314 3244 186320 3256
rect 104032 3216 186320 3244
rect 104032 3204 104038 3216
rect 186314 3204 186320 3216
rect 186372 3204 186378 3256
rect 200390 3204 200396 3256
rect 200448 3244 200454 3256
rect 224218 3244 224224 3256
rect 200448 3216 224224 3244
rect 200448 3204 200454 3216
rect 224218 3204 224224 3216
rect 224276 3204 224282 3256
rect 261018 3204 261024 3256
rect 261076 3244 261082 3256
rect 262122 3244 262128 3256
rect 261076 3216 262128 3244
rect 261076 3204 261082 3216
rect 262122 3204 262128 3216
rect 262180 3204 262186 3256
rect 113542 3136 113548 3188
rect 113600 3176 113606 3188
rect 114462 3176 114468 3188
rect 113600 3148 114468 3176
rect 113600 3136 113606 3148
rect 114462 3136 114468 3148
rect 114520 3136 114526 3188
rect 115934 3136 115940 3188
rect 115992 3176 115998 3188
rect 117130 3176 117136 3188
rect 115992 3148 117136 3176
rect 115992 3136 115998 3148
rect 117130 3136 117136 3148
rect 117188 3136 117194 3188
rect 167638 3176 167644 3188
rect 117976 3148 167644 3176
rect 107562 3068 107568 3120
rect 107620 3108 107626 3120
rect 117976 3108 118004 3148
rect 167638 3136 167644 3148
rect 167696 3136 167702 3188
rect 180058 3136 180064 3188
rect 180116 3176 180122 3188
rect 186130 3176 186136 3188
rect 180116 3148 186136 3176
rect 180116 3136 180122 3148
rect 186130 3136 186136 3148
rect 186188 3136 186194 3188
rect 192018 3136 192024 3188
rect 192076 3176 192082 3188
rect 213178 3176 213184 3188
rect 192076 3148 213184 3176
rect 192076 3136 192082 3148
rect 213178 3136 213184 3148
rect 213236 3136 213242 3188
rect 220538 3136 220544 3188
rect 220596 3176 220602 3188
rect 220596 3148 234660 3176
rect 220596 3136 220602 3148
rect 169018 3108 169024 3120
rect 107620 3080 118004 3108
rect 118160 3080 169024 3108
rect 107620 3068 107626 3080
rect 79042 3000 79048 3052
rect 79100 3040 79106 3052
rect 79962 3040 79968 3052
rect 79100 3012 79968 3040
rect 79100 3000 79106 3012
rect 79962 3000 79968 3012
rect 80020 3000 80026 3052
rect 114738 3000 114744 3052
rect 114796 3040 114802 3052
rect 118160 3040 118188 3080
rect 169018 3068 169024 3080
rect 169076 3068 169082 3120
rect 190822 3068 190828 3120
rect 190880 3108 190886 3120
rect 204254 3108 204260 3120
rect 190880 3080 204260 3108
rect 190880 3068 190886 3080
rect 204254 3068 204260 3080
rect 204312 3068 204318 3120
rect 214650 3068 214656 3120
rect 214708 3108 214714 3120
rect 233878 3108 233884 3120
rect 214708 3080 233884 3108
rect 214708 3068 214714 3080
rect 233878 3068 233884 3080
rect 233936 3068 233942 3120
rect 234632 3108 234660 3148
rect 241974 3136 241980 3188
rect 242032 3176 242038 3188
rect 242802 3176 242808 3188
rect 242032 3148 242808 3176
rect 242032 3136 242038 3148
rect 242802 3136 242808 3148
rect 242860 3136 242866 3188
rect 281350 3136 281356 3188
rect 281408 3176 281414 3188
rect 285950 3176 285956 3188
rect 281408 3148 285956 3176
rect 281408 3136 281414 3148
rect 285950 3136 285956 3148
rect 286008 3136 286014 3188
rect 286060 3176 286088 3284
rect 288342 3272 288348 3324
rect 288400 3312 288406 3324
rect 297910 3312 297916 3324
rect 288400 3284 297916 3312
rect 288400 3272 288406 3284
rect 297910 3272 297916 3284
rect 297968 3272 297974 3324
rect 309042 3204 309048 3256
rect 309100 3244 309106 3256
rect 316696 3244 316724 3420
rect 339494 3408 339500 3420
rect 339552 3408 339558 3460
rect 352466 3408 352472 3460
rect 352524 3448 352530 3460
rect 421558 3448 421564 3460
rect 352524 3420 421564 3448
rect 352524 3408 352530 3420
rect 421558 3408 421564 3420
rect 421616 3408 421622 3460
rect 431218 3408 431224 3460
rect 431276 3448 431282 3460
rect 575014 3448 575020 3460
rect 431276 3420 575020 3448
rect 431276 3408 431282 3420
rect 575014 3408 575020 3420
rect 575072 3408 575078 3460
rect 334618 3340 334624 3392
rect 334676 3380 334682 3392
rect 375190 3380 375196 3392
rect 334676 3352 375196 3380
rect 334676 3340 334682 3352
rect 375190 3340 375196 3352
rect 375248 3340 375254 3392
rect 375282 3340 375288 3392
rect 375340 3380 375346 3392
rect 467926 3380 467932 3392
rect 375340 3352 467932 3380
rect 375340 3340 375346 3352
rect 467926 3340 467932 3352
rect 467984 3340 467990 3392
rect 493318 3340 493324 3392
rect 493376 3380 493382 3392
rect 564342 3380 564348 3392
rect 493376 3352 564348 3380
rect 493376 3340 493382 3352
rect 564342 3340 564348 3352
rect 564400 3340 564406 3392
rect 331950 3272 331956 3324
rect 332008 3312 332014 3324
rect 360930 3312 360936 3324
rect 332008 3284 360936 3312
rect 332008 3272 332014 3284
rect 360930 3272 360936 3284
rect 360988 3272 360994 3324
rect 369118 3272 369124 3324
rect 369176 3312 369182 3324
rect 453666 3312 453672 3324
rect 369176 3284 453672 3312
rect 369176 3272 369182 3284
rect 453666 3272 453672 3284
rect 453724 3272 453730 3324
rect 489546 3272 489552 3324
rect 489604 3312 489610 3324
rect 557166 3312 557172 3324
rect 489604 3284 557172 3312
rect 489604 3272 489610 3284
rect 557166 3272 557172 3284
rect 557224 3272 557230 3324
rect 309100 3216 316724 3244
rect 309100 3204 309106 3216
rect 319438 3204 319444 3256
rect 319496 3244 319502 3256
rect 346670 3244 346676 3256
rect 319496 3216 346676 3244
rect 319496 3204 319502 3216
rect 346670 3204 346676 3216
rect 346728 3204 346734 3256
rect 377398 3204 377404 3256
rect 377456 3244 377462 3256
rect 460842 3244 460848 3256
rect 377456 3216 460848 3244
rect 377456 3204 377462 3216
rect 460842 3204 460848 3216
rect 460900 3204 460906 3256
rect 482186 3204 482192 3256
rect 482244 3244 482250 3256
rect 546494 3244 546500 3256
rect 482244 3216 546500 3244
rect 482244 3204 482250 3216
rect 546494 3204 546500 3216
rect 546552 3204 546558 3256
rect 288342 3176 288348 3188
rect 286060 3148 288348 3176
rect 288342 3136 288348 3148
rect 288400 3136 288406 3188
rect 322198 3136 322204 3188
rect 322256 3176 322262 3188
rect 350258 3176 350264 3188
rect 322256 3148 350264 3176
rect 322256 3136 322262 3148
rect 350258 3136 350264 3148
rect 350316 3136 350322 3188
rect 380158 3136 380164 3188
rect 380216 3176 380222 3188
rect 446582 3176 446588 3188
rect 380216 3148 446588 3176
rect 380216 3136 380222 3148
rect 446582 3136 446588 3148
rect 446640 3136 446646 3188
rect 451274 3136 451280 3188
rect 451332 3176 451338 3188
rect 452470 3176 452476 3188
rect 451332 3148 452476 3176
rect 451332 3136 451338 3148
rect 452470 3136 452476 3148
rect 452528 3136 452534 3188
rect 486418 3136 486424 3188
rect 486476 3176 486482 3188
rect 550082 3176 550088 3188
rect 486476 3148 550088 3176
rect 486476 3136 486482 3148
rect 550082 3136 550088 3148
rect 550140 3136 550146 3188
rect 242158 3108 242164 3120
rect 234632 3080 242164 3108
rect 242158 3068 242164 3080
rect 242216 3068 242222 3120
rect 258626 3068 258632 3120
rect 258684 3108 258690 3120
rect 259362 3108 259368 3120
rect 258684 3080 259368 3108
rect 258684 3068 258690 3080
rect 259362 3068 259368 3080
rect 259420 3068 259426 3120
rect 331858 3068 331864 3120
rect 331916 3108 331922 3120
rect 353754 3108 353760 3120
rect 331916 3080 353760 3108
rect 331916 3068 331922 3080
rect 353754 3068 353760 3080
rect 353812 3068 353818 3120
rect 374638 3068 374644 3120
rect 374696 3108 374702 3120
rect 432322 3108 432328 3120
rect 374696 3080 432328 3108
rect 374696 3068 374702 3080
rect 432322 3068 432328 3080
rect 432380 3068 432386 3120
rect 481266 3068 481272 3120
rect 481324 3108 481330 3120
rect 539318 3108 539324 3120
rect 481324 3080 539324 3108
rect 481324 3068 481330 3080
rect 539318 3068 539324 3080
rect 539376 3068 539382 3120
rect 114796 3012 118188 3040
rect 114796 3000 114802 3012
rect 124214 3000 124220 3052
rect 124272 3040 124278 3052
rect 125502 3040 125508 3052
rect 124272 3012 125508 3040
rect 124272 3000 124278 3012
rect 125502 3000 125508 3012
rect 125560 3000 125566 3052
rect 148042 3000 148048 3052
rect 148100 3040 148106 3052
rect 191098 3040 191104 3052
rect 148100 3012 191104 3040
rect 148100 3000 148106 3012
rect 191098 3000 191104 3012
rect 191156 3000 191162 3052
rect 194410 3000 194416 3052
rect 194468 3040 194474 3052
rect 204346 3040 204352 3052
rect 194468 3012 204352 3040
rect 194468 3000 194474 3012
rect 204346 3000 204352 3012
rect 204404 3000 204410 3052
rect 217042 3000 217048 3052
rect 217100 3040 217106 3052
rect 217962 3040 217968 3052
rect 217100 3012 217968 3040
rect 217100 3000 217106 3012
rect 217962 3000 217968 3012
rect 218020 3000 218026 3052
rect 224126 3000 224132 3052
rect 224184 3040 224190 3052
rect 243538 3040 243544 3052
rect 224184 3012 243544 3040
rect 224184 3000 224190 3012
rect 243538 3000 243544 3012
rect 243596 3000 243602 3052
rect 269298 3000 269304 3052
rect 269356 3040 269362 3052
rect 271138 3040 271144 3052
rect 269356 3012 271144 3040
rect 269356 3000 269362 3012
rect 271138 3000 271144 3012
rect 271196 3000 271202 3052
rect 337378 3000 337384 3052
rect 337436 3040 337442 3052
rect 382366 3040 382372 3052
rect 337436 3012 382372 3040
rect 337436 3000 337442 3012
rect 382366 3000 382372 3012
rect 382424 3000 382430 3052
rect 410518 3000 410524 3052
rect 410576 3040 410582 3052
rect 439406 3040 439412 3052
rect 410576 3012 439412 3040
rect 410576 3000 410582 3012
rect 439406 3000 439412 3012
rect 439464 3000 439470 3052
rect 478138 3000 478144 3052
rect 478196 3040 478202 3052
rect 532234 3040 532240 3052
rect 478196 3012 532240 3040
rect 478196 3000 478202 3012
rect 532234 3000 532240 3012
rect 532292 3000 532298 3052
rect 159910 2932 159916 2984
rect 159968 2972 159974 2984
rect 193306 2972 193312 2984
rect 159968 2944 193312 2972
rect 159968 2932 159974 2944
rect 193306 2932 193312 2944
rect 193364 2932 193370 2984
rect 221734 2932 221740 2984
rect 221792 2972 221798 2984
rect 221792 2944 225184 2972
rect 221792 2932 221798 2944
rect 168190 2864 168196 2916
rect 168248 2904 168254 2916
rect 188062 2904 188068 2916
rect 168248 2876 188068 2904
rect 168248 2864 168254 2876
rect 188062 2864 188068 2876
rect 188120 2864 188126 2916
rect 201494 2864 201500 2916
rect 201552 2904 201558 2916
rect 208302 2904 208308 2916
rect 201552 2876 208308 2904
rect 201552 2864 201558 2876
rect 208302 2864 208308 2876
rect 208360 2864 208366 2916
rect 187234 2796 187240 2848
rect 187292 2836 187298 2848
rect 194594 2836 194600 2848
rect 187292 2808 194600 2836
rect 187292 2796 187298 2808
rect 194594 2796 194600 2808
rect 194652 2796 194658 2848
rect 205082 2796 205088 2848
rect 205140 2836 205146 2848
rect 209222 2836 209228 2848
rect 205140 2808 209228 2836
rect 205140 2796 205146 2808
rect 209222 2796 209228 2808
rect 209280 2796 209286 2848
rect 225156 2836 225184 2944
rect 225230 2932 225236 2984
rect 225288 2972 225294 2984
rect 232590 2972 232596 2984
rect 225288 2944 232596 2972
rect 225288 2932 225294 2944
rect 232590 2932 232596 2944
rect 232648 2932 232654 2984
rect 475378 2932 475384 2984
rect 475436 2972 475442 2984
rect 525058 2972 525064 2984
rect 475436 2944 525064 2972
rect 475436 2932 475442 2944
rect 525058 2932 525064 2944
rect 525116 2932 525122 2984
rect 473998 2864 474004 2916
rect 474056 2904 474062 2916
rect 517882 2904 517888 2916
rect 474056 2876 517888 2904
rect 474056 2864 474062 2876
rect 517882 2864 517888 2876
rect 517940 2864 517946 2916
rect 235258 2836 235264 2848
rect 225156 2808 235264 2836
rect 235258 2796 235264 2808
rect 235316 2796 235322 2848
rect 336918 2796 336924 2848
rect 336976 2836 336982 2848
rect 336976 2808 337056 2836
rect 336976 2796 336982 2808
rect 337028 2780 337056 2808
rect 339678 2796 339684 2848
rect 339736 2796 339742 2848
rect 343910 2796 343916 2848
rect 343968 2796 343974 2848
rect 502334 2796 502340 2848
rect 502392 2836 502398 2848
rect 503622 2836 503628 2848
rect 502392 2808 503628 2836
rect 502392 2796 502398 2808
rect 503622 2796 503628 2808
rect 503680 2796 503686 2848
rect 337010 2728 337016 2780
rect 337068 2728 337074 2780
rect 339696 2768 339724 2796
rect 340138 2768 340144 2780
rect 339696 2740 340144 2768
rect 340138 2728 340144 2740
rect 340196 2728 340202 2780
rect 343928 2768 343956 2796
rect 344002 2768 344008 2780
rect 343928 2740 344008 2768
rect 344002 2728 344008 2740
rect 344060 2728 344066 2780
rect 400950 756 400956 808
rect 401008 796 401014 808
rect 403710 796 403716 808
rect 401008 768 403716 796
rect 401008 756 401014 768
rect 403710 756 403716 768
rect 403768 756 403774 808
rect 92106 552 92112 604
rect 92164 592 92170 604
rect 92382 592 92388 604
rect 92164 564 92388 592
rect 92164 552 92170 564
rect 92382 552 92388 564
rect 92440 552 92446 604
rect 178954 552 178960 604
rect 179012 592 179018 604
rect 179322 592 179328 604
rect 179012 564 179328 592
rect 179012 552 179018 564
rect 179322 552 179328 564
rect 179380 552 179386 604
rect 238386 552 238392 604
rect 238444 592 238450 604
rect 238662 592 238668 604
rect 238444 564 238668 592
rect 238444 552 238450 564
rect 238662 552 238668 564
rect 238720 552 238726 604
rect 275278 552 275284 604
rect 275336 592 275342 604
rect 275370 592 275376 604
rect 275336 564 275376 592
rect 275336 552 275342 564
rect 275370 552 275376 564
rect 275428 552 275434 604
rect 280338 552 280344 604
rect 280396 592 280402 604
rect 281258 592 281264 604
rect 280396 564 281264 592
rect 280396 552 280402 564
rect 281258 552 281264 564
rect 281316 552 281322 604
rect 304994 552 305000 604
rect 305052 592 305058 604
rect 305178 592 305184 604
rect 305052 564 305184 592
rect 305052 552 305058 564
rect 305178 552 305184 564
rect 305236 552 305242 604
rect 307938 552 307944 604
rect 307996 592 308002 604
rect 308582 592 308588 604
rect 307996 564 308588 592
rect 307996 552 308002 564
rect 308582 552 308588 564
rect 308640 552 308646 604
rect 323118 552 323124 604
rect 323176 592 323182 604
rect 324038 592 324044 604
rect 323176 564 324044 592
rect 323176 552 323182 564
rect 324038 552 324044 564
rect 324096 552 324102 604
rect 325878 552 325884 604
rect 325936 592 325942 604
rect 326430 592 326436 604
rect 325936 564 326436 592
rect 325936 552 325942 564
rect 326430 552 326436 564
rect 326488 552 326494 604
rect 332870 552 332876 604
rect 332928 592 332934 604
rect 333606 592 333612 604
rect 332928 564 333612 592
rect 332928 552 332934 564
rect 333606 552 333612 564
rect 333664 552 333670 604
rect 337010 552 337016 604
rect 337068 592 337074 604
rect 337102 592 337108 604
rect 337068 564 337108 592
rect 337068 552 337074 564
rect 337102 552 337108 564
rect 337160 552 337166 604
rect 340138 552 340144 604
rect 340196 592 340202 604
rect 340690 592 340696 604
rect 340196 564 340696 592
rect 340196 552 340202 564
rect 340690 552 340696 564
rect 340748 552 340754 604
rect 344002 552 344008 604
rect 344060 592 344066 604
rect 344278 592 344284 604
rect 344060 564 344284 592
rect 344060 552 344066 564
rect 344278 552 344284 564
rect 344336 552 344342 604
rect 416958 552 416964 604
rect 417016 592 417022 604
rect 417970 592 417976 604
rect 417016 564 417976 592
rect 417016 552 417022 564
rect 417970 552 417976 564
rect 418028 552 418034 604
rect 425146 552 425152 604
rect 425204 592 425210 604
rect 425330 592 425336 604
rect 425204 564 425336 592
rect 425204 552 425210 564
rect 425330 552 425336 564
rect 425388 552 425394 604
rect 441614 552 441620 604
rect 441672 592 441678 604
rect 441798 592 441804 604
rect 441672 564 441804 592
rect 441672 552 441678 564
rect 441798 552 441804 564
rect 441856 552 441862 604
rect 444374 552 444380 604
rect 444432 592 444438 604
rect 445386 592 445392 604
rect 444432 564 445392 592
rect 444432 552 444438 564
rect 445386 552 445392 564
rect 445444 552 445450 604
rect 448514 552 448520 604
rect 448572 592 448578 604
rect 448974 592 448980 604
rect 448572 564 448980 592
rect 448572 552 448578 564
rect 448974 552 448980 564
rect 449032 552 449038 604
rect 455414 552 455420 604
rect 455472 592 455478 604
rect 456058 592 456064 604
rect 455472 564 456064 592
rect 455472 552 455478 564
rect 456058 552 456064 564
rect 456116 552 456122 604
rect 456794 552 456800 604
rect 456852 592 456858 604
rect 457254 592 457260 604
rect 456852 564 457260 592
rect 456852 552 456858 564
rect 457254 552 457260 564
rect 457312 552 457318 604
rect 499574 552 499580 604
rect 499632 592 499638 604
rect 500126 592 500132 604
rect 499632 564 500132 592
rect 499632 552 499638 564
rect 500126 552 500132 564
rect 500184 552 500190 604
rect 506474 552 506480 604
rect 506532 592 506538 604
rect 507210 592 507216 604
rect 506532 564 507216 592
rect 506532 552 506538 564
rect 507210 552 507216 564
rect 507268 552 507274 604
rect 510614 552 510620 604
rect 510672 592 510678 604
rect 510798 592 510804 604
rect 510672 564 510804 592
rect 510672 552 510678 564
rect 510798 552 510804 564
rect 510856 552 510862 604
rect 513374 552 513380 604
rect 513432 592 513438 604
rect 514386 592 514392 604
rect 513432 564 514392 592
rect 513432 552 513438 564
rect 514386 552 514392 564
rect 514444 552 514450 604
<< via1 >>
rect 133880 700952 133932 701004
rect 218980 700952 219032 701004
rect 235172 700952 235224 701004
rect 434076 700952 434128 701004
rect 133604 700884 133656 700936
rect 348792 700884 348844 700936
rect 364984 700884 365036 700936
rect 433984 700884 434036 700936
rect 133236 700816 133288 700868
rect 397460 700816 397512 700868
rect 132224 700748 132276 700800
rect 154120 700748 154172 700800
rect 170312 700748 170364 700800
rect 434168 700748 434220 700800
rect 131120 700680 131172 700732
rect 413652 700680 413704 700732
rect 105452 700612 105504 700664
rect 434352 700612 434404 700664
rect 438124 700612 438176 700664
rect 494796 700612 494848 700664
rect 133420 700544 133472 700596
rect 462320 700544 462372 700596
rect 133696 700476 133748 700528
rect 478512 700476 478564 700528
rect 40500 700408 40552 700460
rect 434444 700408 434496 700460
rect 442264 700408 442316 700460
rect 559656 700408 559708 700460
rect 132592 700340 132644 700392
rect 527180 700340 527232 700392
rect 132500 700272 132552 700324
rect 543464 700272 543516 700324
rect 133328 700204 133380 700256
rect 332508 700204 332560 700256
rect 132316 700136 132368 700188
rect 283840 700136 283892 700188
rect 300124 700136 300176 700188
rect 436100 700136 436152 700188
rect 132040 700068 132092 700120
rect 267648 700068 267700 700120
rect 133144 700000 133196 700052
rect 202788 700000 202840 700052
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 72424 699660 72476 699712
rect 72976 699660 73028 699712
rect 89168 699660 89220 699712
rect 89628 699660 89680 699712
rect 133052 699660 133104 699712
rect 137836 699660 137888 699712
rect 429844 699660 429896 699712
rect 433892 699660 433944 699712
rect 8024 698232 8076 698284
rect 8208 698232 8260 698284
rect 129648 696940 129700 696992
rect 580172 696940 580224 696992
rect 7932 695444 7984 695496
rect 8208 695444 8260 695496
rect 7932 685856 7984 685908
rect 8116 685856 8168 685908
rect 132132 685856 132184 685908
rect 580172 685856 580224 685908
rect 3792 681708 3844 681760
rect 434536 681708 434588 681760
rect 8116 678988 8168 679040
rect 8024 678920 8076 678972
rect 8024 673480 8076 673532
rect 8208 673480 8260 673532
rect 440884 673480 440936 673532
rect 580172 673480 580224 673532
rect 8024 654100 8076 654152
rect 8208 654100 8260 654152
rect 129556 650020 129608 650072
rect 580172 650020 580224 650072
rect 131948 638936 132000 638988
rect 580172 638936 580224 638988
rect 8024 634788 8076 634840
rect 8208 634788 8260 634840
rect 439504 626560 439556 626612
rect 580172 626560 580224 626612
rect 3056 623772 3108 623824
rect 434260 623772 434312 623824
rect 8024 615476 8076 615528
rect 8208 615476 8260 615528
rect 130936 603100 130988 603152
rect 580172 603100 580224 603152
rect 8024 596164 8076 596216
rect 8208 596164 8260 596216
rect 133972 592016 134024 592068
rect 580172 592016 580224 592068
rect 126244 583652 126296 583704
rect 302792 583652 302844 583704
rect 270408 583584 270460 583636
rect 307024 583584 307076 583636
rect 282828 583516 282880 583568
rect 313464 583516 313516 583568
rect 199384 583448 199436 583500
rect 317696 583448 317748 583500
rect 129004 583380 129056 583432
rect 347504 583380 347556 583432
rect 124864 583312 124916 583364
rect 324136 583312 324188 583364
rect 131028 583244 131080 583296
rect 349528 583244 349580 583296
rect 289728 583176 289780 583228
rect 328368 583176 328420 583228
rect 275928 583108 275980 583160
rect 319720 583108 319772 583160
rect 281172 583040 281224 583092
rect 326160 583040 326212 583092
rect 293868 582972 293920 583024
rect 338856 582972 338908 583024
rect 300400 582904 300452 582956
rect 353760 582904 353812 582956
rect 300492 582836 300544 582888
rect 355968 582836 356020 582888
rect 291108 582768 291160 582820
rect 351736 582768 351788 582820
rect 274548 582700 274600 582752
rect 368664 582700 368716 582752
rect 298928 582632 298980 582684
rect 341064 582632 341116 582684
rect 357992 582632 358044 582684
rect 379060 582632 379112 582684
rect 300308 582564 300360 582616
rect 362408 582564 362460 582616
rect 366640 582564 366692 582616
rect 377588 582564 377640 582616
rect 299296 582496 299348 582548
rect 332600 582496 332652 582548
rect 370872 582496 370924 582548
rect 377312 582496 377364 582548
rect 298744 582428 298796 582480
rect 321928 582428 321980 582480
rect 372896 582428 372948 582480
rect 377496 582428 377548 582480
rect 298836 582360 298888 582412
rect 309232 582360 309284 582412
rect 299204 579640 299256 579692
rect 304816 579640 304868 579692
rect 438216 579640 438268 579692
rect 580172 579640 580224 579692
rect 7656 579572 7708 579624
rect 7932 579572 7984 579624
rect 305092 579572 305144 579624
rect 315212 579572 315264 579624
rect 330760 579572 330812 579624
rect 334808 579572 334860 579624
rect 330668 579504 330720 579556
rect 335176 579504 335228 579556
rect 300216 579436 300268 579488
rect 310980 579436 311032 579488
rect 330576 579436 330628 579488
rect 338672 579436 338724 579488
rect 299480 579300 299532 579352
rect 300676 579300 300728 579352
rect 299572 579164 299624 579216
rect 305092 579300 305144 579352
rect 305184 579300 305236 579352
rect 157340 579028 157392 579080
rect 162400 579028 162452 579080
rect 176660 579028 176712 579080
rect 181720 579028 181772 579080
rect 195980 579028 196032 579080
rect 201040 579028 201092 579080
rect 215300 579028 215352 579080
rect 220360 579028 220412 579080
rect 234620 579028 234672 579080
rect 239680 579028 239732 579080
rect 253940 579028 253992 579080
rect 259000 579028 259052 579080
rect 130384 578960 130436 579012
rect 152556 578960 152608 579012
rect 125692 578892 125744 578944
rect 137836 578892 137888 578944
rect 147588 578892 147640 578944
rect 152280 578892 152332 578944
rect 152372 578892 152424 578944
rect 157248 578892 157300 578944
rect 138664 578756 138716 578808
rect 152464 578756 152516 578808
rect 152556 578756 152608 578808
rect 122748 578688 122800 578740
rect 147588 578688 147640 578740
rect 171876 578960 171928 579012
rect 138112 578620 138164 578672
rect 139584 578620 139636 578672
rect 152280 578620 152332 578672
rect 171600 578892 171652 578944
rect 171692 578892 171744 578944
rect 176568 578892 176620 578944
rect 162308 578756 162360 578808
rect 171784 578756 171836 578808
rect 171876 578756 171928 578808
rect 191196 578960 191248 579012
rect 171600 578620 171652 578672
rect 190920 578892 190972 578944
rect 191012 578892 191064 578944
rect 195888 578892 195940 578944
rect 181628 578756 181680 578808
rect 191104 578756 191156 578808
rect 191196 578756 191248 578808
rect 210516 578960 210568 579012
rect 190920 578620 190972 578672
rect 210240 578892 210292 578944
rect 210332 578892 210384 578944
rect 215208 578892 215260 578944
rect 200948 578756 201000 578808
rect 210424 578756 210476 578808
rect 210516 578756 210568 578808
rect 229836 578960 229888 579012
rect 210240 578620 210292 578672
rect 229560 578892 229612 578944
rect 229652 578892 229704 578944
rect 234528 578892 234580 578944
rect 220268 578756 220320 578808
rect 229744 578756 229796 578808
rect 229836 578756 229888 578808
rect 249156 578960 249208 579012
rect 229560 578620 229612 578672
rect 248880 578892 248932 578944
rect 248972 578892 249024 578944
rect 253848 578892 253900 578944
rect 239588 578756 239640 578808
rect 249064 578756 249116 578808
rect 249156 578756 249208 578808
rect 268476 578960 268528 579012
rect 282920 578960 282972 579012
rect 300216 579028 300268 579080
rect 297180 578960 297232 579012
rect 299572 578960 299624 579012
rect 248880 578620 248932 578672
rect 268108 578892 268160 578944
rect 268292 578892 268344 578944
rect 273168 578892 273220 578944
rect 277952 578892 278004 578944
rect 294604 578892 294656 578944
rect 300216 578892 300268 578944
rect 278044 578824 278096 578876
rect 258908 578756 258960 578808
rect 268384 578756 268436 578808
rect 268476 578756 268528 578808
rect 282920 578756 282972 578808
rect 268108 578620 268160 578672
rect 278044 578620 278096 578672
rect 287704 578824 287756 578876
rect 289820 578824 289872 578876
rect 298008 578824 298060 578876
rect 299388 578756 299440 578808
rect 300216 578756 300268 578808
rect 309784 579300 309836 579352
rect 297088 578688 297140 578740
rect 300124 578688 300176 578740
rect 309968 579300 310020 579352
rect 315856 579300 315908 579352
rect 330024 579300 330076 579352
rect 336556 579368 336608 579420
rect 330576 579300 330628 579352
rect 330668 579300 330720 579352
rect 330760 579300 330812 579352
rect 334440 579300 334492 579352
rect 334716 579300 334768 579352
rect 334808 579300 334860 579352
rect 334900 579300 334952 579352
rect 335176 579300 335228 579352
rect 297180 578620 297232 578672
rect 115204 578552 115256 578604
rect 115940 578552 115992 578604
rect 129096 578552 129148 578604
rect 287704 578552 287756 578604
rect 294512 578552 294564 578604
rect 119344 578484 119396 578536
rect 125692 578484 125744 578536
rect 137928 578484 137980 578536
rect 138020 578484 138072 578536
rect 157248 578484 157300 578536
rect 157340 578484 157392 578536
rect 176568 578484 176620 578536
rect 176660 578484 176712 578536
rect 195888 578484 195940 578536
rect 195980 578484 196032 578536
rect 215208 578484 215260 578536
rect 215300 578484 215352 578536
rect 234528 578484 234580 578536
rect 234620 578484 234672 578536
rect 253848 578484 253900 578536
rect 253940 578484 253992 578536
rect 273168 578484 273220 578536
rect 125508 578348 125560 578400
rect 138664 578416 138716 578468
rect 139584 578416 139636 578468
rect 152372 578416 152424 578468
rect 152464 578416 152516 578468
rect 162308 578416 162360 578468
rect 162400 578416 162452 578468
rect 171692 578416 171744 578468
rect 171784 578416 171836 578468
rect 181628 578416 181680 578468
rect 181720 578416 181772 578468
rect 191012 578416 191064 578468
rect 191104 578416 191156 578468
rect 200948 578416 201000 578468
rect 201040 578416 201092 578468
rect 210332 578416 210384 578468
rect 210424 578416 210476 578468
rect 220268 578416 220320 578468
rect 220360 578416 220412 578468
rect 229652 578416 229704 578468
rect 229744 578416 229796 578468
rect 239588 578416 239640 578468
rect 239680 578416 239732 578468
rect 248972 578416 249024 578468
rect 249064 578416 249116 578468
rect 258908 578416 258960 578468
rect 259000 578416 259052 578468
rect 268292 578416 268344 578468
rect 268384 578416 268436 578468
rect 277952 578416 278004 578468
rect 300124 578484 300176 578536
rect 294512 578416 294564 578468
rect 294604 578416 294656 578468
rect 297088 578416 297140 578468
rect 129280 578348 129332 578400
rect 85396 578280 85448 578332
rect 125600 578280 125652 578332
rect 125784 578280 125836 578332
rect 85580 578212 85632 578264
rect 342996 579368 343048 579420
rect 338672 579300 338724 579352
rect 345112 579300 345164 579352
rect 360384 579300 360436 579352
rect 364248 579300 364300 579352
rect 375380 579300 375432 579352
rect 378968 579300 379020 579352
rect 110328 575492 110380 575544
rect 296720 575492 296772 575544
rect 281264 572704 281316 572756
rect 281264 572568 281316 572620
rect 7656 569916 7708 569968
rect 7840 569916 7892 569968
rect 271788 569916 271840 569968
rect 296720 569916 296772 569968
rect 281080 569780 281132 569832
rect 281264 569780 281316 569832
rect 7840 563048 7892 563100
rect 129464 563048 129516 563100
rect 296720 563048 296772 563100
rect 7932 562912 7984 562964
rect 200120 562096 200172 562148
rect 209688 562096 209740 562148
rect 195796 562028 195848 562080
rect 214748 562028 214800 562080
rect 195704 561960 195756 562012
rect 205548 561960 205600 562012
rect 197268 561892 197320 561944
rect 208676 561892 208728 561944
rect 195888 561824 195940 561876
rect 211620 561824 211672 561876
rect 197176 561756 197228 561808
rect 200120 561756 200172 561808
rect 209688 561688 209740 561740
rect 217876 561688 217928 561740
rect 281080 560260 281132 560312
rect 281264 560260 281316 560312
rect 197084 560192 197136 560244
rect 202052 560192 202104 560244
rect 418804 556248 418856 556300
rect 511264 556248 511316 556300
rect 273168 556180 273220 556232
rect 297824 556180 297876 556232
rect 378784 556180 378836 556232
rect 484400 556180 484452 556232
rect 109408 554752 109460 554804
rect 110328 554752 110380 554804
rect 115940 554752 115992 554804
rect 92112 553936 92164 553988
rect 115296 553936 115348 553988
rect 89168 553868 89220 553920
rect 156604 553868 156656 553920
rect 115112 553800 115164 553852
rect 128452 553800 128504 553852
rect 129004 553800 129056 553852
rect 95056 553732 95108 553784
rect 120724 553732 120776 553784
rect 100760 553664 100812 553716
rect 129188 553664 129240 553716
rect 106464 553596 106516 553648
rect 137284 553596 137336 553648
rect 103704 553528 103756 553580
rect 141424 553528 141476 553580
rect 97816 553460 97868 553512
rect 151084 553460 151136 553512
rect 112352 553392 112404 553444
rect 116032 553392 116084 553444
rect 281264 553392 281316 553444
rect 128452 553324 128504 553376
rect 128636 553324 128688 553376
rect 281356 553324 281408 553376
rect 89628 552644 89680 552696
rect 129004 552644 129056 552696
rect 271512 550604 271564 550656
rect 271788 550604 271840 550656
rect 281264 550604 281316 550656
rect 281356 550604 281408 550656
rect 8024 550536 8076 550588
rect 8116 550536 8168 550588
rect 281080 550468 281132 550520
rect 281264 550468 281316 550520
rect 85488 549856 85540 549908
rect 86408 549856 86460 549908
rect 199384 549856 199436 549908
rect 271512 545776 271564 545828
rect 271788 545776 271840 545828
rect 128636 543804 128688 543856
rect 128544 543668 128596 543720
rect 118608 542376 118660 542428
rect 155224 542376 155276 542428
rect 8116 540948 8168 541000
rect 8208 540948 8260 541000
rect 271512 540948 271564 541000
rect 271604 540948 271656 541000
rect 281080 540948 281132 541000
rect 281264 540948 281316 541000
rect 3976 538432 4028 538484
rect 4804 538432 4856 538484
rect 286968 538228 287020 538280
rect 297640 538228 297692 538280
rect 117780 536800 117832 536852
rect 140044 536800 140096 536852
rect 128452 534080 128504 534132
rect 281264 534080 281316 534132
rect 128544 534012 128596 534064
rect 281356 534012 281408 534064
rect 117780 532720 117832 532772
rect 153844 532720 153896 532772
rect 294604 532720 294656 532772
rect 297364 532720 297416 532772
rect 128452 531292 128504 531344
rect 128544 531292 128596 531344
rect 271788 531292 271840 531344
rect 271972 531292 272024 531344
rect 281264 531292 281316 531344
rect 281356 531292 281408 531344
rect 117964 529864 118016 529916
rect 119344 529864 119396 529916
rect 118608 525036 118660 525088
rect 128360 525036 128412 525088
rect 129280 525036 129332 525088
rect 271788 524492 271840 524544
rect 281264 524492 281316 524544
rect 70216 524424 70268 524476
rect 82820 524424 82872 524476
rect 128452 524424 128504 524476
rect 271788 524356 271840 524408
rect 281264 524356 281316 524408
rect 128636 524288 128688 524340
rect 8208 521636 8260 521688
rect 8392 521636 8444 521688
rect 280068 521636 280120 521688
rect 297548 521636 297600 521688
rect 128452 521568 128504 521620
rect 129096 521568 129148 521620
rect 293960 521568 294012 521620
rect 294604 521568 294656 521620
rect 85304 521228 85356 521280
rect 293960 521228 294012 521280
rect 199752 521092 199804 521144
rect 222384 521092 222436 521144
rect 199844 521024 199896 521076
rect 222568 521024 222620 521076
rect 196440 520956 196492 521008
rect 222476 520956 222528 521008
rect 117320 520888 117372 520940
rect 128452 520888 128504 520940
rect 195060 520888 195112 520940
rect 222660 520888 222712 520940
rect 128360 518916 128412 518968
rect 128636 518916 128688 518968
rect 278688 518916 278740 518968
rect 297456 518916 297508 518968
rect 89352 518848 89404 518900
rect 122564 518848 122616 518900
rect 122840 518848 122892 518900
rect 129740 518848 129792 518900
rect 109592 518780 109644 518832
rect 113824 518780 113876 518832
rect 115204 518780 115256 518832
rect 86592 518644 86644 518696
rect 99288 518712 99340 518764
rect 99380 518712 99432 518764
rect 122472 518712 122524 518764
rect 127716 518780 127768 518832
rect 109040 518644 109092 518696
rect 109132 518644 109184 518696
rect 129740 518508 129792 518560
rect 130384 518508 130436 518560
rect 98000 518372 98052 518424
rect 127624 518372 127676 518424
rect 106648 518304 106700 518356
rect 144184 518304 144236 518356
rect 100944 518236 100996 518288
rect 152464 518236 152516 518288
rect 196348 518236 196400 518288
rect 218980 518236 219032 518288
rect 92296 518168 92348 518220
rect 127072 518168 127124 518220
rect 297364 518168 297416 518220
rect 205640 517488 205692 517540
rect 206652 517488 206704 517540
rect 505744 517488 505796 517540
rect 506848 517488 506900 517540
rect 282736 516128 282788 516180
rect 297456 516128 297508 516180
rect 271788 514768 271840 514820
rect 281264 514768 281316 514820
rect 271696 514700 271748 514752
rect 281356 514700 281408 514752
rect 271696 511980 271748 512032
rect 271788 511980 271840 512032
rect 281264 511980 281316 512032
rect 281356 511980 281408 512032
rect 281080 511844 281132 511896
rect 281264 511844 281316 511896
rect 293776 509260 293828 509312
rect 296720 509260 296772 509312
rect 128360 509192 128412 509244
rect 128636 509192 128688 509244
rect 271512 507152 271564 507204
rect 271788 507152 271840 507204
rect 380348 506608 380400 506660
rect 380624 506608 380676 506660
rect 191104 506472 191156 506524
rect 296720 506472 296772 506524
rect 297180 505044 297232 505096
rect 298008 505044 298060 505096
rect 8208 502324 8260 502376
rect 8392 502324 8444 502376
rect 271512 502324 271564 502376
rect 271604 502324 271656 502376
rect 281080 502324 281132 502376
rect 281264 502324 281316 502376
rect 96528 500896 96580 500948
rect 380348 500896 380400 500948
rect 103520 500828 103572 500880
rect 104808 500828 104860 500880
rect 377680 500828 377732 500880
rect 129372 500420 129424 500472
rect 377404 500420 377456 500472
rect 130844 500352 130896 500404
rect 380624 500352 380676 500404
rect 130660 500284 130712 500336
rect 580448 500284 580500 500336
rect 70308 500216 70360 500268
rect 95240 500216 95292 500268
rect 96528 500216 96580 500268
rect 130752 500216 130804 500268
rect 580540 500216 580592 500268
rect 128360 499536 128412 499588
rect 128636 499536 128688 499588
rect 298836 499400 298888 499452
rect 302424 499400 302476 499452
rect 324228 499060 324280 499112
rect 379060 499060 379112 499112
rect 298928 498992 298980 499044
rect 310520 498992 310572 499044
rect 321468 498992 321520 499044
rect 378968 498992 379020 499044
rect 300308 498924 300360 498976
rect 311900 498924 311952 498976
rect 317328 498924 317380 498976
rect 377588 498924 377640 498976
rect 309048 498856 309100 498908
rect 377496 498856 377548 498908
rect 118056 498788 118108 498840
rect 302056 498788 302108 498840
rect 375288 498788 375340 498840
rect 478880 498788 478932 498840
rect 131856 498176 131908 498228
rect 579896 498176 579948 498228
rect 116032 498040 116084 498092
rect 347320 498040 347372 498092
rect 120724 497972 120776 498024
rect 121368 497972 121420 498024
rect 338856 497972 338908 498024
rect 128268 497904 128320 497956
rect 334440 497904 334492 497956
rect 336004 497904 336056 497956
rect 349344 497904 349396 497956
rect 111708 497836 111760 497888
rect 115296 497836 115348 497888
rect 313280 497836 313332 497888
rect 318708 497836 318760 497888
rect 355784 497836 355836 497888
rect 155224 497768 155276 497820
rect 319720 497768 319772 497820
rect 320088 497768 320140 497820
rect 357992 497768 358044 497820
rect 284208 497700 284260 497752
rect 368480 497700 368532 497752
rect 291016 497632 291068 497684
rect 377128 497632 377180 497684
rect 108948 497564 109000 497616
rect 116032 497564 116084 497616
rect 127624 497564 127676 497616
rect 128268 497564 128320 497616
rect 281080 497564 281132 497616
rect 281264 497564 281316 497616
rect 284116 497564 284168 497616
rect 374920 497564 374972 497616
rect 83832 497496 83884 497548
rect 127164 497496 127216 497548
rect 360016 497496 360068 497548
rect 111800 497428 111852 497480
rect 125968 497428 126020 497480
rect 372712 497428 372764 497480
rect 289636 497360 289688 497412
rect 366456 497360 366508 497412
rect 285588 497292 285640 497344
rect 345112 497292 345164 497344
rect 292396 497224 292448 497276
rect 351552 497224 351604 497276
rect 275836 497156 275888 497208
rect 306840 497156 306892 497208
rect 307024 497156 307076 497208
rect 362224 497156 362276 497208
rect 277308 497088 277360 497140
rect 317512 497088 317564 497140
rect 334624 497088 334676 497140
rect 343088 497088 343140 497140
rect 288256 497020 288308 497072
rect 321744 497020 321796 497072
rect 307576 496952 307628 497004
rect 315028 496952 315080 497004
rect 315304 496952 315356 497004
rect 323952 496952 324004 497004
rect 155224 496884 155276 496936
rect 155868 496884 155920 496936
rect 304816 496884 304868 496936
rect 309324 496884 309376 496936
rect 324964 496884 325016 496936
rect 328184 496884 328236 496936
rect 331864 496884 331916 496936
rect 336648 496884 336700 496936
rect 129188 496816 129240 496868
rect 364248 496816 364300 496868
rect 297180 495456 297232 495508
rect 298008 495456 298060 495508
rect 308864 492736 308916 492788
rect 309048 492736 309100 492788
rect 302056 492600 302108 492652
rect 302148 492600 302200 492652
rect 301964 491240 302016 491292
rect 302148 491240 302200 491292
rect 299572 490560 299624 490612
rect 300584 490560 300636 490612
rect 128360 489812 128412 489864
rect 128636 489812 128688 489864
rect 271512 487772 271564 487824
rect 271788 487772 271840 487824
rect 281264 485868 281316 485920
rect 8116 485800 8168 485852
rect 438308 485800 438360 485852
rect 580172 485800 580224 485852
rect 8208 485732 8260 485784
rect 281264 485732 281316 485784
rect 271512 483080 271564 483132
rect 271696 483080 271748 483132
rect 7932 482944 7984 482996
rect 8208 482944 8260 482996
rect 271696 482944 271748 482996
rect 271788 482944 271840 482996
rect 301872 481652 301924 481704
rect 301964 481652 302016 481704
rect 308772 481584 308824 481636
rect 308864 481584 308916 481636
rect 3148 481040 3200 481092
rect 4896 481040 4948 481092
rect 128360 480292 128412 480344
rect 128636 480292 128688 480344
rect 271788 476076 271840 476128
rect 281264 476076 281316 476128
rect 281356 476076 281408 476128
rect 271696 476008 271748 476060
rect 281264 473356 281316 473408
rect 281356 473356 281408 473408
rect 308864 473356 308916 473408
rect 308772 473288 308824 473340
rect 302056 469072 302108 469124
rect 302056 468936 302108 468988
rect 271512 468460 271564 468512
rect 271788 468460 271840 468512
rect 281264 466488 281316 466540
rect 8116 466420 8168 466472
rect 8208 466352 8260 466404
rect 281264 466352 281316 466404
rect 271512 463768 271564 463820
rect 271696 463768 271748 463820
rect 271696 463632 271748 463684
rect 271788 463632 271840 463684
rect 306840 463632 306892 463684
rect 307024 463632 307076 463684
rect 130568 462340 130620 462392
rect 580172 462340 580224 462392
rect 281080 458804 281132 458856
rect 281264 458804 281316 458856
rect 271788 456764 271840 456816
rect 271696 456696 271748 456748
rect 7840 453976 7892 454028
rect 8024 453976 8076 454028
rect 3240 451324 3292 451376
rect 261300 451324 261352 451376
rect 134064 451256 134116 451308
rect 579896 451256 579948 451308
rect 271512 449148 271564 449200
rect 271788 449148 271840 449200
rect 302056 448536 302108 448588
rect 302240 448536 302292 448588
rect 281264 447176 281316 447228
rect 261300 447040 261352 447092
rect 265992 447040 266044 447092
rect 281264 447040 281316 447092
rect 271512 444456 271564 444508
rect 271696 444456 271748 444508
rect 7840 444388 7892 444440
rect 7932 444388 7984 444440
rect 265992 444320 266044 444372
rect 266084 444320 266136 444372
rect 271696 444320 271748 444372
rect 271788 444320 271840 444372
rect 306840 444320 306892 444372
rect 307024 444320 307076 444372
rect 308772 442960 308824 443012
rect 308864 442960 308916 443012
rect 281080 439492 281132 439544
rect 281264 439492 281316 439544
rect 301872 438812 301924 438864
rect 302056 438812 302108 438864
rect 266084 437452 266136 437504
rect 271788 437452 271840 437504
rect 265992 437384 266044 437436
rect 271696 437384 271748 437436
rect 306840 434732 306892 434784
rect 307024 434732 307076 434784
rect 128360 431876 128412 431928
rect 128636 431876 128688 431928
rect 265808 429836 265860 429888
rect 266084 429836 266136 429888
rect 271512 429836 271564 429888
rect 271788 429836 271840 429888
rect 301872 429156 301924 429208
rect 302056 429156 302108 429208
rect 281264 427864 281316 427916
rect 8116 427796 8168 427848
rect 302148 427796 302200 427848
rect 8208 427728 8260 427780
rect 281264 427728 281316 427780
rect 302056 427728 302108 427780
rect 265808 425144 265860 425196
rect 265992 425144 266044 425196
rect 271512 425144 271564 425196
rect 271696 425144 271748 425196
rect 7932 425008 7984 425060
rect 8208 425008 8260 425060
rect 265992 425008 266044 425060
rect 266176 425008 266228 425060
rect 271696 425008 271748 425060
rect 271788 425008 271840 425060
rect 308772 423648 308824 423700
rect 308864 423648 308916 423700
rect 281264 423580 281316 423632
rect 281540 423580 281592 423632
rect 128360 422356 128412 422408
rect 128636 422356 128688 422408
rect 302056 418140 302108 418192
rect 302056 418004 302108 418056
rect 7932 415420 7984 415472
rect 8116 415420 8168 415472
rect 132960 415420 133012 415472
rect 579804 415420 579856 415472
rect 281632 413924 281684 413976
rect 281816 413924 281868 413976
rect 265716 411136 265768 411188
rect 265900 411136 265952 411188
rect 254584 411068 254636 411120
rect 269580 411068 269632 411120
rect 254676 411000 254728 411052
rect 266360 411000 266412 411052
rect 258724 410932 258776 410984
rect 267004 410932 267056 410984
rect 226156 410864 226208 410916
rect 270776 410864 270828 410916
rect 223396 410796 223448 410848
rect 266544 410796 266596 410848
rect 246028 410728 246080 410780
rect 270684 410728 270736 410780
rect 211988 410660 212040 410712
rect 258724 410660 258776 410712
rect 258816 410660 258868 410712
rect 266728 410660 266780 410712
rect 206284 410592 206336 410644
rect 270500 410592 270552 410644
rect 203340 410524 203392 410576
rect 254584 410524 254636 410576
rect 257252 410524 257304 410576
rect 269212 410524 269264 410576
rect 240324 410456 240376 410508
rect 266452 410456 266504 410508
rect 237564 410388 237616 410440
rect 258816 410388 258868 410440
rect 260380 410388 260432 410440
rect 267280 410388 267332 410440
rect 234620 410320 234672 410372
rect 257252 410320 257304 410372
rect 257344 410320 257396 410372
rect 269304 410320 269356 410372
rect 231860 410252 231912 410304
rect 270868 410252 270920 410304
rect 228916 410184 228968 410236
rect 270592 410184 270644 410236
rect 200028 410116 200080 410168
rect 217692 410116 217744 410168
rect 251732 410116 251784 410168
rect 257344 410116 257396 410168
rect 257436 410116 257488 410168
rect 269396 410116 269448 410168
rect 195520 410048 195572 410100
rect 220452 410048 220504 410100
rect 195612 409980 195664 410032
rect 214748 409980 214800 410032
rect 248972 409980 249024 410032
rect 269488 410048 269540 410100
rect 199936 409912 199988 409964
rect 209044 409912 209096 409964
rect 243268 409912 243320 409964
rect 266636 409980 266688 410032
rect 263140 409912 263192 409964
rect 267372 409912 267424 409964
rect 196992 409844 197044 409896
rect 200580 409844 200632 409896
rect 265900 409844 265952 409896
rect 268752 409844 268804 409896
rect 196808 409640 196860 409692
rect 202880 409640 202932 409692
rect 196900 409572 196952 409624
rect 205640 409572 205692 409624
rect 195428 409504 195480 409556
rect 209780 409504 209832 409556
rect 195152 409436 195204 409488
rect 212540 409436 212592 409488
rect 196624 409368 196676 409420
rect 215300 409368 215352 409420
rect 196716 409300 196768 409352
rect 219440 409300 219492 409352
rect 195336 409232 195388 409284
rect 219532 409232 219584 409284
rect 196532 409164 196584 409216
rect 222200 409164 222252 409216
rect 195244 409096 195296 409148
rect 222292 409096 222344 409148
rect 8116 408484 8168 408536
rect 271604 408484 271656 408536
rect 271972 408484 272024 408536
rect 8208 408348 8260 408400
rect 265716 408348 265768 408400
rect 266084 408348 266136 408400
rect 188344 407804 188396 407856
rect 380532 407804 380584 407856
rect 70124 407736 70176 407788
rect 104808 407736 104860 407788
rect 416780 407736 416832 407788
rect 155224 407600 155276 407652
rect 155868 407600 155920 407652
rect 155868 407192 155920 407244
rect 416872 407192 416924 407244
rect 127808 407124 127860 407176
rect 411260 407124 411312 407176
rect 197728 406512 197780 406564
rect 293960 406512 294012 406564
rect 199384 406444 199436 406496
rect 402980 406444 403032 406496
rect 293960 406376 294012 406428
rect 294604 406376 294656 406428
rect 308772 404336 308824 404388
rect 308864 404336 308916 404388
rect 301780 401616 301832 401668
rect 302056 401616 302108 401668
rect 8208 400868 8260 400920
rect 8392 400868 8444 400920
rect 120908 398896 120960 398948
rect 121368 398896 121420 398948
rect 125692 398896 125744 398948
rect 71688 398828 71740 398880
rect 85488 398828 85540 398880
rect 110972 398828 111024 398880
rect 111708 398828 111760 398880
rect 126060 398828 126112 398880
rect 113548 398760 113600 398812
rect 113824 398760 113876 398812
rect 126980 398760 127032 398812
rect 127808 398760 127860 398812
rect 271604 398760 271656 398812
rect 271788 398760 271840 398812
rect 85488 398692 85540 398744
rect 90272 398692 90324 398744
rect 125600 398216 125652 398268
rect 128268 398216 128320 398268
rect 138020 398216 138072 398268
rect 100668 398148 100720 398200
rect 113548 398148 113600 398200
rect 75828 398080 75880 398132
rect 115940 398080 115992 398132
rect 127256 398080 127308 398132
rect 128268 398080 128320 398132
rect 155224 398080 155276 398132
rect 80796 397740 80848 397792
rect 124128 397740 124180 397792
rect 106004 397672 106056 397724
rect 130108 397672 130160 397724
rect 95884 397604 95936 397656
rect 126244 397604 126296 397656
rect 85948 397536 86000 397588
rect 128268 397536 128320 397588
rect 115848 397468 115900 397520
rect 127624 397468 127676 397520
rect 124128 397400 124180 397452
rect 124864 397400 124916 397452
rect 125784 397400 125836 397452
rect 71504 396720 71556 396772
rect 117964 396720 118016 396772
rect 126336 396720 126388 396772
rect 8024 396040 8076 396092
rect 8392 396040 8444 396092
rect 83924 395972 83976 396024
rect 84568 395972 84620 396024
rect 71596 395700 71648 395752
rect 96620 395836 96672 395888
rect 83740 395632 83792 395684
rect 72332 395496 72384 395548
rect 84108 395700 84160 395752
rect 84568 395700 84620 395752
rect 84016 395632 84068 395684
rect 99288 395700 99340 395752
rect 108948 395700 109000 395752
rect 125876 395700 125928 395752
rect 126888 395632 126940 395684
rect 168656 395564 168708 395616
rect 179512 395496 179564 395548
rect 8024 394680 8076 394732
rect 8116 394680 8168 394732
rect 308588 394544 308640 394596
rect 308864 394544 308916 394596
rect 128360 393252 128412 393304
rect 128636 393252 128688 393304
rect 402980 393252 403032 393304
rect 403900 393252 403952 393304
rect 266176 392572 266228 392624
rect 436192 392572 436244 392624
rect 301872 391960 301924 392012
rect 302056 391960 302108 392012
rect 126888 391892 126940 391944
rect 199384 391892 199436 391944
rect 458824 389376 458876 389428
rect 475844 389376 475896 389428
rect 416688 389308 416740 389360
rect 464252 389308 464304 389360
rect 418068 389240 418120 389292
rect 487436 389240 487488 389292
rect 8116 389172 8168 389224
rect 416596 389172 416648 389224
rect 499028 389172 499080 389224
rect 271512 389104 271564 389156
rect 271604 389104 271656 389156
rect 297180 389104 297232 389156
rect 298008 389104 298060 389156
rect 8208 389036 8260 389088
rect 126888 386316 126940 386368
rect 130384 386316 130436 386368
rect 281356 386316 281408 386368
rect 281540 386316 281592 386368
rect 306840 386316 306892 386368
rect 307024 386316 307076 386368
rect 344928 385704 344980 385756
rect 408868 385704 408920 385756
rect 294604 385636 294656 385688
rect 388260 385636 388312 385688
rect 365628 385568 365680 385620
rect 392860 385568 392912 385620
rect 349068 385500 349120 385552
rect 385868 385500 385920 385552
rect 355876 385432 355928 385484
rect 399668 385432 399720 385484
rect 353208 385364 353260 385416
rect 402060 385364 402112 385416
rect 357348 385296 357400 385348
rect 406660 385296 406712 385348
rect 347688 385228 347740 385280
rect 397460 385228 397512 385280
rect 343548 385160 343600 385212
rect 395068 385160 395120 385212
rect 355968 385092 356020 385144
rect 413468 385092 413520 385144
rect 367008 385024 367060 385076
rect 390468 385024 390520 385076
rect 126336 384956 126388 385008
rect 130292 384956 130344 385008
rect 271512 384208 271564 384260
rect 271696 384208 271748 384260
rect 128360 383664 128412 383716
rect 128636 383664 128688 383716
rect 301504 381488 301556 381540
rect 301964 381488 302016 381540
rect 380900 381488 380952 381540
rect 8208 379516 8260 379568
rect 297180 379516 297232 379568
rect 298008 379516 298060 379568
rect 8024 379448 8076 379500
rect 271696 379448 271748 379500
rect 271788 379448 271840 379500
rect 281172 376796 281224 376848
rect 281540 376796 281592 376848
rect 306840 376728 306892 376780
rect 307024 376728 307076 376780
rect 308588 376728 308640 376780
rect 308680 376728 308732 376780
rect 351828 376728 351880 376780
rect 380900 376728 380952 376780
rect 281080 376660 281132 376712
rect 281172 376660 281224 376712
rect 7840 375300 7892 375352
rect 8024 375300 8076 375352
rect 129096 374076 129148 374128
rect 128820 374008 128872 374060
rect 364248 374008 364300 374060
rect 380900 374008 380952 374060
rect 414664 374008 414716 374060
rect 456800 374008 456852 374060
rect 128360 373940 128412 373992
rect 128544 373940 128596 373992
rect 347596 369860 347648 369912
rect 380900 369860 380952 369912
rect 128544 369792 128596 369844
rect 128636 369724 128688 369776
rect 281080 367140 281132 367192
rect 281356 367140 281408 367192
rect 281080 367004 281132 367056
rect 281356 367004 281408 367056
rect 306840 367004 306892 367056
rect 307024 367004 307076 367056
rect 2964 366120 3016 366172
rect 4988 366120 5040 366172
rect 308680 365780 308732 365832
rect 308864 365780 308916 365832
rect 7840 365712 7892 365764
rect 8116 365712 8168 365764
rect 128912 365644 128964 365696
rect 197728 365644 197780 365696
rect 308680 365644 308732 365696
rect 308864 365644 308916 365696
rect 333888 362924 333940 362976
rect 380900 362924 380952 362976
rect 8116 360204 8168 360256
rect 128820 360204 128872 360256
rect 129096 360204 129148 360256
rect 271696 360204 271748 360256
rect 271788 360204 271840 360256
rect 8208 360136 8260 360188
rect 281080 357484 281132 357536
rect 281172 357484 281224 357536
rect 306840 357416 306892 357468
rect 307024 357416 307076 357468
rect 308680 357416 308732 357468
rect 281080 357348 281132 357400
rect 281172 357348 281224 357400
rect 308864 357348 308916 357400
rect 185584 355988 185636 356040
rect 188344 355988 188396 356040
rect 8208 354628 8260 354680
rect 8392 354628 8444 354680
rect 354588 353268 354640 353320
rect 380900 353268 380952 353320
rect 129740 350548 129792 350600
rect 130476 350548 130528 350600
rect 128728 347896 128780 347948
rect 281080 347828 281132 347880
rect 281356 347828 281408 347880
rect 128636 347760 128688 347812
rect 128728 347760 128780 347812
rect 129096 347760 129148 347812
rect 281080 347692 281132 347744
rect 281356 347692 281408 347744
rect 306840 347692 306892 347744
rect 306932 347692 306984 347744
rect 365536 347692 365588 347744
rect 386788 347692 386840 347744
rect 360108 347624 360160 347676
rect 391388 347624 391440 347676
rect 358728 347556 358780 347608
rect 393596 347556 393648 347608
rect 362868 347488 362920 347540
rect 398196 347488 398248 347540
rect 362776 347420 362828 347472
rect 402796 347420 402848 347472
rect 350540 347352 350592 347404
rect 395988 347352 396040 347404
rect 342168 347284 342220 347336
rect 388996 347284 389048 347336
rect 361488 347216 361540 347268
rect 407396 347216 407448 347268
rect 354496 347148 354548 347200
rect 400588 347148 400640 347200
rect 361396 347080 361448 347132
rect 414388 347080 414440 347132
rect 274456 347012 274508 347064
rect 310612 347012 310664 347064
rect 333796 347012 333848 347064
rect 411996 347012 412048 347064
rect 130292 346468 130344 346520
rect 132776 346468 132828 346520
rect 308680 346400 308732 346452
rect 308772 346400 308824 346452
rect 128728 345516 128780 345568
rect 129096 345516 129148 345568
rect 8208 345040 8260 345092
rect 8392 345040 8444 345092
rect 504824 345040 504876 345092
rect 579988 345040 580040 345092
rect 135260 342864 135312 342916
rect 191104 342864 191156 342916
rect 199660 342728 199712 342780
rect 200212 342728 200264 342780
rect 128820 342456 128872 342508
rect 135260 342456 135312 342508
rect 503812 341980 503864 342032
rect 504180 341980 504232 342032
rect 126060 340824 126112 340876
rect 408500 340824 408552 340876
rect 127256 340756 127308 340808
rect 404360 340756 404412 340808
rect 503904 340756 503956 340808
rect 504732 340824 504784 340876
rect 127716 340688 127768 340740
rect 381636 340688 381688 340740
rect 130476 340620 130528 340672
rect 381544 340620 381596 340672
rect 132776 340552 132828 340604
rect 383660 340552 383712 340604
rect 130200 340416 130252 340468
rect 138020 340416 138072 340468
rect 154580 340416 154632 340468
rect 173900 340484 173952 340536
rect 157340 340348 157392 340400
rect 183468 340416 183520 340468
rect 202788 340416 202840 340468
rect 240140 340484 240192 340536
rect 215208 340416 215260 340468
rect 240048 340416 240100 340468
rect 249708 340416 249760 340468
rect 269028 340484 269080 340536
rect 259460 340416 259512 340468
rect 269120 340416 269172 340468
rect 273260 340416 273312 340468
rect 280160 340484 280212 340536
rect 333244 340416 333296 340468
rect 193220 340348 193272 340400
rect 224960 340348 225012 340400
rect 230480 340348 230532 340400
rect 173992 340280 174044 340332
rect 183468 340280 183520 340332
rect 215392 340280 215444 340332
rect 224868 340280 224920 340332
rect 280160 340280 280212 340332
rect 292488 340348 292540 340400
rect 292672 340280 292724 340332
rect 318892 340348 318944 340400
rect 331128 340348 331180 340400
rect 318800 340280 318852 340332
rect 357440 340348 357492 340400
rect 362224 340348 362276 340400
rect 381728 340348 381780 340400
rect 114468 340212 114520 340264
rect 126060 340212 126112 340264
rect 331128 340212 331180 340264
rect 333244 340212 333296 340264
rect 357440 340212 357492 340264
rect 362224 340212 362276 340264
rect 110328 340144 110380 340196
rect 127256 340144 127308 340196
rect 196348 338988 196400 339040
rect 209780 338988 209832 339040
rect 199752 338920 199804 338972
rect 213920 338920 213972 338972
rect 199844 338852 199896 338904
rect 215300 338852 215352 338904
rect 196440 338784 196492 338836
rect 222200 338784 222252 338836
rect 257988 338784 258040 338836
rect 267280 338784 267332 338836
rect 195060 338716 195112 338768
rect 220820 338716 220872 338768
rect 237288 338716 237340 338768
rect 267372 338716 267424 338768
rect 262128 338580 262180 338632
rect 268752 338580 268804 338632
rect 281080 338104 281132 338156
rect 281264 338104 281316 338156
rect 306840 338104 306892 338156
rect 307024 338104 307076 338156
rect 308772 338104 308824 338156
rect 350264 338104 350316 338156
rect 350540 338104 350592 338156
rect 107568 338036 107620 338088
rect 97908 337968 97960 338020
rect 127072 337968 127124 338020
rect 231860 337968 231912 338020
rect 244832 337968 244884 338020
rect 250996 337968 251048 338020
rect 260196 337968 260248 338020
rect 301504 338036 301556 338088
rect 308864 337968 308916 338020
rect 112812 337900 112864 337952
rect 113088 337900 113140 337952
rect 127164 337900 127216 337952
rect 226156 337900 226208 337952
rect 248512 337900 248564 337952
rect 253756 337900 253808 337952
rect 263140 337900 263192 337952
rect 122656 337832 122708 337884
rect 127716 337832 127768 337884
rect 220452 337832 220504 337884
rect 239404 337832 239456 337884
rect 211804 337764 211856 337816
rect 240784 337764 240836 337816
rect 242164 337764 242216 337816
rect 246028 337764 246080 337816
rect 249064 337764 249116 337816
rect 257436 337764 257488 337816
rect 92756 337696 92808 337748
rect 93768 337696 93820 337748
rect 102876 337696 102928 337748
rect 103428 337696 103480 337748
rect 203340 337696 203392 337748
rect 207664 337696 207716 337748
rect 214748 337696 214800 337748
rect 258724 337696 258776 337748
rect 206100 337628 206152 337680
rect 255596 337628 255648 337680
rect 117964 337560 118016 337612
rect 128176 337560 128228 337612
rect 297272 337560 297324 337612
rect 401508 337560 401560 337612
rect 460572 337560 460624 337612
rect 72884 337492 72936 337544
rect 130292 337492 130344 337544
rect 299572 337492 299624 337544
rect 411168 337492 411220 337544
rect 472164 337492 472216 337544
rect 77852 337424 77904 337476
rect 99288 337424 99340 337476
rect 329840 337424 329892 337476
rect 408408 337424 408460 337476
rect 483756 337424 483808 337476
rect 87788 337356 87840 337408
rect 117228 337356 117280 337408
rect 380440 337356 380492 337408
rect 413928 337356 413980 337408
rect 495348 337356 495400 337408
rect 223212 337288 223264 337340
rect 237656 337288 237708 337340
rect 239404 337288 239456 337340
rect 246304 337288 246356 337340
rect 228916 337220 228968 337272
rect 236000 337220 236052 337272
rect 242808 337220 242860 337272
rect 249064 337220 249116 337272
rect 251732 337220 251784 337272
rect 260104 337220 260156 337272
rect 271788 336880 271840 336932
rect 200580 336812 200632 336864
rect 201408 336812 201460 336864
rect 234620 336812 234672 336864
rect 237472 336812 237524 336864
rect 237564 336812 237616 336864
rect 239404 336812 239456 336864
rect 240048 336812 240100 336864
rect 243084 336812 243136 336864
rect 247684 336812 247736 336864
rect 248788 336812 248840 336864
rect 254492 336812 254544 336864
rect 258448 336812 258500 336864
rect 265900 336812 265952 336864
rect 269672 336812 269724 336864
rect 271696 336812 271748 336864
rect 2964 336744 3016 336796
rect 434720 336744 434772 336796
rect 82728 336676 82780 336728
rect 125968 336676 126020 336728
rect 258172 336676 258224 336728
rect 258448 336676 258500 336728
rect 128728 335996 128780 336048
rect 129096 335996 129148 336048
rect 503628 331168 503680 331220
rect 503996 331168 504048 331220
rect 271420 330488 271472 330540
rect 271604 330488 271656 330540
rect 244832 328448 244884 328500
rect 248696 328448 248748 328500
rect 281172 328448 281224 328500
rect 281264 328448 281316 328500
rect 307024 328380 307076 328432
rect 503536 328380 503588 328432
rect 503720 328380 503772 328432
rect 307024 328244 307076 328296
rect 308772 327156 308824 327208
rect 258172 327088 258224 327140
rect 258356 327088 258408 327140
rect 308864 327088 308916 327140
rect 128728 327020 128780 327072
rect 129096 327020 129148 327072
rect 8024 325660 8076 325712
rect 8208 325660 8260 325712
rect 128360 325660 128412 325712
rect 128452 325660 128504 325712
rect 271420 325660 271472 325712
rect 271512 325660 271564 325712
rect 503996 323552 504048 323604
rect 504180 323552 504232 323604
rect 2964 322940 3016 322992
rect 5080 322940 5132 322992
rect 271512 322872 271564 322924
rect 271696 322872 271748 322924
rect 130016 321580 130068 321632
rect 580172 321580 580224 321632
rect 122564 321512 122616 321564
rect 122748 321512 122800 321564
rect 132684 321512 132736 321564
rect 132868 321512 132920 321564
rect 281264 321512 281316 321564
rect 281356 321512 281408 321564
rect 255780 318792 255832 318844
rect 255872 318792 255924 318844
rect 503536 318792 503588 318844
rect 503720 318792 503772 318844
rect 503996 318792 504048 318844
rect 504180 318792 504232 318844
rect 122472 318724 122524 318776
rect 122748 318724 122800 318776
rect 132408 318724 132460 318776
rect 132868 318724 132920 318776
rect 257712 318724 257764 318776
rect 257988 318724 258040 318776
rect 281080 318724 281132 318776
rect 281356 318724 281408 318776
rect 504364 318724 504416 318776
rect 504456 318724 504508 318776
rect 258172 317432 258224 317484
rect 258632 317432 258684 317484
rect 503444 313896 503496 313948
rect 503720 313896 503772 313948
rect 503628 311856 503680 311908
rect 503996 311856 504048 311908
rect 503628 311720 503680 311772
rect 503996 311720 504048 311772
rect 128728 311584 128780 311636
rect 129096 311584 129148 311636
rect 131764 310496 131816 310548
rect 580172 310496 580224 310548
rect 504364 309204 504416 309256
rect 504456 309204 504508 309256
rect 122472 309136 122524 309188
rect 122656 309136 122708 309188
rect 132408 309136 132460 309188
rect 132776 309136 132828 309188
rect 257712 309136 257764 309188
rect 257804 309136 257856 309188
rect 281080 309136 281132 309188
rect 281264 309136 281316 309188
rect 307024 309136 307076 309188
rect 503444 309136 503496 309188
rect 503812 309136 503864 309188
rect 307116 309068 307168 309120
rect 504180 309068 504232 309120
rect 504364 309068 504416 309120
rect 2964 307776 3016 307828
rect 5172 307776 5224 307828
rect 307116 307776 307168 307828
rect 307208 307776 307260 307828
rect 128728 307028 128780 307080
rect 129096 307028 129148 307080
rect 8024 306348 8076 306400
rect 8208 306348 8260 306400
rect 271788 303560 271840 303612
rect 271972 303560 272024 303612
rect 281264 302200 281316 302252
rect 281356 302132 281408 302184
rect 128636 299480 128688 299532
rect 128820 299480 128872 299532
rect 307024 299480 307076 299532
rect 307208 299480 307260 299532
rect 308680 299480 308732 299532
rect 308772 299480 308824 299532
rect 504180 299480 504232 299532
rect 504456 299480 504508 299532
rect 255504 299412 255556 299464
rect 255596 299412 255648 299464
rect 257712 299412 257764 299464
rect 257896 299412 257948 299464
rect 258264 299412 258316 299464
rect 258356 299412 258408 299464
rect 281080 299412 281132 299464
rect 281356 299412 281408 299464
rect 504456 298052 504508 298104
rect 504732 298052 504784 298104
rect 128728 297372 128780 297424
rect 129096 297372 129148 297424
rect 2964 293972 3016 294024
rect 434812 293972 434864 294024
rect 308680 292544 308732 292596
rect 308864 292544 308916 292596
rect 322848 291932 322900 291984
rect 378692 291932 378744 291984
rect 300768 291864 300820 291916
rect 378600 291864 378652 291916
rect 198924 291796 198976 291848
rect 231860 291796 231912 291848
rect 300676 291796 300728 291848
rect 378876 291796 378928 291848
rect 128452 290436 128504 290488
rect 128636 290436 128688 290488
rect 255504 289892 255556 289944
rect 258264 289892 258316 289944
rect 255596 289824 255648 289876
rect 257712 289824 257764 289876
rect 257804 289824 257856 289876
rect 258356 289824 258408 289876
rect 281080 289824 281132 289876
rect 281264 289824 281316 289876
rect 504548 288396 504600 288448
rect 504732 288396 504784 288448
rect 128728 287716 128780 287768
rect 129096 287716 129148 287768
rect 8024 287036 8076 287088
rect 8208 287036 8260 287088
rect 271788 284248 271840 284300
rect 271972 284248 272024 284300
rect 308588 283568 308640 283620
rect 308864 283568 308916 283620
rect 503720 283024 503772 283076
rect 503812 282956 503864 283008
rect 132684 282888 132736 282940
rect 132868 282888 132920 282940
rect 257804 282888 257856 282940
rect 257988 282888 258040 282940
rect 281264 282888 281316 282940
rect 281356 282820 281408 282872
rect 128452 280100 128504 280152
rect 128636 280100 128688 280152
rect 281356 280100 281408 280152
rect 281632 280100 281684 280152
rect 308588 278740 308640 278792
rect 308680 278740 308732 278792
rect 504456 278672 504508 278724
rect 504548 278672 504600 278724
rect 258264 275952 258316 276004
rect 258356 275952 258408 276004
rect 131580 274660 131632 274712
rect 579988 274660 580040 274712
rect 128728 274252 128780 274304
rect 129096 274252 129148 274304
rect 503628 273300 503680 273352
rect 503996 273300 504048 273352
rect 503628 273164 503680 273216
rect 503996 273164 504048 273216
rect 281356 270580 281408 270632
rect 281632 270580 281684 270632
rect 128452 270512 128504 270564
rect 128636 270512 128688 270564
rect 307024 270512 307076 270564
rect 281080 270444 281132 270496
rect 281356 270444 281408 270496
rect 306932 270444 306984 270496
rect 308680 269084 308732 269136
rect 308864 269084 308916 269136
rect 306748 269016 306800 269068
rect 306932 269016 306984 269068
rect 128728 268404 128780 268456
rect 129096 268404 129148 268456
rect 8024 267724 8076 267776
rect 8208 267724 8260 267776
rect 2872 264936 2924 264988
rect 5264 264936 5316 264988
rect 271604 264868 271656 264920
rect 271788 264868 271840 264920
rect 503720 263644 503772 263696
rect 503996 263644 504048 263696
rect 131672 263576 131724 263628
rect 580172 263576 580224 263628
rect 503720 263508 503772 263560
rect 503996 263508 504048 263560
rect 255688 260856 255740 260908
rect 281080 260856 281132 260908
rect 281264 260856 281316 260908
rect 128084 260788 128136 260840
rect 128544 260788 128596 260840
rect 504272 260788 504324 260840
rect 504548 260788 504600 260840
rect 255688 260720 255740 260772
rect 306748 259428 306800 259480
rect 307024 259428 307076 259480
rect 128728 258748 128780 258800
rect 129096 258748 129148 258800
rect 271420 255212 271472 255264
rect 271788 255212 271840 255264
rect 503628 253988 503680 254040
rect 503996 253988 504048 254040
rect 503628 253852 503680 253904
rect 503996 253852 504048 253904
rect 504272 253784 504324 253836
rect 504548 253784 504600 253836
rect 307024 251472 307076 251524
rect 307024 251336 307076 251388
rect 2872 251200 2924 251252
rect 434904 251200 434956 251252
rect 7748 251132 7800 251184
rect 7932 251132 7984 251184
rect 504088 251132 504140 251184
rect 504272 251132 504324 251184
rect 128728 249092 128780 249144
rect 129096 249092 129148 249144
rect 258448 249092 258500 249144
rect 258448 248956 258500 249008
rect 271420 245624 271472 245676
rect 271512 245624 271564 245676
rect 308588 245352 308640 245404
rect 308864 245352 308916 245404
rect 503720 244400 503772 244452
rect 503812 244332 503864 244384
rect 271512 242156 271564 242208
rect 271788 242156 271840 242208
rect 307024 241544 307076 241596
rect 307208 241544 307260 241596
rect 7748 241476 7800 241528
rect 8024 241476 8076 241528
rect 281080 241476 281132 241528
rect 281264 241476 281316 241528
rect 504088 241476 504140 241528
rect 504456 241476 504508 241528
rect 281080 241340 281132 241392
rect 281264 241340 281316 241392
rect 258264 240116 258316 240168
rect 258448 240116 258500 240168
rect 128728 239436 128780 239488
rect 129096 239436 129148 239488
rect 258264 238688 258316 238740
rect 258448 238688 258500 238740
rect 255412 236648 255464 236700
rect 255596 236648 255648 236700
rect 308588 235288 308640 235340
rect 308772 235288 308824 235340
rect 8024 234676 8076 234728
rect 503628 234676 503680 234728
rect 503996 234676 504048 234728
rect 504456 234676 504508 234728
rect 7932 234540 7984 234592
rect 503628 234540 503680 234592
rect 503996 234540 504048 234592
rect 504364 234540 504416 234592
rect 128636 231820 128688 231872
rect 128820 231820 128872 231872
rect 257988 231820 258040 231872
rect 258172 231820 258224 231872
rect 281080 231820 281132 231872
rect 281264 231820 281316 231872
rect 306932 231820 306984 231872
rect 7748 231752 7800 231804
rect 7932 231752 7984 231804
rect 307024 231752 307076 231804
rect 504180 231752 504232 231804
rect 504364 231752 504416 231804
rect 306932 230460 306984 230512
rect 307024 230460 307076 230512
rect 128728 229712 128780 229764
rect 129096 229712 129148 229764
rect 132684 227740 132736 227792
rect 580080 227740 580132 227792
rect 271696 227672 271748 227724
rect 271880 227672 271932 227724
rect 503720 225088 503772 225140
rect 503812 225020 503864 225072
rect 122564 224884 122616 224936
rect 122748 224884 122800 224936
rect 2780 222504 2832 222556
rect 6184 222504 6236 222556
rect 7748 222164 7800 222216
rect 8024 222164 8076 222216
rect 255596 222164 255648 222216
rect 255688 222164 255740 222216
rect 281080 222164 281132 222216
rect 281172 222164 281224 222216
rect 308680 222164 308732 222216
rect 504180 222164 504232 222216
rect 504456 222164 504508 222216
rect 213920 222096 213972 222148
rect 214196 222096 214248 222148
rect 307024 222096 307076 222148
rect 307116 222096 307168 222148
rect 308772 222096 308824 222148
rect 308680 220804 308732 220856
rect 308772 220804 308824 220856
rect 128728 220056 128780 220108
rect 129096 220056 129148 220108
rect 271696 218016 271748 218068
rect 271972 218016 272024 218068
rect 132776 216656 132828 216708
rect 579804 216656 579856 216708
rect 308312 215976 308364 216028
rect 308680 215976 308732 216028
rect 8024 215364 8076 215416
rect 122748 215364 122800 215416
rect 128452 215364 128504 215416
rect 258540 215364 258592 215416
rect 503628 215364 503680 215416
rect 503996 215364 504048 215416
rect 281172 215296 281224 215348
rect 7932 215228 7984 215280
rect 122656 215228 122708 215280
rect 128452 215228 128504 215280
rect 258448 215228 258500 215280
rect 504456 215364 504508 215416
rect 297272 215228 297324 215280
rect 298008 215228 298060 215280
rect 503628 215228 503680 215280
rect 503996 215228 504048 215280
rect 504272 215228 504324 215280
rect 281264 215160 281316 215212
rect 214196 212508 214248 212560
rect 214380 212508 214432 212560
rect 255596 212508 255648 212560
rect 255688 212508 255740 212560
rect 257804 212508 257856 212560
rect 257988 212508 258040 212560
rect 271512 212508 271564 212560
rect 271972 212508 272024 212560
rect 275652 212508 275704 212560
rect 275928 212508 275980 212560
rect 307024 212508 307076 212560
rect 307208 212508 307260 212560
rect 255596 211488 255648 211540
rect 256148 211488 256200 211540
rect 297824 211080 297876 211132
rect 303896 211080 303948 211132
rect 2780 210400 2832 210452
rect 3056 210400 3108 210452
rect 128728 210400 128780 210452
rect 129096 210400 129148 210452
rect 132868 210400 132920 210452
rect 133512 210400 133564 210452
rect 268476 210400 268528 210452
rect 268844 210400 268896 210452
rect 290924 210400 290976 210452
rect 291108 210400 291160 210452
rect 297732 210400 297784 210452
rect 311992 210400 312044 210452
rect 3056 207000 3108 207052
rect 434996 207000 435048 207052
rect 503720 205776 503772 205828
rect 503812 205708 503864 205760
rect 297272 205640 297324 205692
rect 297824 205640 297876 205692
rect 503720 205640 503772 205692
rect 503996 205640 504048 205692
rect 504180 205640 504232 205692
rect 8024 205572 8076 205624
rect 308404 205572 308456 205624
rect 308588 205572 308640 205624
rect 504272 205572 504324 205624
rect 8116 205504 8168 205556
rect 196624 205096 196676 205148
rect 230572 205096 230624 205148
rect 195152 205028 195204 205080
rect 229560 205028 229612 205080
rect 195244 204960 195296 205012
rect 231216 204960 231268 205012
rect 294880 204960 294932 205012
rect 378324 204960 378376 205012
rect 196532 204892 196584 204944
rect 233240 204892 233292 204944
rect 237472 204892 237524 204944
rect 237748 204892 237800 204944
rect 286232 204892 286284 204944
rect 378232 204892 378284 204944
rect 199476 204212 199528 204264
rect 244740 204212 244792 204264
rect 255780 204212 255832 204264
rect 266912 204212 266964 204264
rect 319168 204212 319220 204264
rect 380072 204212 380124 204264
rect 197636 204144 197688 204196
rect 245660 204144 245712 204196
rect 250536 204144 250588 204196
rect 267832 204144 267884 204196
rect 313556 204144 313608 204196
rect 378140 204144 378192 204196
rect 197452 204076 197504 204128
rect 251916 204076 251968 204128
rect 253572 204076 253624 204128
rect 268660 204076 268712 204128
rect 314936 204076 314988 204128
rect 380164 204076 380216 204128
rect 199384 204008 199436 204060
rect 254032 204008 254084 204060
rect 255964 204008 256016 204060
rect 268384 204008 268436 204060
rect 308404 204008 308456 204060
rect 377220 204008 377272 204060
rect 199200 203940 199252 203992
rect 258448 203940 258500 203992
rect 306656 203940 306708 203992
rect 380716 203940 380768 203992
rect 197728 203872 197780 203924
rect 257160 203872 257212 203924
rect 259828 203872 259880 203924
rect 267188 203872 267240 203924
rect 301412 203872 301464 203924
rect 379520 203872 379572 203924
rect 197912 203804 197964 203856
rect 260380 203804 260432 203856
rect 299388 203804 299440 203856
rect 380256 203804 380308 203856
rect 198188 203736 198240 203788
rect 262772 203736 262824 203788
rect 292488 203736 292540 203788
rect 379796 203736 379848 203788
rect 197544 203668 197596 203720
rect 262956 203668 263008 203720
rect 287520 203668 287572 203720
rect 379612 203668 379664 203720
rect 197820 203600 197872 203652
rect 265440 203600 265492 203652
rect 271788 203600 271840 203652
rect 369860 203600 369912 203652
rect 198004 203532 198056 203584
rect 267188 203532 267240 203584
rect 280528 203532 280580 203584
rect 379888 203532 379940 203584
rect 198096 203464 198148 203516
rect 238760 203464 238812 203516
rect 240968 203464 241020 203516
rect 268568 203464 268620 203516
rect 296168 203464 296220 203516
rect 353300 203464 353352 203516
rect 209688 203396 209740 203448
rect 243176 203396 243228 203448
rect 294420 203396 294472 203448
rect 340880 203396 340932 203448
rect 198372 203328 198424 203380
rect 225144 203328 225196 203380
rect 302884 203328 302936 203380
rect 331220 203328 331272 203380
rect 297916 203260 297968 203312
rect 325148 203260 325200 203312
rect 315212 203192 315264 203244
rect 336004 203192 336056 203244
rect 308956 203124 309008 203176
rect 321744 203124 321796 203176
rect 128452 202852 128504 202904
rect 128636 202852 128688 202904
rect 196716 202784 196768 202836
rect 195336 202716 195388 202768
rect 220636 202716 220688 202768
rect 220820 202784 220872 202836
rect 221280 202784 221332 202836
rect 239680 202784 239732 202836
rect 240140 202784 240192 202836
rect 240508 202784 240560 202836
rect 242164 202784 242216 202836
rect 242256 202784 242308 202836
rect 242808 202784 242860 202836
rect 251456 202784 251508 202836
rect 258816 202852 258868 202904
rect 504180 202852 504232 202904
rect 504272 202852 504324 202904
rect 226892 202716 226944 202768
rect 236368 202716 236420 202768
rect 259000 202784 259052 202836
rect 260104 202784 260156 202836
rect 263600 202784 263652 202836
rect 266268 202784 266320 202836
rect 269396 202784 269448 202836
rect 289268 202784 289320 202836
rect 289728 202784 289780 202836
rect 290556 202784 290608 202836
rect 291016 202784 291068 202836
rect 291384 202784 291436 202836
rect 292396 202784 292448 202836
rect 293132 202784 293184 202836
rect 293868 202784 293920 202836
rect 295800 202784 295852 202836
rect 296444 202784 296496 202836
rect 300124 202784 300176 202836
rect 300676 202784 300728 202836
rect 258724 202716 258776 202768
rect 263876 202716 263928 202768
rect 264888 202716 264940 202768
rect 269488 202716 269540 202768
rect 299480 202716 299532 202768
rect 307116 202784 307168 202836
rect 311900 202784 311952 202836
rect 312544 202784 312596 202836
rect 312636 202784 312688 202836
rect 319168 202784 319220 202836
rect 319260 202784 319312 202836
rect 320088 202784 320140 202836
rect 351000 202784 351052 202836
rect 351828 202784 351880 202836
rect 352748 202784 352800 202836
rect 353208 202784 353260 202836
rect 353300 202784 353352 202836
rect 413008 202784 413060 202836
rect 413100 202784 413152 202836
rect 414664 202784 414716 202836
rect 415032 202784 415084 202836
rect 417424 202784 417476 202836
rect 417516 202784 417568 202836
rect 418068 202784 418120 202836
rect 301044 202716 301096 202768
rect 307208 202716 307260 202768
rect 310428 202716 310480 202768
rect 375656 202716 375708 202768
rect 375748 202716 375800 202768
rect 378784 202716 378836 202768
rect 400588 202716 400640 202768
rect 401508 202716 401560 202768
rect 401600 202716 401652 202768
rect 458824 202716 458876 202768
rect 200028 202648 200080 202700
rect 238208 202648 238260 202700
rect 240784 202648 240836 202700
rect 242348 202648 242400 202700
rect 250904 202648 250956 202700
rect 269212 202648 269264 202700
rect 299112 202648 299164 202700
rect 305000 202648 305052 202700
rect 306932 202648 306984 202700
rect 320640 202648 320692 202700
rect 344008 202648 344060 202700
rect 156604 202580 156656 202632
rect 169116 202580 169168 202632
rect 198280 202580 198332 202632
rect 202880 202580 202932 202632
rect 207664 202580 207716 202632
rect 239312 202580 239364 202632
rect 239404 202580 239456 202632
rect 243820 202580 243872 202632
rect 248972 202580 249024 202632
rect 268108 202580 268160 202632
rect 283932 202580 283984 202632
rect 284208 202580 284260 202632
rect 299020 202580 299072 202632
rect 305644 202580 305696 202632
rect 307208 202580 307260 202632
rect 309508 202580 309560 202632
rect 311164 202580 311216 202632
rect 331864 202580 331916 202632
rect 342076 202580 342128 202632
rect 153844 202512 153896 202564
rect 178040 202512 178092 202564
rect 196992 202512 197044 202564
rect 241520 202512 241572 202564
rect 247500 202512 247552 202564
rect 130108 202444 130160 202496
rect 134432 202444 134484 202496
rect 152464 202444 152516 202496
rect 176936 202444 176988 202496
rect 195520 202444 195572 202496
rect 241060 202444 241112 202496
rect 243728 202444 243780 202496
rect 252652 202444 252704 202496
rect 253848 202512 253900 202564
rect 267924 202512 267976 202564
rect 299296 202512 299348 202564
rect 302240 202512 302292 202564
rect 302332 202512 302384 202564
rect 302976 202512 303028 202564
rect 307300 202512 307352 202564
rect 325700 202512 325752 202564
rect 151084 202376 151136 202428
rect 182180 202376 182232 202428
rect 199936 202376 199988 202428
rect 246488 202376 246540 202428
rect 137284 202308 137336 202360
rect 168380 202308 168432 202360
rect 195612 202308 195664 202360
rect 245200 202308 245252 202360
rect 247592 202308 247644 202360
rect 253480 202308 253532 202360
rect 254124 202444 254176 202496
rect 266268 202444 266320 202496
rect 267648 202444 267700 202496
rect 269304 202444 269356 202496
rect 273996 202444 274048 202496
rect 274548 202444 274600 202496
rect 280988 202444 281040 202496
rect 281264 202444 281316 202496
rect 282276 202444 282328 202496
rect 282736 202444 282788 202496
rect 288808 202444 288860 202496
rect 315304 202444 315356 202496
rect 333152 202444 333204 202496
rect 333888 202444 333940 202496
rect 341432 202444 341484 202496
rect 342168 202444 342220 202496
rect 343180 202444 343232 202496
rect 343548 202444 343600 202496
rect 346676 202444 346728 202496
rect 347596 202444 347648 202496
rect 349988 202648 350040 202700
rect 350448 202648 350500 202700
rect 351736 202648 351788 202700
rect 353300 202648 353352 202700
rect 348332 202580 348384 202632
rect 412916 202648 412968 202700
rect 413008 202648 413060 202700
rect 417332 202648 417384 202700
rect 353484 202580 353536 202632
rect 417148 202580 417200 202632
rect 416872 202512 416924 202564
rect 412824 202444 412876 202496
rect 412916 202444 412968 202496
rect 417240 202444 417292 202496
rect 253940 202376 253992 202428
rect 268016 202376 268068 202428
rect 299204 202376 299256 202428
rect 306932 202376 306984 202428
rect 307024 202376 307076 202428
rect 307576 202376 307628 202428
rect 310520 202376 310572 202428
rect 311256 202376 311308 202428
rect 311348 202376 311400 202428
rect 325700 202376 325752 202428
rect 332508 202376 332560 202428
rect 415032 202376 415084 202428
rect 415768 202376 415820 202428
rect 416688 202376 416740 202428
rect 266084 202308 266136 202360
rect 266176 202308 266228 202360
rect 269580 202308 269632 202360
rect 297548 202308 297600 202360
rect 302240 202308 302292 202360
rect 305552 202308 305604 202360
rect 140044 202240 140096 202292
rect 178684 202240 178736 202292
rect 201408 202240 201460 202292
rect 258540 202240 258592 202292
rect 103428 202172 103480 202224
rect 142528 202172 142580 202224
rect 144184 202172 144236 202224
rect 181260 202172 181312 202224
rect 199108 202172 199160 202224
rect 256516 202172 256568 202224
rect 93768 202104 93820 202156
rect 134708 202104 134760 202156
rect 141424 202104 141476 202156
rect 180340 202104 180392 202156
rect 199292 202104 199344 202156
rect 269764 202240 269816 202292
rect 292304 202240 292356 202292
rect 375656 202308 375708 202360
rect 377312 202308 377364 202360
rect 410156 202308 410208 202360
rect 411168 202308 411220 202360
rect 417148 202308 417200 202360
rect 503904 202308 503956 202360
rect 259000 202172 259052 202224
rect 266728 202172 266780 202224
rect 270960 202172 271012 202224
rect 374368 202172 374420 202224
rect 374460 202172 374512 202224
rect 375288 202172 375340 202224
rect 378508 202240 378560 202292
rect 411076 202240 411128 202292
rect 503812 202240 503864 202292
rect 379704 202172 379756 202224
rect 409236 202172 409288 202224
rect 503720 202172 503772 202224
rect 258908 202104 258960 202156
rect 268292 202104 268344 202156
rect 283564 202104 283616 202156
rect 196900 202036 196952 202088
rect 216864 202036 216916 202088
rect 217968 202036 218020 202088
rect 195428 201968 195480 202020
rect 223028 201968 223080 202020
rect 195888 201900 195940 201952
rect 218060 201900 218112 201952
rect 220636 201900 220688 201952
rect 227812 201900 227864 201952
rect 199660 201832 199712 201884
rect 219532 201832 219584 201884
rect 196808 201764 196860 201816
rect 218612 201764 218664 201816
rect 239220 202036 239272 202088
rect 240048 202036 240100 202088
rect 251824 202036 251876 202088
rect 267740 202036 267792 202088
rect 297456 202036 297508 202088
rect 303896 202036 303948 202088
rect 306932 202036 306984 202088
rect 315304 202036 315356 202088
rect 246304 201968 246356 202020
rect 243084 201900 243136 201952
rect 247684 201900 247736 201952
rect 253112 201968 253164 202020
rect 253664 201968 253716 202020
rect 253756 201968 253808 202020
rect 258724 201968 258776 202020
rect 258816 201968 258868 202020
rect 266452 201968 266504 202020
rect 300492 201968 300544 202020
rect 317144 201968 317196 202020
rect 320548 201968 320600 202020
rect 321468 201968 321520 202020
rect 324044 201968 324096 202020
rect 324964 201968 325016 202020
rect 345756 202104 345808 202156
rect 353484 202104 353536 202156
rect 353576 202104 353628 202156
rect 354588 202104 354640 202156
rect 364892 202104 364944 202156
rect 365536 202104 365588 202156
rect 366180 202104 366232 202156
rect 367008 202104 367060 202156
rect 376484 202104 376536 202156
rect 505744 202104 505796 202156
rect 357900 202036 357952 202088
rect 334624 201968 334676 202020
rect 366916 201968 366968 202020
rect 414664 201968 414716 202020
rect 414940 202036 414992 202088
rect 417148 202036 417200 202088
rect 416964 201968 417016 202020
rect 260840 201900 260892 201952
rect 265348 201900 265400 201952
rect 266820 201900 266872 201952
rect 267004 201900 267056 201952
rect 268200 201900 268252 201952
rect 299204 201900 299256 201952
rect 304264 201900 304316 201952
rect 239312 201832 239364 201884
rect 247776 201832 247828 201884
rect 257068 201832 257120 201884
rect 265992 201832 266044 201884
rect 266084 201832 266136 201884
rect 270684 201832 270736 201884
rect 297272 201832 297324 201884
rect 305552 201832 305604 201884
rect 246028 201764 246080 201816
rect 256516 201764 256568 201816
rect 259920 201764 259972 201816
rect 198740 201696 198792 201748
rect 216036 201696 216088 201748
rect 250076 201696 250128 201748
rect 250996 201696 251048 201748
rect 254860 201696 254912 201748
rect 266452 201764 266504 201816
rect 262680 201696 262732 201748
rect 265900 201696 265952 201748
rect 265992 201696 266044 201748
rect 270868 201764 270920 201816
rect 300400 201764 300452 201816
rect 315580 201900 315632 201952
rect 374368 201900 374420 201952
rect 379980 201900 380032 201952
rect 412272 201900 412324 201952
rect 457444 201900 457496 201952
rect 412824 201832 412876 201884
rect 417056 201832 417108 201884
rect 307116 201764 307168 201816
rect 313648 201764 313700 201816
rect 414664 201764 414716 201816
rect 418804 201764 418856 201816
rect 268108 201696 268160 201748
rect 270592 201696 270644 201748
rect 272248 201696 272300 201748
rect 273168 201696 273220 201748
rect 273628 201696 273680 201748
rect 274456 201696 274508 201748
rect 275284 201696 275336 201748
rect 275836 201696 275888 201748
rect 279240 201696 279292 201748
rect 280068 201696 280120 201748
rect 298376 201696 298428 201748
rect 301044 201696 301096 201748
rect 198556 201628 198608 201680
rect 212540 201628 212592 201680
rect 244648 201628 244700 201680
rect 253848 201628 253900 201680
rect 258356 201628 258408 201680
rect 266728 201628 266780 201680
rect 127624 201560 127676 201612
rect 134156 201560 134208 201612
rect 198464 201560 198516 201612
rect 211160 201560 211212 201612
rect 258724 201560 258776 201612
rect 266360 201560 266412 201612
rect 270776 201628 270828 201680
rect 297364 201628 297416 201680
rect 311348 201696 311400 201748
rect 301872 201628 301924 201680
rect 312636 201628 312688 201680
rect 198832 201492 198884 201544
rect 211712 201492 211764 201544
rect 8024 201424 8076 201476
rect 8116 201424 8168 201476
rect 252744 201424 252796 201476
rect 266452 201492 266504 201544
rect 265900 201424 265952 201476
rect 267096 201560 267148 201612
rect 270500 201560 270552 201612
rect 298744 201560 298796 201612
rect 307300 201560 307352 201612
rect 266636 201492 266688 201544
rect 268016 201492 268068 201544
rect 297640 201492 297692 201544
rect 306932 201492 306984 201544
rect 355324 201492 355376 201544
rect 355968 201492 356020 201544
rect 359648 201492 359700 201544
rect 360108 201492 360160 201544
rect 360568 201492 360620 201544
rect 361396 201492 361448 201544
rect 362316 201492 362368 201544
rect 362776 201492 362828 201544
rect 400956 201492 401008 201544
rect 401508 201492 401560 201544
rect 504180 201220 504232 201272
rect 504456 201220 504508 201272
rect 4068 201152 4120 201204
rect 436652 201152 436704 201204
rect 3884 201084 3936 201136
rect 436560 201084 436612 201136
rect 2780 201016 2832 201068
rect 436744 201016 436796 201068
rect 132408 200948 132460 201000
rect 580724 200948 580776 201000
rect 131304 200880 131356 200932
rect 580356 200880 580408 200932
rect 131396 200812 131448 200864
rect 580632 200812 580684 200864
rect 131488 200744 131540 200796
rect 580908 200744 580960 200796
rect 248696 200200 248748 200252
rect 249386 200200 249438 200252
rect 254998 200200 255050 200252
rect 258908 200200 258960 200252
rect 308542 200200 308594 200252
rect 308772 200200 308824 200252
rect 133788 200132 133840 200184
rect 579988 200132 580040 200184
rect 133512 200064 133564 200116
rect 135260 200064 135312 200116
rect 238760 199860 238812 199912
rect 239496 199860 239548 199912
rect 2780 199792 2832 199844
rect 436284 199792 436336 199844
rect 3884 198704 3936 198756
rect 131212 198704 131264 198756
rect 4068 197344 4120 197396
rect 131212 197344 131264 197396
rect 131304 196324 131356 196376
rect 14464 196052 14516 196104
rect 5356 195984 5408 196036
rect 131212 195984 131264 196036
rect 122748 195848 122800 195900
rect 122932 195848 122984 195900
rect 128360 195848 128412 195900
rect 128544 195848 128596 195900
rect 128728 195576 128780 195628
rect 129096 195576 129148 195628
rect 8944 194556 8996 194608
rect 131212 194556 131264 194608
rect 6184 194420 6236 194472
rect 131212 194420 131264 194472
rect 5172 193128 5224 193180
rect 5264 193060 5316 193112
rect 131212 193060 131264 193112
rect 131212 192788 131264 192840
rect 436284 192924 436336 192976
rect 436836 192924 436888 192976
rect 4988 191768 5040 191820
rect 131212 191768 131264 191820
rect 128728 191088 128780 191140
rect 129096 191088 129148 191140
rect 3240 190408 3292 190460
rect 131212 190408 131264 190460
rect 133512 189864 133564 189916
rect 133512 189728 133564 189780
rect 133788 189728 133840 189780
rect 133788 189592 133840 189644
rect 4896 188980 4948 189032
rect 131212 188980 131264 189032
rect 4804 188844 4856 188896
rect 9680 188844 9732 188896
rect 19248 188844 19300 188896
rect 22100 188844 22152 188896
rect 22192 188844 22244 188896
rect 41512 188708 41564 188760
rect 60740 188708 60792 188760
rect 67640 188776 67692 188828
rect 77208 188708 77260 188760
rect 79968 188708 80020 188760
rect 80060 188708 80112 188760
rect 86960 188776 87012 188828
rect 115940 188776 115992 188828
rect 41328 188640 41380 188692
rect 48320 188640 48372 188692
rect 57888 188640 57940 188692
rect 60648 188640 60700 188692
rect 96528 188640 96580 188692
rect 99380 188640 99432 188692
rect 99472 188640 99524 188692
rect 125508 188708 125560 188760
rect 131212 188572 131264 188624
rect 48320 188504 48372 188556
rect 57888 188504 57940 188556
rect 3700 187620 3752 187672
rect 131212 187620 131264 187672
rect 3516 186260 3568 186312
rect 131212 186260 131264 186312
rect 132868 185172 132920 185224
rect 133144 185172 133196 185224
rect 132868 184968 132920 185020
rect 133052 184968 133104 185020
rect 8300 184832 8352 184884
rect 131212 184832 131264 184884
rect 128360 183540 128412 183592
rect 128544 183540 128596 183592
rect 72424 183472 72476 183524
rect 131212 183472 131264 183524
rect 132592 181228 132644 181280
rect 133236 181228 133288 181280
rect 3700 179460 3752 179512
rect 8944 179460 8996 179512
rect 128728 177352 128780 177404
rect 129096 177352 129148 177404
rect 122748 176672 122800 176724
rect 128544 176672 128596 176724
rect 122656 176536 122708 176588
rect 128636 176536 128688 176588
rect 128728 175584 128780 175636
rect 129096 175584 129148 175636
rect 129648 175176 129700 175228
rect 131212 175176 131264 175228
rect 129556 175108 129608 175160
rect 132040 175108 132092 175160
rect 504456 173884 504508 173936
rect 504640 173884 504692 173936
rect 128360 169056 128412 169108
rect 128544 169056 128596 169108
rect 133052 168648 133104 168700
rect 133052 168444 133104 168496
rect 130016 166812 130068 166864
rect 132040 166812 132092 166864
rect 504180 164160 504232 164212
rect 504364 164160 504416 164212
rect 128728 162120 128780 162172
rect 129096 162120 129148 162172
rect 122564 161440 122616 161492
rect 122748 161440 122800 161492
rect 4804 158720 4856 158772
rect 131212 158720 131264 158772
rect 4160 155932 4212 155984
rect 131212 155932 131264 155984
rect 3056 155864 3108 155916
rect 131212 155796 131264 155848
rect 436100 155592 436152 155644
rect 438124 155592 438176 155644
rect 2872 154504 2924 154556
rect 131212 154504 131264 154556
rect 2964 153144 3016 153196
rect 131212 153144 131264 153196
rect 5080 153076 5132 153128
rect 6920 153076 6972 153128
rect 82820 153076 82872 153128
rect 82912 153076 82964 153128
rect 16488 152940 16540 152992
rect 116308 152940 116360 152992
rect 116308 152804 116360 152856
rect 131212 152804 131264 152856
rect 437388 151920 437440 151972
rect 442264 151920 442316 151972
rect 3148 151716 3200 151768
rect 131212 151716 131264 151768
rect 3332 150356 3384 150408
rect 131212 150356 131264 150408
rect 437020 150288 437072 150340
rect 440884 150288 440936 150340
rect 128728 149812 128780 149864
rect 129096 149812 129148 149864
rect 3976 148996 4028 149048
rect 131212 148996 131264 149048
rect 115940 148860 115992 148912
rect 436192 148860 436244 148912
rect 439504 148860 439556 148912
rect 70400 148792 70452 148844
rect 22192 148724 22244 148776
rect 41512 148724 41564 148776
rect 50988 148724 51040 148776
rect 56600 148724 56652 148776
rect 64880 148724 64932 148776
rect 79968 148724 80020 148776
rect 80060 148724 80112 148776
rect 84200 148792 84252 148844
rect 3792 148656 3844 148708
rect 22008 148656 22060 148708
rect 26240 148656 26292 148708
rect 35808 148656 35860 148708
rect 41328 148656 41380 148708
rect 51080 148656 51132 148708
rect 56508 148656 56560 148708
rect 93768 148656 93820 148708
rect 99380 148656 99432 148708
rect 99472 148656 99524 148708
rect 116032 148588 116084 148640
rect 131212 148588 131264 148640
rect 26240 148520 26292 148572
rect 35808 148520 35860 148572
rect 130936 148180 130988 148232
rect 131212 148180 131264 148232
rect 3608 147568 3660 147620
rect 132224 147568 132276 147620
rect 132316 147568 132368 147620
rect 122564 147500 122616 147552
rect 122748 147500 122800 147552
rect 132224 146548 132276 146600
rect 130936 146344 130988 146396
rect 131120 146344 131172 146396
rect 3424 146208 3476 146260
rect 131120 146208 131172 146260
rect 436100 146208 436152 146260
rect 438216 146208 438268 146260
rect 24768 144848 24820 144900
rect 131120 144848 131172 144900
rect 437388 144848 437440 144900
rect 580264 144848 580316 144900
rect 131028 144440 131080 144492
rect 131028 144100 131080 144152
rect 128820 143488 128872 143540
rect 129096 143488 129148 143540
rect 436100 142060 436152 142112
rect 438308 142060 438360 142112
rect 437388 140700 437440 140752
rect 580448 140700 580500 140752
rect 122564 137980 122616 138032
rect 437388 137912 437440 137964
rect 580540 137912 580592 137964
rect 122656 137844 122708 137896
rect 437020 136552 437072 136604
rect 504456 136552 504508 136604
rect 2780 136348 2832 136400
rect 5356 136348 5408 136400
rect 128636 135192 128688 135244
rect 128728 135192 128780 135244
rect 128820 135192 128872 135244
rect 129096 135192 129148 135244
rect 132868 135192 132920 135244
rect 132960 135124 133012 135176
rect 437388 133832 437440 133884
rect 580816 133832 580868 133884
rect 436836 132404 436888 132456
rect 580172 132404 580224 132456
rect 128820 130364 128872 130416
rect 129096 130364 129148 130416
rect 437388 129684 437440 129736
rect 580080 129684 580132 129736
rect 128728 128324 128780 128376
rect 128636 128256 128688 128308
rect 436100 128256 436152 128308
rect 580632 128256 580684 128308
rect 128728 125536 128780 125588
rect 128820 125536 128872 125588
rect 129096 125536 129148 125588
rect 129188 125536 129240 125588
rect 129096 125400 129148 125452
rect 129188 125400 129240 125452
rect 134064 120776 134116 120828
rect 580908 120776 580960 120828
rect 133972 120708 134024 120760
rect 580356 120708 580408 120760
rect 132408 120640 132460 120692
rect 580264 120640 580316 120692
rect 3240 120572 3292 120624
rect 436468 120572 436520 120624
rect 187792 119756 187844 119808
rect 188758 119756 188810 119808
rect 205180 119756 205232 119808
rect 210194 119756 210246 119808
rect 130200 119348 130252 119400
rect 139400 119348 139452 119400
rect 143632 119348 143684 119400
rect 144368 119348 144420 119400
rect 130844 119076 130896 119128
rect 142252 119076 142304 119128
rect 142528 119076 142580 119128
rect 137192 118940 137244 118992
rect 138296 118940 138348 118992
rect 129464 118872 129516 118924
rect 145012 118872 145064 118924
rect 131028 118804 131080 118856
rect 147772 118804 147824 118856
rect 129372 118736 129424 118788
rect 149060 118736 149112 118788
rect 128268 118668 128320 118720
rect 154672 118668 154724 118720
rect 155316 118668 155368 118720
rect 69848 118600 69900 118652
rect 70308 118600 70360 118652
rect 138204 118600 138256 118652
rect 138296 118600 138348 118652
rect 143080 118600 143132 118652
rect 146760 118600 146812 118652
rect 157340 118600 157392 118652
rect 170404 118600 170456 118652
rect 198188 118600 198240 118652
rect 200028 118600 200080 118652
rect 236184 118600 236236 118652
rect 239404 118600 239456 118652
rect 249800 118600 249852 118652
rect 249892 118600 249944 118652
rect 258264 118600 258316 118652
rect 298652 118600 298704 118652
rect 318984 118600 319036 118652
rect 349436 118600 349488 118652
rect 416964 118600 417016 118652
rect 424784 118600 424836 118652
rect 493324 118600 493376 118652
rect 97908 118532 97960 118584
rect 181076 118532 181128 118584
rect 195888 118532 195940 118584
rect 234712 118532 234764 118584
rect 240048 118532 240100 118584
rect 256976 118532 257028 118584
rect 301136 118532 301188 118584
rect 323124 118532 323176 118584
rect 364064 118532 364116 118584
rect 380164 118532 380216 118584
rect 408224 118532 408276 118584
rect 478144 118532 478196 118584
rect 82728 118464 82780 118516
rect 164516 118464 164568 118516
rect 188988 118464 189040 118516
rect 230664 118464 230716 118516
rect 237288 118464 237340 118516
rect 255320 118464 255372 118516
rect 299296 118464 299348 118516
rect 320364 118464 320416 118516
rect 342168 118464 342220 118516
rect 400956 118464 401008 118516
rect 404268 118464 404320 118516
rect 475384 118464 475436 118516
rect 120724 118396 120776 118448
rect 125692 118396 125744 118448
rect 170036 118396 170088 118448
rect 186228 118396 186280 118448
rect 229468 118396 229520 118448
rect 235908 118396 235960 118448
rect 254584 118396 254636 118448
rect 302148 118396 302200 118448
rect 325884 118396 325936 118448
rect 336004 118396 336056 118448
rect 348424 118396 348476 118448
rect 369676 118396 369728 118448
rect 374644 118396 374696 118448
rect 417424 118396 417476 118448
rect 422852 118396 422904 118448
rect 431776 118396 431828 118448
rect 500224 118396 500276 118448
rect 71596 118328 71648 118380
rect 88340 118328 88392 118380
rect 110328 118328 110380 118380
rect 145564 118328 145616 118380
rect 146852 118328 146904 118380
rect 153476 118328 153528 118380
rect 182180 118328 182232 118380
rect 187792 118328 187844 118380
rect 194508 118328 194560 118380
rect 233240 118328 233292 118380
rect 56508 118260 56560 118312
rect 125876 118260 125928 118312
rect 126888 118260 126940 118312
rect 128912 118260 128964 118312
rect 135444 118260 135496 118312
rect 137192 118260 137244 118312
rect 137284 118260 137336 118312
rect 182916 118260 182968 118312
rect 183468 118260 183520 118312
rect 227720 118260 227772 118312
rect 231124 118260 231176 118312
rect 238116 118328 238168 118380
rect 238668 118328 238720 118380
rect 256700 118328 256752 118380
rect 260748 118328 260800 118380
rect 267740 118328 267792 118380
rect 304172 118328 304224 118380
rect 330024 118328 330076 118380
rect 338488 118328 338540 118380
rect 396264 118328 396316 118380
rect 400864 118328 400916 118380
rect 474004 118328 474056 118380
rect 237196 118260 237248 118312
rect 255780 118260 255832 118312
rect 256608 118260 256660 118312
rect 265532 118260 265584 118312
rect 306012 118260 306064 118312
rect 332876 118260 332928 118312
rect 337844 118260 337896 118312
rect 351184 118260 351236 118312
rect 362316 118260 362368 118312
rect 443000 118260 443052 118312
rect 31668 118192 31720 118244
rect 107568 118192 107620 118244
rect 113088 118192 113140 118244
rect 175556 118192 175608 118244
rect 184848 118192 184900 118244
rect 229192 118192 229244 118244
rect 233148 118192 233200 118244
rect 253296 118192 253348 118244
rect 253848 118192 253900 118244
rect 263692 118192 263744 118244
rect 300492 118192 300544 118244
rect 28908 118124 28960 118176
rect 114468 118124 114520 118176
rect 129280 118124 129332 118176
rect 177396 118124 177448 118176
rect 179328 118124 179380 118176
rect 225788 118124 225840 118176
rect 234528 118124 234580 118176
rect 253940 118124 253992 118176
rect 257988 118124 258040 118176
rect 266360 118124 266412 118176
rect 267648 118124 267700 118176
rect 271052 118124 271104 118176
rect 291108 118124 291160 118176
rect 305184 118124 305236 118176
rect 307668 118192 307720 118244
rect 336924 118192 336976 118244
rect 339408 118192 339460 118244
rect 353944 118192 353996 118244
rect 356796 118192 356848 118244
rect 23388 118056 23440 118108
rect 110328 118056 110380 118108
rect 115204 118056 115256 118108
rect 126980 118056 127032 118108
rect 128176 118056 128228 118108
rect 133144 118056 133196 118108
rect 133236 118056 133288 118108
rect 173900 118056 173952 118108
rect 176568 118056 176620 118108
rect 223948 118056 224000 118108
rect 231768 118056 231820 118108
rect 252744 118056 252796 118108
rect 255228 118056 255280 118108
rect 264980 118056 265032 118108
rect 293132 118056 293184 118108
rect 307944 118056 307996 118108
rect 60648 117988 60700 118040
rect 82728 117988 82780 118040
rect 88340 117988 88392 118040
rect 179420 117988 179472 118040
rect 182088 117988 182140 118040
rect 226984 117988 227036 118040
rect 229008 117988 229060 118040
rect 251272 117988 251324 118040
rect 253756 117988 253808 118040
rect 264336 117988 264388 118040
rect 266268 117988 266320 118040
rect 270500 117988 270552 118040
rect 294972 117988 295024 118040
rect 9588 117920 9640 117972
rect 69848 117920 69900 117972
rect 122840 117920 122892 117972
rect 107568 117852 107620 117904
rect 149888 117852 149940 117904
rect 96528 117784 96580 117836
rect 99196 117784 99248 117836
rect 122104 117784 122156 117836
rect 122656 117784 122708 117836
rect 160836 117784 160888 117836
rect 71688 117716 71740 117768
rect 73804 117716 73856 117768
rect 79968 117716 80020 117768
rect 99472 117716 99524 117768
rect 80152 117648 80204 117700
rect 86960 117648 87012 117700
rect 122840 117716 122892 117768
rect 126888 117716 126940 117768
rect 162860 117716 162912 117768
rect 127624 117648 127676 117700
rect 128176 117648 128228 117700
rect 129096 117648 129148 117700
rect 129372 117648 129424 117700
rect 137284 117648 137336 117700
rect 130476 117580 130528 117632
rect 137652 117648 137704 117700
rect 166264 117648 166316 117700
rect 158996 117580 159048 117632
rect 177948 117920 178000 117972
rect 225144 117920 225196 117972
rect 226248 117920 226300 117972
rect 239404 117920 239456 117972
rect 197268 117852 197320 117904
rect 234988 117852 235040 117904
rect 238116 117852 238168 117904
rect 241704 117920 241756 117972
rect 251088 117920 251140 117972
rect 262496 117920 262548 117972
rect 264888 117920 264940 117972
rect 269856 117920 269908 117972
rect 279056 117920 279108 117972
rect 280344 117920 280396 117972
rect 280896 117920 280948 117972
rect 281448 117920 281500 117972
rect 241428 117852 241480 117904
rect 257620 117852 257672 117904
rect 263508 117852 263560 117904
rect 268660 117852 268712 117904
rect 296536 117852 296588 117904
rect 316684 118124 316736 118176
rect 339684 118124 339736 118176
rect 359280 118124 359332 118176
rect 360108 118124 360160 118176
rect 316592 118056 316644 118108
rect 343916 118056 343968 118108
rect 354956 118056 355008 118108
rect 364984 118056 365036 118108
rect 365996 118192 366048 118244
rect 449900 118192 449952 118244
rect 374644 118124 374696 118176
rect 456800 118124 456852 118176
rect 313188 117988 313240 118040
rect 347964 117988 348016 118040
rect 373356 118056 373408 118108
rect 463700 118056 463752 118108
rect 374644 117988 374696 118040
rect 377036 117988 377088 118040
rect 470600 117988 470652 118040
rect 321744 117920 321796 117972
rect 380716 117920 380768 117972
rect 477500 117920 477552 117972
rect 167736 117784 167788 117836
rect 189080 117784 189132 117836
rect 213828 117784 213880 117836
rect 243636 117784 243688 117836
rect 245752 117784 245804 117836
rect 260012 117784 260064 117836
rect 263416 117784 263468 117836
rect 269212 117784 269264 117836
rect 296168 117784 296220 117836
rect 191104 117716 191156 117768
rect 205180 117716 205232 117768
rect 217968 117716 218020 117768
rect 245660 117716 245712 117768
rect 246948 117716 247000 117768
rect 260840 117716 260892 117768
rect 262128 117716 262180 117768
rect 268016 117716 268068 117768
rect 277860 117716 277912 117768
rect 278688 117716 278740 117768
rect 169024 117648 169076 117700
rect 192668 117648 192720 117700
rect 213184 117648 213236 117700
rect 232504 117648 232556 117700
rect 233884 117648 233936 117700
rect 244280 117648 244332 117700
rect 245568 117648 245620 117700
rect 259460 117648 259512 117700
rect 311900 117852 311952 117904
rect 314568 117852 314620 117904
rect 322204 117852 322256 117904
rect 316408 117784 316460 117836
rect 331864 117852 331916 117904
rect 345848 117852 345900 117904
rect 407764 117852 407816 117904
rect 420828 117852 420880 117904
rect 489184 117852 489236 117904
rect 331128 117784 331180 117836
rect 337384 117784 337436 117836
rect 314660 117716 314712 117768
rect 315212 117716 315264 117768
rect 315948 117716 316000 117768
rect 320732 117716 320784 117768
rect 321376 117716 321428 117768
rect 321928 117716 321980 117768
rect 357992 117716 358044 117768
rect 171876 117580 171928 117632
rect 196624 117580 196676 117632
rect 211712 117580 211764 117632
rect 224224 117580 224276 117632
rect 236828 117580 236880 117632
rect 237288 117580 237340 117632
rect 240416 117580 240468 117632
rect 244188 117580 244240 117632
rect 258816 117580 258868 117632
rect 259276 117580 259328 117632
rect 263140 117580 263192 117632
rect 86960 117512 87012 117564
rect 96528 117512 96580 117564
rect 128820 117512 128872 117564
rect 137652 117512 137704 117564
rect 138664 117512 138716 117564
rect 139400 117512 139452 117564
rect 146760 117512 146812 117564
rect 235264 117512 235316 117564
rect 247776 117512 247828 117564
rect 248328 117512 248380 117564
rect 261300 117512 261352 117564
rect 67548 117444 67600 117496
rect 71044 117444 71096 117496
rect 168380 117444 168432 117496
rect 229744 117444 229796 117496
rect 238852 117444 238904 117496
rect 114468 117376 114520 117428
rect 148048 117376 148100 117428
rect 182180 117376 182232 117428
rect 186504 117376 186556 117428
rect 232504 117376 232556 117428
rect 92388 117308 92440 117360
rect 97908 117308 97960 117360
rect 109684 117308 109736 117360
rect 113088 117308 113140 117360
rect 133144 117308 133196 117360
rect 190460 117308 190512 117360
rect 190552 117308 190604 117360
rect 192116 117308 192168 117360
rect 225604 117308 225656 117360
rect 231308 117308 231360 117360
rect 232596 117308 232648 117360
rect 237288 117308 237340 117360
rect 240232 117444 240284 117496
rect 243544 117444 243596 117496
rect 249064 117444 249116 117496
rect 249708 117444 249760 117496
rect 262220 117444 262272 117496
rect 271788 117444 271840 117496
rect 273260 117444 273312 117496
rect 305368 117648 305420 117700
rect 312636 117648 312688 117700
rect 312728 117648 312780 117700
rect 319352 117648 319404 117700
rect 320088 117648 320140 117700
rect 308496 117580 308548 117632
rect 308956 117580 309008 117632
rect 311532 117580 311584 117632
rect 316592 117580 316644 117632
rect 360476 117648 360528 117700
rect 422852 117784 422904 117836
rect 486424 117784 486476 117836
rect 394700 117716 394752 117768
rect 394884 117716 394936 117768
rect 380256 117648 380308 117700
rect 393228 117648 393280 117700
rect 411904 117716 411956 117768
rect 480904 117716 480956 117768
rect 404360 117648 404412 117700
rect 415308 117648 415360 117700
rect 482284 117648 482336 117700
rect 331956 117580 332008 117632
rect 353116 117580 353168 117632
rect 425336 117580 425388 117632
rect 428464 117580 428516 117632
rect 496084 117580 496136 117632
rect 307208 117512 307260 117564
rect 309692 117512 309744 117564
rect 316684 117512 316736 117564
rect 419264 117512 419316 117564
rect 420184 117512 420236 117564
rect 430304 117512 430356 117564
rect 431224 117512 431276 117564
rect 242164 117376 242216 117428
rect 247224 117376 247276 117428
rect 269028 117376 269080 117428
rect 271880 117376 271932 117428
rect 272524 117376 272576 117428
rect 273536 117376 273588 117428
rect 284576 117376 284628 117428
rect 285496 117376 285548 117428
rect 303436 117376 303488 117428
rect 305644 117376 305696 117428
rect 239404 117308 239456 117360
rect 242256 117308 242308 117360
rect 242808 117308 242860 117360
rect 249892 117308 249944 117360
rect 250444 117308 250496 117360
rect 251456 117308 251508 117360
rect 252468 117308 252520 117360
rect 259276 117308 259328 117360
rect 259368 117308 259420 117360
rect 266820 117308 266872 117360
rect 271144 117308 271196 117360
rect 272340 117308 272392 117360
rect 273168 117308 273220 117360
rect 274180 117308 274232 117360
rect 279700 117308 279752 117360
rect 280068 117308 280120 117360
rect 282092 117308 282144 117360
rect 282828 117308 282880 117360
rect 283380 117308 283432 117360
rect 284024 117308 284076 117360
rect 285220 117308 285272 117360
rect 285588 117308 285640 117360
rect 286416 117308 286468 117360
rect 286968 117308 287020 117360
rect 287612 117308 287664 117360
rect 288348 117308 288400 117360
rect 288900 117308 288952 117360
rect 289544 117308 289596 117360
rect 290096 117308 290148 117360
rect 290740 117308 290792 117360
rect 291936 117308 291988 117360
rect 292396 117308 292448 117360
rect 294328 117308 294380 117360
rect 295248 117308 295300 117360
rect 295616 117308 295668 117360
rect 296628 117308 296680 117360
rect 297456 117308 297508 117360
rect 297916 117308 297968 117360
rect 299848 117308 299900 117360
rect 300768 117308 300820 117360
rect 301688 117308 301740 117360
rect 302884 117308 302936 117360
rect 302976 117308 303028 117360
rect 303528 117308 303580 117360
rect 306656 117308 306708 117360
rect 307668 117308 307720 117360
rect 314108 117444 314160 117496
rect 327448 117444 327500 117496
rect 334624 117444 334676 117496
rect 336648 117444 336700 117496
rect 341156 117444 341208 117496
rect 380256 117444 380308 117496
rect 383660 117444 383712 117496
rect 413744 117444 413796 117496
rect 414664 117444 414716 117496
rect 426348 117444 426400 117496
rect 429844 117444 429896 117496
rect 310888 117376 310940 117428
rect 315304 117376 315356 117428
rect 332968 117376 333020 117428
rect 333888 117376 333940 117428
rect 334808 117376 334860 117428
rect 338764 117376 338816 117428
rect 340328 117376 340380 117428
rect 342904 117376 342956 117428
rect 344008 117376 344060 117428
rect 345664 117376 345716 117428
rect 347596 117376 347648 117428
rect 349804 117376 349856 117428
rect 367836 117376 367888 117428
rect 369124 117376 369176 117428
rect 371516 117376 371568 117428
rect 377404 117376 377456 117428
rect 399668 117376 399720 117428
rect 400128 117376 400180 117428
rect 421748 117376 421800 117428
rect 422208 117376 422260 117428
rect 312544 117308 312596 117360
rect 313924 117308 313976 117360
rect 314568 117308 314620 117360
rect 318248 117308 318300 117360
rect 318708 117308 318760 117360
rect 319444 117308 319496 117360
rect 320088 117308 320140 117360
rect 322572 117308 322624 117360
rect 322848 117308 322900 117360
rect 323768 117308 323820 117360
rect 324228 117308 324280 117360
rect 324964 117308 325016 117360
rect 325516 117308 325568 117360
rect 326252 117308 326304 117360
rect 326988 117308 327040 117360
rect 328092 117308 328144 117360
rect 328368 117308 328420 117360
rect 329288 117308 329340 117360
rect 329748 117308 329800 117360
rect 330484 117308 330536 117360
rect 331128 117308 331180 117360
rect 331680 117308 331732 117360
rect 332508 117308 332560 117360
rect 333520 117308 333572 117360
rect 333796 117308 333848 117360
rect 337200 117308 337252 117360
rect 338028 117308 338080 117360
rect 341524 117308 341576 117360
rect 342168 117308 342220 117360
rect 342720 117308 342772 117360
rect 343548 117308 343600 117360
rect 344560 117308 344612 117360
rect 344928 117308 344980 117360
rect 347044 117308 347096 117360
rect 347688 117308 347740 117360
rect 348240 117308 348292 117360
rect 349068 117308 349120 117360
rect 350080 117308 350132 117360
rect 350448 117308 350500 117360
rect 351276 117308 351328 117360
rect 352472 117308 352524 117360
rect 352564 117308 352616 117360
rect 353208 117308 353260 117360
rect 353760 117308 353812 117360
rect 354588 117308 354640 117360
rect 355600 117308 355652 117360
rect 355968 117308 356020 117360
rect 358084 117308 358136 117360
rect 358636 117308 358688 117360
rect 361120 117308 361172 117360
rect 361488 117308 361540 117360
rect 363604 117308 363656 117360
rect 364248 117308 364300 117360
rect 364800 117308 364852 117360
rect 365628 117308 365680 117360
rect 366640 117308 366692 117360
rect 367008 117308 367060 117360
rect 369032 117308 369084 117360
rect 369768 117308 369820 117360
rect 370320 117308 370372 117360
rect 371148 117308 371200 117360
rect 372160 117308 372212 117360
rect 372528 117308 372580 117360
rect 374552 117308 374604 117360
rect 375196 117308 375248 117360
rect 375840 117308 375892 117360
rect 376668 117308 376720 117360
rect 377680 117308 377732 117360
rect 378048 117308 378100 117360
rect 378876 117308 378928 117360
rect 379428 117308 379480 117360
rect 380072 117308 380124 117360
rect 380808 117308 380860 117360
rect 381360 117308 381412 117360
rect 382188 117308 382240 117360
rect 382556 117308 382608 117360
rect 383568 117308 383620 117360
rect 384396 117308 384448 117360
rect 384856 117308 384908 117360
rect 385592 117308 385644 117360
rect 386328 117308 386380 117360
rect 386788 117308 386840 117360
rect 387616 117308 387668 117360
rect 388076 117308 388128 117360
rect 388904 117308 388956 117360
rect 389916 117308 389968 117360
rect 390376 117308 390428 117360
rect 391112 117308 391164 117360
rect 391848 117308 391900 117360
rect 392308 117308 392360 117360
rect 393136 117308 393188 117360
rect 393596 117308 393648 117360
rect 394424 117308 394476 117360
rect 395436 117308 395488 117360
rect 395896 117308 395948 117360
rect 396632 117308 396684 117360
rect 397368 117308 397420 117360
rect 397828 117308 397880 117360
rect 398656 117308 398708 117360
rect 399116 117308 399168 117360
rect 399944 117308 399996 117360
rect 402152 117308 402204 117360
rect 402796 117308 402848 117360
rect 403348 117308 403400 117360
rect 404268 117308 404320 117360
rect 405188 117308 405240 117360
rect 405648 117308 405700 117360
rect 406384 117308 406436 117360
rect 407028 117308 407080 117360
rect 407672 117308 407724 117360
rect 408408 117308 408460 117360
rect 408868 117308 408920 117360
rect 409696 117308 409748 117360
rect 410708 117308 410760 117360
rect 411168 117308 411220 117360
rect 413192 117308 413244 117360
rect 413928 117308 413980 117360
rect 414388 117308 414440 117360
rect 415308 117308 415360 117360
rect 416228 117308 416280 117360
rect 416688 117308 416740 117360
rect 418620 117308 418672 117360
rect 419448 117308 419500 117360
rect 419908 117308 419960 117360
rect 420828 117308 420880 117360
rect 422944 117308 422996 117360
rect 423588 117308 423640 117360
rect 424140 117308 424192 117360
rect 424968 117308 425020 117360
rect 425428 117308 425480 117360
rect 426348 117308 426400 117360
rect 427268 117308 427320 117360
rect 427728 117308 427780 117360
rect 429660 117308 429712 117360
rect 430488 117308 430540 117360
rect 430948 117308 431000 117360
rect 431868 117308 431920 117360
rect 432788 117308 432840 117360
rect 433248 117308 433300 117360
rect 433984 117308 434036 117360
rect 439504 117308 439556 117360
rect 133788 117240 133840 117292
rect 130292 117172 130344 117224
rect 133880 117172 133932 117224
rect 143448 117172 143500 117224
rect 154488 117172 154540 117224
rect 133880 117036 133932 117088
rect 143448 117036 143500 117088
rect 161388 117036 161440 117088
rect 171140 117172 171192 117224
rect 180708 117036 180760 117088
rect 182180 117172 182232 117224
rect 404360 117172 404412 117224
rect 410524 117172 410576 117224
rect 154488 116900 154540 116952
rect 161388 116900 161440 116952
rect 208492 116628 208544 116680
rect 209228 116628 209280 116680
rect 205640 116560 205692 116612
rect 206192 116560 206244 116612
rect 208400 116560 208452 116612
rect 208676 116560 208728 116612
rect 212540 116560 212592 116612
rect 212908 116560 212960 116612
rect 214012 116560 214064 116612
rect 214748 116560 214800 116612
rect 420276 115948 420328 116000
rect 420460 115948 420512 116000
rect 128728 115880 128780 115932
rect 129004 115880 129056 115932
rect 143632 115880 143684 115932
rect 143724 115880 143776 115932
rect 144920 115880 144972 115932
rect 145288 115880 145340 115932
rect 168472 115880 168524 115932
rect 168564 115880 168616 115932
rect 238944 115880 238996 115932
rect 239128 115880 239180 115932
rect 248236 115880 248288 115932
rect 248328 115880 248380 115932
rect 253756 115880 253808 115932
rect 253940 115880 253992 115932
rect 314016 115880 314068 115932
rect 314108 115880 314160 115932
rect 339684 115880 339736 115932
rect 339868 115880 339920 115932
rect 341248 115880 341300 115932
rect 341432 115880 341484 115932
rect 343916 115880 343968 115932
rect 344100 115880 344152 115932
rect 409328 114588 409380 114640
rect 409604 114588 409656 114640
rect 147956 114520 148008 114572
rect 148600 114520 148652 114572
rect 157432 114520 157484 114572
rect 157800 114520 157852 114572
rect 179604 114520 179656 114572
rect 179972 114520 180024 114572
rect 245384 114520 245436 114572
rect 245752 114520 245804 114572
rect 250076 114520 250128 114572
rect 250352 114520 250404 114572
rect 276112 114520 276164 114572
rect 276204 114520 276256 114572
rect 382924 114520 382976 114572
rect 383108 114520 383160 114572
rect 403716 114520 403768 114572
rect 403900 114520 403952 114572
rect 161664 114452 161716 114504
rect 161848 114452 161900 114504
rect 185032 114452 185084 114504
rect 185124 114452 185176 114504
rect 189080 114452 189132 114504
rect 189264 114452 189316 114504
rect 409420 114452 409472 114504
rect 409604 114452 409656 114504
rect 425980 114452 426032 114504
rect 431592 114452 431644 114504
rect 431684 114452 431736 114504
rect 147956 114384 148008 114436
rect 148232 114384 148284 114436
rect 426164 114384 426216 114436
rect 133880 113840 133932 113892
rect 134524 113840 134576 113892
rect 135260 113840 135312 113892
rect 135720 113840 135772 113892
rect 136732 113840 136784 113892
rect 137008 113840 137060 113892
rect 139492 113840 139544 113892
rect 140044 113840 140096 113892
rect 167000 113840 167052 113892
rect 167644 113840 167696 113892
rect 169852 113840 169904 113892
rect 170680 113840 170732 113892
rect 178040 113840 178092 113892
rect 178592 113840 178644 113892
rect 186320 113840 186372 113892
rect 187148 113840 187200 113892
rect 194600 113840 194652 113892
rect 195152 113840 195204 113892
rect 201500 113840 201552 113892
rect 201868 113840 201920 113892
rect 136640 113772 136692 113824
rect 137560 113772 137612 113824
rect 222200 113704 222252 113756
rect 222660 113704 222712 113756
rect 233424 113160 233476 113212
rect 233700 113160 233752 113212
rect 414756 113160 414808 113212
rect 415216 113160 415268 113212
rect 175372 111732 175424 111784
rect 176200 111732 176252 111784
rect 436928 111732 436980 111784
rect 579804 111732 579856 111784
rect 200120 111460 200172 111512
rect 200672 111460 200724 111512
rect 198740 110576 198792 110628
rect 199476 110576 199528 110628
rect 245752 109964 245804 110016
rect 246580 109964 246632 110016
rect 153292 109760 153344 109812
rect 154120 109760 154172 109812
rect 172520 109080 172572 109132
rect 173072 109080 173124 109132
rect 179604 109080 179656 109132
rect 159088 109012 159140 109064
rect 168564 109012 168616 109064
rect 190736 109080 190788 109132
rect 196072 109080 196124 109132
rect 383108 109080 383160 109132
rect 314108 109012 314160 109064
rect 388812 109012 388864 109064
rect 388996 109012 389048 109064
rect 394332 109012 394384 109064
rect 394516 109012 394568 109064
rect 403900 109012 403952 109064
rect 3240 108944 3292 108996
rect 131212 108944 131264 108996
rect 158996 108944 159048 108996
rect 168472 108944 168524 108996
rect 179604 108944 179656 108996
rect 190644 108944 190696 108996
rect 196072 108944 196124 108996
rect 314016 108944 314068 108996
rect 383108 108944 383160 108996
rect 403992 108944 404044 108996
rect 217048 106428 217100 106480
rect 317052 106360 317104 106412
rect 317236 106360 317288 106412
rect 143632 106292 143684 106344
rect 143724 106292 143776 106344
rect 216956 106292 217008 106344
rect 245384 106292 245436 106344
rect 245476 106292 245528 106344
rect 248236 106292 248288 106344
rect 248328 106292 248380 106344
rect 253756 106292 253808 106344
rect 253940 106292 253992 106344
rect 339684 106292 339736 106344
rect 339868 106292 339920 106344
rect 343916 106292 343968 106344
rect 344100 106292 344152 106344
rect 415216 106292 415268 106344
rect 431684 106292 431736 106344
rect 140780 106224 140832 106276
rect 140964 106224 141016 106276
rect 156144 106224 156196 106276
rect 156512 106224 156564 106276
rect 251272 106224 251324 106276
rect 251456 106224 251508 106276
rect 341432 106224 341484 106276
rect 341524 106224 341576 106276
rect 400588 106224 400640 106276
rect 400864 106224 400916 106276
rect 403992 106224 404044 106276
rect 404084 106224 404136 106276
rect 431592 106224 431644 106276
rect 415216 106156 415268 106208
rect 189080 104932 189132 104984
rect 189172 104932 189224 104984
rect 161664 104864 161716 104916
rect 161848 104864 161900 104916
rect 218244 104864 218296 104916
rect 218336 104864 218388 104916
rect 233332 104864 233384 104916
rect 233516 104864 233568 104916
rect 409328 104864 409380 104916
rect 409420 104864 409472 104916
rect 140964 104796 141016 104848
rect 141148 104796 141200 104848
rect 143632 104796 143684 104848
rect 143908 104796 143960 104848
rect 148048 104796 148100 104848
rect 148232 104796 148284 104848
rect 152096 104796 152148 104848
rect 152188 104796 152240 104848
rect 221280 104796 221332 104848
rect 221464 104796 221516 104848
rect 253572 104796 253624 104848
rect 253756 104796 253808 104848
rect 275928 104796 275980 104848
rect 276112 104796 276164 104848
rect 316868 104796 316920 104848
rect 317052 104796 317104 104848
rect 420552 104796 420604 104848
rect 420644 104796 420696 104848
rect 425980 104796 426032 104848
rect 426164 104796 426216 104848
rect 431408 104796 431460 104848
rect 431684 104796 431736 104848
rect 179604 103436 179656 103488
rect 179696 103436 179748 103488
rect 189172 103436 189224 103488
rect 189540 103436 189592 103488
rect 233332 103436 233384 103488
rect 233516 103436 233568 103488
rect 414940 103436 414992 103488
rect 415124 103436 415176 103488
rect 133144 99424 133196 99476
rect 138112 99424 138164 99476
rect 162952 99424 163004 99476
rect 216956 99424 217008 99476
rect 168380 99356 168432 99408
rect 168564 99356 168616 99408
rect 179604 99356 179656 99408
rect 227904 99424 227956 99476
rect 249892 99356 249944 99408
rect 313924 99356 313976 99408
rect 314108 99356 314160 99408
rect 133144 99288 133196 99340
rect 138112 99288 138164 99340
rect 162952 99288 163004 99340
rect 179696 99288 179748 99340
rect 216956 99288 217008 99340
rect 227812 99288 227864 99340
rect 383292 99424 383344 99476
rect 249984 99288 250036 99340
rect 383200 99288 383252 99340
rect 173808 98676 173860 98728
rect 173992 98676 174044 98728
rect 251272 96636 251324 96688
rect 251456 96636 251508 96688
rect 341524 96636 341576 96688
rect 400588 96636 400640 96688
rect 400772 96636 400824 96688
rect 168380 96568 168432 96620
rect 168564 96568 168616 96620
rect 180984 96568 181036 96620
rect 181168 96568 181220 96620
rect 186044 96568 186096 96620
rect 186228 96568 186280 96620
rect 203064 96568 203116 96620
rect 203248 96568 203300 96620
rect 204628 96568 204680 96620
rect 204812 96568 204864 96620
rect 209964 96568 210016 96620
rect 210148 96568 210200 96620
rect 274456 96568 274508 96620
rect 274732 96568 274784 96620
rect 341432 96568 341484 96620
rect 343916 96568 343968 96620
rect 344100 96568 344152 96620
rect 382924 96568 382976 96620
rect 383200 96568 383252 96620
rect 403716 96568 403768 96620
rect 403992 96568 404044 96620
rect 190644 96500 190696 96552
rect 190736 96500 190788 96552
rect 148048 95208 148100 95260
rect 148232 95208 148284 95260
rect 150716 95208 150768 95260
rect 150992 95208 151044 95260
rect 151820 95208 151872 95260
rect 152096 95208 152148 95260
rect 215576 95208 215628 95260
rect 215944 95208 215996 95260
rect 216956 95208 217008 95260
rect 217048 95208 217100 95260
rect 218336 95208 218388 95260
rect 218428 95208 218480 95260
rect 233516 95208 233568 95260
rect 253572 95208 253624 95260
rect 253756 95208 253808 95260
rect 275928 95208 275980 95260
rect 276020 95208 276072 95260
rect 316868 95208 316920 95260
rect 317052 95208 317104 95260
rect 341432 95208 341484 95260
rect 341524 95208 341576 95260
rect 409328 95208 409380 95260
rect 409604 95208 409656 95260
rect 420552 95208 420604 95260
rect 420736 95208 420788 95260
rect 185952 95140 186004 95192
rect 186044 95140 186096 95192
rect 431408 95140 431460 95192
rect 431500 95140 431552 95192
rect 189356 95072 189408 95124
rect 189540 95072 189592 95124
rect 233516 95072 233568 95124
rect 276020 95072 276072 95124
rect 276296 95072 276348 95124
rect 173808 93848 173860 93900
rect 173992 93848 174044 93900
rect 3424 93780 3476 93832
rect 14464 93780 14516 93832
rect 150532 91740 150584 91792
rect 150716 91740 150768 91792
rect 400772 91740 400824 91792
rect 401048 91740 401100 91792
rect 185032 89768 185084 89820
rect 227812 89700 227864 89752
rect 341340 89700 341392 89752
rect 341524 89700 341576 89752
rect 409512 89700 409564 89752
rect 180984 89632 181036 89684
rect 181168 89632 181220 89684
rect 184940 89632 184992 89684
rect 415124 89700 415176 89752
rect 251272 89632 251324 89684
rect 409604 89632 409656 89684
rect 227904 89564 227956 89616
rect 251364 89564 251416 89616
rect 415124 89564 415176 89616
rect 133512 88272 133564 88324
rect 580172 88272 580224 88324
rect 140872 86980 140924 87032
rect 140964 86980 141016 87032
rect 143632 86980 143684 87032
rect 143908 86980 143960 87032
rect 147864 86980 147916 87032
rect 148048 86980 148100 87032
rect 343916 86980 343968 87032
rect 344100 86980 344152 87032
rect 382924 86980 382976 87032
rect 383108 86980 383160 87032
rect 403716 86980 403768 87032
rect 403900 86980 403952 87032
rect 151820 86912 151872 86964
rect 151912 86912 151964 86964
rect 184756 86912 184808 86964
rect 184940 86912 184992 86964
rect 203248 86912 203300 86964
rect 203432 86912 203484 86964
rect 215484 86912 215536 86964
rect 215576 86912 215628 86964
rect 216956 86912 217008 86964
rect 217048 86912 217100 86964
rect 218244 86912 218296 86964
rect 218336 86912 218388 86964
rect 219716 86912 219768 86964
rect 219808 86912 219860 86964
rect 274640 86912 274692 86964
rect 274824 86912 274876 86964
rect 316960 86912 317012 86964
rect 317144 86912 317196 86964
rect 420552 86912 420604 86964
rect 420644 86912 420696 86964
rect 403900 86844 403952 86896
rect 403992 86844 404044 86896
rect 185952 85552 186004 85604
rect 186228 85552 186280 85604
rect 189264 85552 189316 85604
rect 189356 85552 189408 85604
rect 431500 85552 431552 85604
rect 431592 85552 431644 85604
rect 143632 85484 143684 85536
rect 143816 85484 143868 85536
rect 144828 85484 144880 85536
rect 145104 85484 145156 85536
rect 218244 85484 218296 85536
rect 218428 85484 218480 85536
rect 227536 85484 227588 85536
rect 227904 85484 227956 85536
rect 253572 85484 253624 85536
rect 253756 85484 253808 85536
rect 276112 85484 276164 85536
rect 276204 85484 276256 85536
rect 313924 85484 313976 85536
rect 314016 85484 314068 85536
rect 339132 85484 339184 85536
rect 339224 85484 339276 85536
rect 400772 85484 400824 85536
rect 400956 85484 401008 85536
rect 173808 84124 173860 84176
rect 173992 84124 174044 84176
rect 276020 84124 276072 84176
rect 276204 84124 276256 84176
rect 314016 84124 314068 84176
rect 314200 84124 314252 84176
rect 338948 84124 339000 84176
rect 339132 84124 339184 84176
rect 415032 84124 415084 84176
rect 415124 84124 415176 84176
rect 164516 82084 164568 82136
rect 164608 82016 164660 82068
rect 426072 80656 426124 80708
rect 426164 80656 426216 80708
rect 196164 80180 196216 80232
rect 240324 80112 240376 80164
rect 249892 80112 249944 80164
rect 196164 80044 196216 80096
rect 240232 80044 240284 80096
rect 249800 80044 249852 80096
rect 431592 80044 431644 80096
rect 431776 80044 431828 80096
rect 3148 79976 3200 80028
rect 436376 79976 436428 80028
rect 420552 77324 420604 77376
rect 420736 77324 420788 77376
rect 183652 77256 183704 77308
rect 183744 77256 183796 77308
rect 184756 77256 184808 77308
rect 185032 77256 185084 77308
rect 189080 77256 189132 77308
rect 189264 77256 189316 77308
rect 203064 77256 203116 77308
rect 203432 77256 203484 77308
rect 204352 77256 204404 77308
rect 204628 77256 204680 77308
rect 316960 77256 317012 77308
rect 317236 77256 317288 77308
rect 128912 77188 128964 77240
rect 129004 77188 129056 77240
rect 132316 77188 132368 77240
rect 580172 77188 580224 77240
rect 186228 75964 186280 76016
rect 186320 75964 186372 76016
rect 186412 75964 186464 76016
rect 186504 75964 186556 76016
rect 143632 75896 143684 75948
rect 143816 75896 143868 75948
rect 144828 75896 144880 75948
rect 145012 75896 145064 75948
rect 218244 75896 218296 75948
rect 218428 75896 218480 75948
rect 227536 75896 227588 75948
rect 227720 75896 227772 75948
rect 244280 75896 244332 75948
rect 244464 75896 244516 75948
rect 253572 75896 253624 75948
rect 253756 75896 253808 75948
rect 341708 75896 341760 75948
rect 341892 75896 341944 75948
rect 186228 75828 186280 75880
rect 186320 75828 186372 75880
rect 186412 75828 186464 75880
rect 186504 75828 186556 75880
rect 189080 75828 189132 75880
rect 189172 75828 189224 75880
rect 221004 75828 221056 75880
rect 221280 75828 221332 75880
rect 249800 75828 249852 75880
rect 249892 75828 249944 75880
rect 431592 75828 431644 75880
rect 431776 75828 431828 75880
rect 233240 74604 233292 74656
rect 233700 74604 233752 74656
rect 173808 74536 173860 74588
rect 173900 74536 173952 74588
rect 186228 74536 186280 74588
rect 186596 74536 186648 74588
rect 275928 74536 275980 74588
rect 276020 74536 276072 74588
rect 414940 74536 414992 74588
rect 415032 74536 415084 74588
rect 426072 74468 426124 74520
rect 426440 74468 426492 74520
rect 274732 72428 274784 72480
rect 275100 72428 275152 72480
rect 138112 71068 138164 71120
rect 138296 71068 138348 71120
rect 162952 71068 163004 71120
rect 163136 71068 163188 71120
rect 184756 71068 184808 71120
rect 185032 71068 185084 71120
rect 189172 70388 189224 70440
rect 249892 70388 249944 70440
rect 400956 70388 401008 70440
rect 203064 70320 203116 70372
rect 249984 70320 250036 70372
rect 401048 70320 401100 70372
rect 189172 70252 189224 70304
rect 203156 70252 203208 70304
rect 179604 67668 179656 67720
rect 181076 67668 181128 67720
rect 133144 67600 133196 67652
rect 133236 67600 133288 67652
rect 161572 67600 161624 67652
rect 161664 67600 161716 67652
rect 128820 67532 128872 67584
rect 129096 67532 129148 67584
rect 179696 67464 179748 67516
rect 209872 67600 209924 67652
rect 209964 67600 210016 67652
rect 274916 67600 274968 67652
rect 275100 67600 275152 67652
rect 341524 67600 341576 67652
rect 341892 67600 341944 67652
rect 383292 67600 383344 67652
rect 383660 67600 383712 67652
rect 400956 67600 401008 67652
rect 401048 67600 401100 67652
rect 409512 67600 409564 67652
rect 409604 67600 409656 67652
rect 420644 67600 420696 67652
rect 421012 67600 421064 67652
rect 203064 67532 203116 67584
rect 203156 67532 203208 67584
rect 238944 67532 238996 67584
rect 239128 67532 239180 67584
rect 181168 67464 181220 67516
rect 186228 66308 186280 66360
rect 186596 66308 186648 66360
rect 339224 66308 339276 66360
rect 339316 66308 339368 66360
rect 138112 66240 138164 66292
rect 138296 66240 138348 66292
rect 144828 66240 144880 66292
rect 145104 66240 145156 66292
rect 162952 66240 163004 66292
rect 163136 66240 163188 66292
rect 219624 66240 219676 66292
rect 219716 66240 219768 66292
rect 244372 66240 244424 66292
rect 244648 66240 244700 66292
rect 251272 66240 251324 66292
rect 251364 66240 251416 66292
rect 403808 66240 403860 66292
rect 404084 66240 404136 66292
rect 143632 66172 143684 66224
rect 143816 66172 143868 66224
rect 186136 66172 186188 66224
rect 186228 66172 186280 66224
rect 221004 66172 221056 66224
rect 221096 66172 221148 66224
rect 249892 66172 249944 66224
rect 409420 66172 409472 66224
rect 409512 66172 409564 66224
rect 414756 66172 414808 66224
rect 414940 66172 414992 66224
rect 250168 66104 250220 66156
rect 3332 64812 3384 64864
rect 131580 64812 131632 64864
rect 164516 64812 164568 64864
rect 164792 64812 164844 64864
rect 173808 64812 173860 64864
rect 173992 64812 174044 64864
rect 221004 64812 221056 64864
rect 221188 64812 221240 64864
rect 339132 64812 339184 64864
rect 339500 64812 339552 64864
rect 425980 64812 426032 64864
rect 426072 64812 426124 64864
rect 431408 64812 431460 64864
rect 431592 64812 431644 64864
rect 436836 64812 436888 64864
rect 579804 64812 579856 64864
rect 383292 60800 383344 60852
rect 420736 60732 420788 60784
rect 128820 60664 128872 60716
rect 129096 60664 129148 60716
rect 189172 60664 189224 60716
rect 189356 60664 189408 60716
rect 227812 60664 227864 60716
rect 227996 60664 228048 60716
rect 383200 60664 383252 60716
rect 420644 60664 420696 60716
rect 203064 57944 203116 57996
rect 203248 57944 203300 57996
rect 238944 57944 238996 57996
rect 239128 57944 239180 57996
rect 314016 57944 314068 57996
rect 132960 57876 133012 57928
rect 133236 57876 133288 57928
rect 181076 57876 181128 57928
rect 181168 57876 181220 57928
rect 209688 57876 209740 57928
rect 209964 57876 210016 57928
rect 227720 57876 227772 57928
rect 227996 57876 228048 57928
rect 233332 57876 233384 57928
rect 233516 57876 233568 57928
rect 276112 57876 276164 57928
rect 276204 57876 276256 57928
rect 383016 57876 383068 57928
rect 383200 57876 383252 57928
rect 420460 57876 420512 57928
rect 420736 57876 420788 57928
rect 314016 57808 314068 57860
rect 159088 56652 159140 56704
rect 219624 56652 219676 56704
rect 219808 56652 219860 56704
rect 143632 56584 143684 56636
rect 143816 56584 143868 56636
rect 145104 56584 145156 56636
rect 145196 56584 145248 56636
rect 159180 56584 159232 56636
rect 183744 56584 183796 56636
rect 183836 56584 183888 56636
rect 184756 56584 184808 56636
rect 184940 56584 184992 56636
rect 186136 56584 186188 56636
rect 186228 56584 186280 56636
rect 244280 56584 244332 56636
rect 244556 56584 244608 56636
rect 250076 56584 250128 56636
rect 250168 56584 250220 56636
rect 253664 56584 253716 56636
rect 253756 56584 253808 56636
rect 400772 56584 400824 56636
rect 400956 56584 401008 56636
rect 409328 56584 409380 56636
rect 409420 56584 409472 56636
rect 414756 56584 414808 56636
rect 415216 56584 415268 56636
rect 162952 56516 163004 56568
rect 163136 56516 163188 56568
rect 179512 56516 179564 56568
rect 179604 56516 179656 56568
rect 180984 56516 181036 56568
rect 181076 56516 181128 56568
rect 218152 56516 218204 56568
rect 218244 56516 218296 56568
rect 403808 56516 403860 56568
rect 403992 56516 404044 56568
rect 425980 55292 426032 55344
rect 426072 55292 426124 55344
rect 173808 55224 173860 55276
rect 174084 55224 174136 55276
rect 221004 55224 221056 55276
rect 221188 55224 221240 55276
rect 431408 55224 431460 55276
rect 431592 55224 431644 55276
rect 425796 55156 425848 55208
rect 426072 55156 426124 55208
rect 274732 53116 274784 53168
rect 275100 53116 275152 53168
rect 145196 51076 145248 51128
rect 189356 51076 189408 51128
rect 314016 51076 314068 51128
rect 145104 51008 145156 51060
rect 196072 51008 196124 51060
rect 189356 50940 189408 50992
rect 409328 51008 409380 51060
rect 409512 51008 409564 51060
rect 196164 50940 196216 50992
rect 314016 50940 314068 50992
rect 253664 48356 253716 48408
rect 253756 48356 253808 48408
rect 276112 48356 276164 48408
rect 276204 48356 276256 48408
rect 129096 48288 129148 48340
rect 159088 48288 159140 48340
rect 161572 48288 161624 48340
rect 161756 48288 161808 48340
rect 227720 48288 227772 48340
rect 227904 48288 227956 48340
rect 233332 48288 233384 48340
rect 233608 48288 233660 48340
rect 274916 48288 274968 48340
rect 275100 48288 275152 48340
rect 317144 48288 317196 48340
rect 317236 48288 317288 48340
rect 383016 48288 383068 48340
rect 383292 48288 383344 48340
rect 414940 48288 414992 48340
rect 415216 48288 415268 48340
rect 129004 48220 129056 48272
rect 159180 48220 159232 48272
rect 238760 48220 238812 48272
rect 238944 48220 238996 48272
rect 420552 48220 420604 48272
rect 420644 48220 420696 48272
rect 158996 46928 159048 46980
rect 159180 46928 159232 46980
rect 162952 46928 163004 46980
rect 163136 46928 163188 46980
rect 164608 46928 164660 46980
rect 164792 46928 164844 46980
rect 168472 46928 168524 46980
rect 168564 46928 168616 46980
rect 173900 46928 173952 46980
rect 174084 46928 174136 46980
rect 179512 46928 179564 46980
rect 179696 46928 179748 46980
rect 180984 46928 181036 46980
rect 181168 46928 181220 46980
rect 218152 46928 218204 46980
rect 218428 46928 218480 46980
rect 341248 46928 341300 46980
rect 341340 46928 341392 46980
rect 403808 46928 403860 46980
rect 404084 46928 404136 46980
rect 129096 46860 129148 46912
rect 253480 46860 253532 46912
rect 253756 46860 253808 46912
rect 276112 46860 276164 46912
rect 276204 46860 276256 46912
rect 341248 46792 341300 46844
rect 341432 46792 341484 46844
rect 129096 46724 129148 46776
rect 339224 45568 339276 45620
rect 339500 45568 339552 45620
rect 425796 45568 425848 45620
rect 425980 45568 426032 45620
rect 173716 45500 173768 45552
rect 173900 45500 173952 45552
rect 179420 45500 179472 45552
rect 179696 45500 179748 45552
rect 219716 45500 219768 45552
rect 219900 45500 219952 45552
rect 221004 45500 221056 45552
rect 221280 45500 221332 45552
rect 431500 45500 431552 45552
rect 431592 45500 431644 45552
rect 425796 45432 425848 45484
rect 425980 45432 426032 45484
rect 313740 43460 313792 43512
rect 314016 43460 314068 43512
rect 227904 41556 227956 41608
rect 132040 41352 132092 41404
rect 227904 41420 227956 41472
rect 580172 41352 580224 41404
rect 157340 38632 157392 38684
rect 157432 38632 157484 38684
rect 161572 38632 161624 38684
rect 161664 38632 161716 38684
rect 189080 38632 189132 38684
rect 189356 38632 189408 38684
rect 233240 38632 233292 38684
rect 233608 38632 233660 38684
rect 244280 38632 244332 38684
rect 244556 38632 244608 38684
rect 249800 38632 249852 38684
rect 250076 38632 250128 38684
rect 313740 38632 313792 38684
rect 313924 38632 313976 38684
rect 132960 38564 133012 38616
rect 133236 38564 133288 38616
rect 168380 38564 168432 38616
rect 168564 38564 168616 38616
rect 184940 38564 184992 38616
rect 185032 38564 185084 38616
rect 251180 38564 251232 38616
rect 251364 38564 251416 38616
rect 274732 38564 274784 38616
rect 275100 38564 275152 38616
rect 383016 38564 383068 38616
rect 383200 38564 383252 38616
rect 400588 38564 400640 38616
rect 400772 38564 400824 38616
rect 409328 38564 409380 38616
rect 409604 38564 409656 38616
rect 253480 37272 253532 37324
rect 253572 37272 253624 37324
rect 339224 37340 339276 37392
rect 158720 37204 158772 37256
rect 158996 37204 159048 37256
rect 244096 37204 244148 37256
rect 244280 37204 244332 37256
rect 249800 37204 249852 37256
rect 250168 37204 250220 37256
rect 339132 37204 339184 37256
rect 173716 35912 173768 35964
rect 173992 35912 174044 35964
rect 179420 35912 179472 35964
rect 179604 35912 179656 35964
rect 219716 35912 219768 35964
rect 219992 35912 220044 35964
rect 431408 35912 431460 35964
rect 431500 35912 431552 35964
rect 3424 35844 3476 35896
rect 436284 35844 436336 35896
rect 143816 34484 143868 34536
rect 144000 34484 144052 34536
rect 425980 34484 426032 34536
rect 426072 34484 426124 34536
rect 128820 33804 128872 33856
rect 129096 33804 129148 33856
rect 420460 33804 420512 33856
rect 420644 33804 420696 33856
rect 138112 31832 138164 31884
rect 138296 31832 138348 31884
rect 227904 31764 227956 31816
rect 251180 31764 251232 31816
rect 190644 31696 190696 31748
rect 190828 31696 190880 31748
rect 404084 31764 404136 31816
rect 415124 31764 415176 31816
rect 251272 31696 251324 31748
rect 415032 31696 415084 31748
rect 227904 31628 227956 31680
rect 404084 31628 404136 31680
rect 132132 30268 132184 30320
rect 580172 30268 580224 30320
rect 161664 29044 161716 29096
rect 161572 28976 161624 29028
rect 209596 28976 209648 29028
rect 209964 28976 210016 29028
rect 218244 28976 218296 29028
rect 218428 28976 218480 29028
rect 219992 29044 220044 29096
rect 253572 29044 253624 29096
rect 253756 29044 253808 29096
rect 276112 29044 276164 29096
rect 276204 29044 276256 29096
rect 227812 28976 227864 29028
rect 227904 28976 227956 29028
rect 274916 28976 274968 29028
rect 275100 28976 275152 29028
rect 317144 28976 317196 29028
rect 317236 28976 317288 29028
rect 383016 28976 383068 29028
rect 383292 28976 383344 29028
rect 400588 28976 400640 29028
rect 400864 28976 400916 29028
rect 409328 28976 409380 29028
rect 409420 28976 409472 29028
rect 415032 28976 415084 29028
rect 415216 28976 415268 29028
rect 150532 28908 150584 28960
rect 150624 28908 150676 28960
rect 151820 28908 151872 28960
rect 151912 28908 151964 28960
rect 156052 28908 156104 28960
rect 156144 28908 156196 28960
rect 157340 28908 157392 28960
rect 157432 28908 157484 28960
rect 168472 28908 168524 28960
rect 168656 28908 168708 28960
rect 173992 28908 174044 28960
rect 179604 28908 179656 28960
rect 179696 28908 179748 28960
rect 204352 28908 204404 28960
rect 204536 28908 204588 28960
rect 219808 28908 219860 28960
rect 420552 28908 420604 28960
rect 420644 28908 420696 28960
rect 233332 28840 233384 28892
rect 233516 28840 233568 28892
rect 313648 28840 313700 28892
rect 313924 28840 313976 28892
rect 173992 28772 174044 28824
rect 158720 27616 158772 27668
rect 158996 27616 159048 27668
rect 183376 27616 183428 27668
rect 183836 27616 183888 27668
rect 221096 27616 221148 27668
rect 221280 27616 221332 27668
rect 244096 27616 244148 27668
rect 244372 27616 244424 27668
rect 249892 27616 249944 27668
rect 250168 27616 250220 27668
rect 431408 27616 431460 27668
rect 431684 27616 431736 27668
rect 180708 27548 180760 27600
rect 181168 27548 181220 27600
rect 253572 27548 253624 27600
rect 253756 27548 253808 27600
rect 275928 27548 275980 27600
rect 276112 27548 276164 27600
rect 138112 26256 138164 26308
rect 138296 26256 138348 26308
rect 426072 24760 426124 24812
rect 426164 24760 426216 24812
rect 238944 24148 238996 24200
rect 239128 24148 239180 24200
rect 238024 22040 238076 22092
rect 244372 22040 244424 22092
rect 244556 22040 244608 22092
rect 249892 22040 249944 22092
rect 250076 22040 250128 22092
rect 341524 22040 341576 22092
rect 341708 22040 341760 22092
rect 238116 21972 238168 22024
rect 2780 21428 2832 21480
rect 4804 21428 4856 21480
rect 143724 19320 143776 19372
rect 143816 19320 143868 19372
rect 157340 19320 157392 19372
rect 157432 19320 157484 19372
rect 161572 19320 161624 19372
rect 161664 19320 161716 19372
rect 162952 19320 163004 19372
rect 204352 19320 204404 19372
rect 204444 19320 204496 19372
rect 209596 19320 209648 19372
rect 209780 19320 209832 19372
rect 238944 19320 238996 19372
rect 239128 19320 239180 19372
rect 313648 19320 313700 19372
rect 313924 19320 313976 19372
rect 409420 19320 409472 19372
rect 409604 19320 409656 19372
rect 128728 19252 128780 19304
rect 129096 19252 129148 19304
rect 140872 19252 140924 19304
rect 145012 19252 145064 19304
rect 145196 19252 145248 19304
rect 163044 19252 163096 19304
rect 168196 19252 168248 19304
rect 168380 19252 168432 19304
rect 173992 19252 174044 19304
rect 174176 19252 174228 19304
rect 183744 19252 183796 19304
rect 183928 19252 183980 19304
rect 400772 19252 400824 19304
rect 401048 19252 401100 19304
rect 140964 19184 141016 19236
rect 163044 17960 163096 18012
rect 163136 17960 163188 18012
rect 180708 17960 180760 18012
rect 181076 17960 181128 18012
rect 219716 17960 219768 18012
rect 219808 17960 219860 18012
rect 221004 17960 221056 18012
rect 221096 17960 221148 18012
rect 247960 17960 248012 18012
rect 248328 17960 248380 18012
rect 253480 17960 253532 18012
rect 253572 17960 253624 18012
rect 275928 17960 275980 18012
rect 276112 17960 276164 18012
rect 339316 17960 339368 18012
rect 339408 17960 339460 18012
rect 154856 17892 154908 17944
rect 161664 17892 161716 17944
rect 436744 17892 436796 17944
rect 579804 17892 579856 17944
rect 158720 17824 158772 17876
rect 158996 17824 159048 17876
rect 420460 14492 420512 14544
rect 420644 14492 420696 14544
rect 204444 12452 204496 12504
rect 276112 12452 276164 12504
rect 204352 12384 204404 12436
rect 314660 12384 314712 12436
rect 315764 12384 315816 12436
rect 276480 12316 276532 12368
rect 386236 12180 386288 12232
rect 488540 12180 488592 12232
rect 388904 12112 388956 12164
rect 492680 12112 492732 12164
rect 390376 12044 390428 12096
rect 495440 12044 495492 12096
rect 391756 11976 391808 12028
rect 499580 11976 499632 12028
rect 394424 11908 394476 11960
rect 502340 11908 502392 11960
rect 395896 11840 395948 11892
rect 506480 11840 506532 11892
rect 397276 11772 397328 11824
rect 510620 11772 510672 11824
rect 399944 11704 399996 11756
rect 513380 11704 513432 11756
rect 366916 10956 366968 11008
rect 451280 10956 451332 11008
rect 369768 10888 369820 10940
rect 455420 10888 455472 10940
rect 371056 10820 371108 10872
rect 459652 10820 459704 10872
rect 372436 10752 372488 10804
rect 462320 10752 462372 10804
rect 114468 10684 114520 10736
rect 190552 10684 190604 10736
rect 375196 10684 375248 10736
rect 466460 10684 466512 10736
rect 86868 10616 86920 10668
rect 178132 10616 178184 10668
rect 376576 10616 376628 10668
rect 469220 10616 469272 10668
rect 79968 10548 80020 10600
rect 174176 10548 174228 10600
rect 377956 10548 378008 10600
rect 473360 10548 473412 10600
rect 72976 10480 73028 10532
rect 169852 10480 169904 10532
rect 380808 10480 380860 10532
rect 477592 10480 477644 10532
rect 64788 10412 64840 10464
rect 167092 10412 167144 10464
rect 382096 10412 382148 10464
rect 480260 10412 480312 10464
rect 38568 10344 38620 10396
rect 146484 10344 146536 10396
rect 384856 10344 384908 10396
rect 485780 10344 485832 10396
rect 42708 10276 42760 10328
rect 154672 10276 154724 10328
rect 433156 10276 433208 10328
rect 581092 10276 581144 10328
rect 365536 10208 365588 10260
rect 448520 10208 448572 10260
rect 361396 10140 361448 10192
rect 441620 10140 441672 10192
rect 364248 10072 364300 10124
rect 444380 10072 444432 10124
rect 360016 10004 360068 10056
rect 437480 10004 437532 10056
rect 358636 9936 358688 9988
rect 434628 9936 434680 9988
rect 128728 9664 128780 9716
rect 128912 9664 128964 9716
rect 162860 9664 162912 9716
rect 163136 9664 163188 9716
rect 168196 9664 168248 9716
rect 168472 9664 168524 9716
rect 185860 9664 185912 9716
rect 186044 9664 186096 9716
rect 253480 9664 253532 9716
rect 253664 9664 253716 9716
rect 275008 9664 275060 9716
rect 275284 9664 275336 9716
rect 339132 9664 339184 9716
rect 339408 9664 339460 9716
rect 400772 9664 400824 9716
rect 400956 9664 401008 9716
rect 420460 9664 420512 9716
rect 420644 9664 420696 9716
rect 94504 9596 94556 9648
rect 182272 9596 182324 9648
rect 183652 9596 183704 9648
rect 183836 9596 183888 9648
rect 184296 9596 184348 9648
rect 185032 9596 185084 9648
rect 232872 9596 232924 9648
rect 238944 9596 238996 9648
rect 245384 9596 245436 9648
rect 246764 9596 246816 9648
rect 247960 9596 248012 9648
rect 368388 9596 368440 9648
rect 454868 9596 454920 9648
rect 45744 9528 45796 9580
rect 138664 9528 138716 9580
rect 143264 9528 143316 9580
rect 207112 9528 207164 9580
rect 245476 9528 245528 9580
rect 339132 9528 339184 9580
rect 343088 9528 343140 9580
rect 371148 9528 371200 9580
rect 458456 9528 458508 9580
rect 62396 9460 62448 9512
rect 165712 9460 165764 9512
rect 246764 9460 246816 9512
rect 247960 9460 248012 9512
rect 372528 9460 372580 9512
rect 462044 9460 462096 9512
rect 58808 9392 58860 9444
rect 164332 9392 164384 9444
rect 393136 9392 393188 9444
rect 501236 9392 501288 9444
rect 55220 9324 55272 9376
rect 154856 9324 154908 9376
rect 394516 9324 394568 9376
rect 504824 9324 504876 9376
rect 51632 9256 51684 9308
rect 160192 9256 160244 9308
rect 395988 9256 396040 9308
rect 508412 9256 508464 9308
rect 40960 9188 41012 9240
rect 154580 9188 154632 9240
rect 398656 9188 398708 9240
rect 512000 9188 512052 9240
rect 33876 9120 33928 9172
rect 150624 9120 150676 9172
rect 426164 9120 426216 9172
rect 566740 9120 566792 9172
rect 13636 9052 13688 9104
rect 133052 9052 133104 9104
rect 134892 9052 134944 9104
rect 202972 9052 203024 9104
rect 409512 9052 409564 9104
rect 409788 9052 409840 9104
rect 430488 9052 430540 9104
rect 573824 9052 573876 9104
rect 6460 8984 6512 9036
rect 136732 8984 136784 9036
rect 139676 8984 139728 9036
rect 205732 8984 205784 9036
rect 354496 8984 354548 9036
rect 427544 8984 427596 9036
rect 427636 8984 427688 9036
rect 570236 8984 570288 9036
rect 5264 8916 5316 8968
rect 136824 8916 136876 8968
rect 138480 8916 138532 8968
rect 204352 8916 204404 8968
rect 355876 8916 355928 8968
rect 431132 8916 431184 8968
rect 431684 8916 431736 8968
rect 577412 8916 577464 8968
rect 98092 8848 98144 8900
rect 183836 8848 183888 8900
rect 367008 8848 367060 8900
rect 451372 8848 451424 8900
rect 77852 8780 77904 8832
rect 84936 8712 84988 8764
rect 129004 8780 129056 8832
rect 200212 8780 200264 8832
rect 365628 8780 365680 8832
rect 447784 8780 447836 8832
rect 95700 8644 95752 8696
rect 129188 8712 129240 8764
rect 131396 8712 131448 8764
rect 201592 8712 201644 8764
rect 362868 8712 362920 8764
rect 444196 8712 444248 8764
rect 120632 8576 120684 8628
rect 129280 8644 129332 8696
rect 132592 8644 132644 8696
rect 201500 8644 201552 8696
rect 361488 8644 361540 8696
rect 440608 8644 440660 8696
rect 136088 8576 136140 8628
rect 203156 8576 203208 8628
rect 360108 8576 360160 8628
rect 437020 8576 437072 8628
rect 129372 8508 129424 8560
rect 126244 8440 126296 8492
rect 34980 8236 35032 8288
rect 115204 8236 115256 8288
rect 118240 8236 118292 8288
rect 194692 8236 194744 8288
rect 388996 8236 389048 8288
rect 494152 8236 494204 8288
rect 96896 8168 96948 8220
rect 183560 8168 183612 8220
rect 390468 8168 390520 8220
rect 497740 8168 497792 8220
rect 89720 8100 89772 8152
rect 179604 8100 179656 8152
rect 409604 8100 409656 8152
rect 534540 8100 534592 8152
rect 82636 8032 82688 8084
rect 175372 8032 175424 8084
rect 411076 8032 411128 8084
rect 538128 8032 538180 8084
rect 75460 7964 75512 8016
rect 172612 7964 172664 8016
rect 342168 7964 342220 8016
rect 402520 7964 402572 8016
rect 413928 7964 413980 8016
rect 541716 7964 541768 8016
rect 68284 7896 68336 7948
rect 168472 7896 168524 7948
rect 343456 7896 343508 7948
rect 406108 7896 406160 7948
rect 415124 7896 415176 7948
rect 545304 7896 545356 7948
rect 48136 7828 48188 7880
rect 158812 7828 158864 7880
rect 344836 7828 344888 7880
rect 409696 7828 409748 7880
rect 416596 7828 416648 7880
rect 548892 7828 548944 7880
rect 7656 7760 7708 7812
rect 136640 7760 136692 7812
rect 171784 7760 171836 7812
rect 222292 7760 222344 7812
rect 347688 7760 347740 7812
rect 413284 7760 413336 7812
rect 419448 7760 419500 7812
rect 552388 7760 552440 7812
rect 1676 7692 1728 7744
rect 133880 7692 133932 7744
rect 140872 7692 140924 7744
rect 205640 7692 205692 7744
rect 348976 7692 349028 7744
rect 416872 7692 416924 7744
rect 420644 7692 420696 7744
rect 555976 7692 556028 7744
rect 2872 7624 2924 7676
rect 135352 7624 135404 7676
rect 144460 7624 144512 7676
rect 208584 7624 208636 7676
rect 350356 7624 350408 7676
rect 420368 7624 420420 7676
rect 422116 7624 422168 7676
rect 559564 7624 559616 7676
rect 572 7556 624 7608
rect 133972 7556 134024 7608
rect 137284 7556 137336 7608
rect 204260 7556 204312 7608
rect 353208 7556 353260 7608
rect 423956 7556 424008 7608
rect 424968 7556 425020 7608
rect 563152 7556 563204 7608
rect 98000 7488 98052 7540
rect 99288 7488 99340 7540
rect 111156 7488 111208 7540
rect 190644 7488 190696 7540
rect 376392 7488 376444 7540
rect 376668 7488 376720 7540
rect 387616 7488 387668 7540
rect 490564 7488 490616 7540
rect 121828 7420 121880 7472
rect 195980 7420 196032 7472
rect 384948 7420 385000 7472
rect 486976 7420 487028 7472
rect 126612 7352 126664 7404
rect 198832 7352 198884 7404
rect 383384 7352 383436 7404
rect 483480 7352 483532 7404
rect 109960 7284 110012 7336
rect 127624 7284 127676 7336
rect 127808 7284 127860 7336
rect 198740 7284 198792 7336
rect 357348 7284 357400 7336
rect 433524 7284 433576 7336
rect 63592 7216 63644 7268
rect 128912 7216 128964 7268
rect 133788 7216 133840 7268
rect 202880 7216 202932 7268
rect 358728 7216 358780 7268
rect 435824 7216 435876 7268
rect 130200 7148 130252 7200
rect 200120 7148 200172 7200
rect 138020 6876 138072 6928
rect 138204 6876 138256 6928
rect 360200 6876 360252 6928
rect 101588 6808 101640 6860
rect 186412 6808 186464 6860
rect 321376 6808 321428 6860
rect 362132 6808 362184 6860
rect 376760 6876 376812 6928
rect 389088 6808 389140 6860
rect 495348 6808 495400 6860
rect 61200 6740 61252 6792
rect 164516 6740 164568 6792
rect 321468 6740 321520 6792
rect 363328 6740 363380 6792
rect 379612 6740 379664 6792
rect 387248 6740 387300 6792
rect 57612 6672 57664 6724
rect 162860 6672 162912 6724
rect 197176 6672 197228 6724
rect 212632 6672 212684 6724
rect 354496 6672 354548 6724
rect 360200 6672 360252 6724
rect 391756 6672 391808 6724
rect 498936 6740 498988 6792
rect 393228 6672 393280 6724
rect 502432 6672 502484 6724
rect 54024 6604 54076 6656
rect 161480 6604 161532 6656
rect 194600 6604 194652 6656
rect 214104 6604 214156 6656
rect 322756 6604 322808 6656
rect 366916 6604 366968 6656
rect 394608 6604 394660 6656
rect 506020 6604 506072 6656
rect 50528 6536 50580 6588
rect 158720 6536 158772 6588
rect 193312 6536 193364 6588
rect 215484 6536 215536 6588
rect 315948 6536 316000 6588
rect 351092 6536 351144 6588
rect 351184 6536 351236 6588
rect 395436 6536 395488 6588
rect 397368 6536 397420 6588
rect 509608 6536 509660 6588
rect 46940 6468 46992 6520
rect 157340 6468 157392 6520
rect 188620 6468 188672 6520
rect 218244 6468 218296 6520
rect 325516 6468 325568 6520
rect 370412 6468 370464 6520
rect 387248 6468 387300 6520
rect 391848 6468 391900 6520
rect 398748 6468 398800 6520
rect 513196 6468 513248 6520
rect 44548 6400 44600 6452
rect 156144 6400 156196 6452
rect 188068 6400 188120 6452
rect 219716 6400 219768 6452
rect 326896 6400 326948 6452
rect 374000 6400 374052 6452
rect 400036 6400 400088 6452
rect 516784 6400 516836 6452
rect 39764 6332 39816 6384
rect 153292 6332 153344 6384
rect 157524 6332 157576 6384
rect 214012 6332 214064 6384
rect 328276 6332 328328 6384
rect 377588 6332 377640 6384
rect 402796 6332 402848 6384
rect 520280 6332 520332 6384
rect 18328 6264 18380 6316
rect 135444 6264 135496 6316
rect 161112 6264 161164 6316
rect 216772 6264 216824 6316
rect 331128 6264 331180 6316
rect 381176 6264 381228 6316
rect 404176 6264 404228 6316
rect 523868 6264 523920 6316
rect 32680 6196 32732 6248
rect 84200 6196 84252 6248
rect 103428 6196 103480 6248
rect 113180 6196 113232 6248
rect 122748 6196 122800 6248
rect 128360 6196 128412 6248
rect 153936 6196 153988 6248
rect 212540 6196 212592 6248
rect 332416 6196 332468 6248
rect 384672 6196 384724 6248
rect 408408 6196 408460 6248
rect 531044 6196 531096 6248
rect 4068 6128 4120 6180
rect 135260 6128 135312 6180
rect 135352 6128 135404 6180
rect 150348 6128 150400 6180
rect 150440 6128 150492 6180
rect 211252 6128 211304 6180
rect 333704 6128 333756 6180
rect 388260 6128 388312 6180
rect 405556 6128 405608 6180
rect 527456 6128 527508 6180
rect 102784 6060 102836 6112
rect 186504 6060 186556 6112
rect 318616 6060 318668 6112
rect 358544 6060 358596 6112
rect 387708 6060 387760 6112
rect 491760 6060 491812 6112
rect 84200 5992 84252 6044
rect 103428 5992 103480 6044
rect 105176 5992 105228 6044
rect 187700 5992 187752 6044
rect 317328 5992 317380 6044
rect 356152 5992 356204 6044
rect 383476 5992 383528 6044
rect 484584 5992 484636 6044
rect 106372 5924 106424 5976
rect 187792 5924 187844 5976
rect 320088 5924 320140 5976
rect 359740 5924 359792 5976
rect 386328 5924 386380 5976
rect 488172 5924 488224 5976
rect 108764 5856 108816 5908
rect 189356 5856 189408 5908
rect 317052 5856 317104 5908
rect 354956 5856 355008 5908
rect 379336 5856 379388 5908
rect 476304 5856 476356 5908
rect 81440 5788 81492 5840
rect 109684 5788 109736 5840
rect 112352 5788 112404 5840
rect 191932 5788 191984 5840
rect 315856 5788 315908 5840
rect 352564 5788 352616 5840
rect 382188 5788 382240 5840
rect 479892 5788 479944 5840
rect 116032 5720 116084 5772
rect 193220 5720 193272 5772
rect 348424 5720 348476 5772
rect 354496 5720 354548 5772
rect 378048 5720 378100 5772
rect 472716 5720 472768 5772
rect 119436 5652 119488 5704
rect 194692 5652 194744 5704
rect 373908 5652 373960 5704
rect 465632 5652 465684 5704
rect 113180 5584 113232 5636
rect 122748 5584 122800 5636
rect 123024 5584 123076 5636
rect 197544 5584 197596 5636
rect 376392 5584 376444 5636
rect 469128 5584 469180 5636
rect 128360 5516 128412 5568
rect 135352 5516 135404 5568
rect 353944 5516 353996 5568
rect 399024 5516 399076 5568
rect 80244 5448 80296 5500
rect 175464 5448 175516 5500
rect 209228 5448 209280 5500
rect 232872 5448 232924 5500
rect 335268 5448 335320 5500
rect 390652 5448 390704 5500
rect 415308 5448 415360 5500
rect 544108 5448 544160 5500
rect 76656 5380 76708 5432
rect 172520 5380 172572 5432
rect 208308 5380 208360 5432
rect 237472 5380 237524 5432
rect 343088 5380 343140 5432
rect 397828 5380 397880 5432
rect 416688 5380 416740 5432
rect 547696 5380 547748 5432
rect 73068 5312 73120 5364
rect 171232 5312 171284 5364
rect 173900 5312 173952 5364
rect 213920 5312 213972 5364
rect 340788 5312 340840 5364
rect 401324 5312 401376 5364
rect 418068 5312 418120 5364
rect 551192 5312 551244 5364
rect 69480 5244 69532 5296
rect 169944 5244 169996 5296
rect 174176 5244 174228 5296
rect 223672 5244 223724 5296
rect 343548 5244 343600 5296
rect 404912 5244 404964 5296
rect 420828 5244 420880 5296
rect 554780 5244 554832 5296
rect 65984 5176 66036 5228
rect 167000 5176 167052 5228
rect 170588 5176 170640 5228
rect 221004 5176 221056 5228
rect 303528 5176 303580 5228
rect 327632 5176 327684 5228
rect 344928 5176 344980 5228
rect 408500 5176 408552 5228
rect 422208 5176 422260 5228
rect 558368 5176 558420 5228
rect 37372 5108 37424 5160
rect 153384 5108 153436 5160
rect 160008 5108 160060 5160
rect 209872 5108 209924 5160
rect 307668 5108 307720 5160
rect 334716 5108 334768 5160
rect 346308 5108 346360 5160
rect 412088 5108 412140 5160
rect 426348 5108 426400 5160
rect 565544 5108 565596 5160
rect 30288 5040 30340 5092
rect 149060 5040 149112 5092
rect 167092 5040 167144 5092
rect 219532 5040 219584 5092
rect 304908 5040 304960 5092
rect 331220 5040 331272 5092
rect 349068 5040 349120 5092
rect 415676 5040 415728 5092
rect 423496 5040 423548 5092
rect 561956 5040 562008 5092
rect 26700 4972 26752 5024
rect 147772 4972 147824 5024
rect 163504 4972 163556 5024
rect 218060 4972 218112 5024
rect 219348 4972 219400 5024
rect 245752 4972 245804 5024
rect 308956 4972 309008 5024
rect 338304 4972 338356 5024
rect 350448 4972 350500 5024
rect 419172 4972 419224 5024
rect 427728 4972 427780 5024
rect 569040 4972 569092 5024
rect 21916 4904 21968 4956
rect 145012 4904 145064 4956
rect 158720 4904 158772 4956
rect 215300 4904 215352 4956
rect 215852 4904 215904 4956
rect 244556 4904 244608 4956
rect 310428 4904 310480 4956
rect 341892 4904 341944 4956
rect 351828 4904 351880 4956
rect 422760 4904 422812 4956
rect 429108 4904 429160 4956
rect 572628 4904 572680 4956
rect 17224 4836 17276 4888
rect 142252 4836 142304 4888
rect 145656 4836 145708 4888
rect 208400 4836 208452 4888
rect 208676 4836 208728 4888
rect 240140 4836 240192 4888
rect 311808 4836 311860 4888
rect 345480 4836 345532 4888
rect 354588 4836 354640 4888
rect 426348 4836 426400 4888
rect 431868 4836 431920 4888
rect 576216 4836 576268 4888
rect 12440 4768 12492 4820
rect 139492 4768 139544 4820
rect 142068 4768 142120 4820
rect 207020 4768 207072 4820
rect 212264 4768 212316 4820
rect 242992 4768 243044 4820
rect 314568 4768 314620 4820
rect 349068 4768 349120 4820
rect 355968 4768 356020 4820
rect 429936 4768 429988 4820
rect 433248 4768 433300 4820
rect 579804 4768 579856 4820
rect 83832 4700 83884 4752
rect 176752 4700 176804 4752
rect 206928 4700 206980 4752
rect 234712 4700 234764 4752
rect 338028 4700 338080 4752
rect 394240 4700 394292 4752
rect 412548 4700 412600 4752
rect 540520 4700 540572 4752
rect 90916 4632 90968 4684
rect 180892 4632 180944 4684
rect 204352 4632 204404 4684
rect 233516 4632 233568 4684
rect 333796 4632 333848 4684
rect 387064 4632 387116 4684
rect 411168 4632 411220 4684
rect 536932 4632 536984 4684
rect 87328 4564 87380 4616
rect 178040 4564 178092 4616
rect 204260 4564 204312 4616
rect 231952 4564 232004 4616
rect 329656 4564 329708 4616
rect 379980 4564 380032 4616
rect 409788 4564 409840 4616
rect 533436 4564 533488 4616
rect 49332 4496 49384 4548
rect 130476 4496 130528 4548
rect 162124 4496 162176 4548
rect 208492 4496 208544 4548
rect 332508 4496 332560 4548
rect 383568 4496 383620 4548
rect 406936 4496 406988 4548
rect 529848 4496 529900 4548
rect 52828 4428 52880 4480
rect 122104 4428 122156 4480
rect 202972 4428 203024 4480
rect 229192 4428 229244 4480
rect 328368 4428 328420 4480
rect 376392 4428 376444 4480
rect 405648 4428 405700 4480
rect 526260 4428 526312 4480
rect 70676 4360 70728 4412
rect 120724 4360 120776 4412
rect 120816 4360 120868 4412
rect 146392 4360 146444 4412
rect 202880 4360 202932 4412
rect 227996 4360 228048 4412
rect 326988 4360 327040 4412
rect 372804 4360 372856 4412
rect 404268 4360 404320 4412
rect 522672 4360 522724 4412
rect 324136 4292 324188 4344
rect 369216 4292 369268 4344
rect 401508 4292 401560 4344
rect 519084 4292 519136 4344
rect 322848 4224 322900 4276
rect 365720 4224 365772 4276
rect 400128 4224 400180 4276
rect 515588 4224 515640 4276
rect 25504 4088 25556 4140
rect 120816 4088 120868 4140
rect 125416 4088 125468 4140
rect 170404 4088 170456 4140
rect 175372 4088 175424 4140
rect 176568 4088 176620 4140
rect 181352 4088 181404 4140
rect 182088 4088 182140 4140
rect 182548 4088 182600 4140
rect 183468 4088 183520 4140
rect 188436 4088 188488 4140
rect 188988 4088 189040 4140
rect 196808 4088 196860 4140
rect 197268 4088 197320 4140
rect 199200 4088 199252 4140
rect 200028 4088 200080 4140
rect 203892 4088 203944 4140
rect 229744 4088 229796 4140
rect 231308 4088 231360 4140
rect 231768 4088 231820 4140
rect 232504 4088 232556 4140
rect 233148 4088 233200 4140
rect 233700 4088 233752 4140
rect 234528 4088 234580 4140
rect 234804 4088 234856 4140
rect 235908 4088 235960 4140
rect 236000 4088 236052 4140
rect 237288 4088 237340 4140
rect 239588 4088 239640 4140
rect 240048 4088 240100 4140
rect 240784 4088 240836 4140
rect 241428 4088 241480 4140
rect 243176 4088 243228 4140
rect 244188 4088 244240 4140
rect 244372 4088 244424 4140
rect 245568 4088 245620 4140
rect 249156 4088 249208 4140
rect 249708 4088 249760 4140
rect 251456 4088 251508 4140
rect 252468 4088 252520 4140
rect 252652 4088 252704 4140
rect 253848 4088 253900 4140
rect 274088 4088 274140 4140
rect 274548 4088 274600 4140
rect 277308 4088 277360 4140
rect 277676 4088 277728 4140
rect 278596 4088 278648 4140
rect 280068 4088 280120 4140
rect 284116 4088 284168 4140
rect 289544 4088 289596 4140
rect 289728 4088 289780 4140
rect 301412 4088 301464 4140
rect 312544 4088 312596 4140
rect 314568 4088 314620 4140
rect 324228 4088 324280 4140
rect 368020 4088 368072 4140
rect 379428 4088 379480 4140
rect 475108 4088 475160 4140
rect 477500 4088 477552 4140
rect 478696 4088 478748 4140
rect 480904 4088 480956 4140
rect 481272 4088 481324 4140
rect 489184 4088 489236 4140
rect 489552 4088 489604 4140
rect 496084 4088 496136 4140
rect 503536 4088 503588 4140
rect 503812 4088 503864 4140
rect 571432 4088 571484 4140
rect 42156 4020 42208 4072
rect 42708 4020 42760 4072
rect 43352 4020 43404 4072
rect 155960 4020 156012 4072
rect 164700 4020 164752 4072
rect 188620 4020 188672 4072
rect 189632 4020 189684 4072
rect 225604 4020 225656 4072
rect 253664 4020 253716 4072
rect 279976 4020 280028 4072
rect 282460 4020 282512 4072
rect 291108 4020 291160 4072
rect 303804 4020 303856 4072
rect 325608 4020 325660 4072
rect 371608 4020 371660 4072
rect 383476 4020 383528 4072
rect 482284 4020 482336 4072
rect 500224 4020 500276 4072
rect 578608 4020 578660 4072
rect 36176 3952 36228 4004
rect 151912 3952 151964 4004
rect 156328 3952 156380 4004
rect 194600 3952 194652 4004
rect 209872 3952 209924 4004
rect 238116 3952 238168 4004
rect 253848 3952 253900 4004
rect 286968 3952 287020 4004
rect 295524 3952 295576 4004
rect 297916 3952 297968 4004
rect 316960 3952 317012 4004
rect 329748 3952 329800 4004
rect 378784 3952 378836 4004
rect 29092 3884 29144 3936
rect 147956 3884 148008 3936
rect 152740 3884 152792 3936
rect 197176 3884 197228 3936
rect 202696 3884 202748 3936
rect 231124 3884 231176 3936
rect 293868 3884 293920 3936
rect 309784 3884 309836 3936
rect 312636 3884 312688 3936
rect 332416 3884 332468 3936
rect 338764 3884 338816 3936
rect 389456 3884 389508 3936
rect 402888 3884 402940 3936
rect 521476 3952 521528 4004
rect 407028 3884 407080 3936
rect 528652 3884 528704 3936
rect 24308 3816 24360 3868
rect 146300 3816 146352 3868
rect 151544 3816 151596 3868
rect 196624 3816 196676 3868
rect 198004 3816 198056 3868
rect 206928 3816 206980 3868
rect 211068 3816 211120 3868
rect 239404 3816 239456 3868
rect 285588 3816 285640 3868
rect 293132 3816 293184 3868
rect 295248 3816 295300 3868
rect 310980 3816 311032 3868
rect 313924 3816 313976 3868
rect 335912 3816 335964 3868
rect 341708 3816 341760 3868
rect 393044 3816 393096 3868
rect 409512 3816 409564 3868
rect 535736 3816 535788 3868
rect 20720 3748 20772 3800
rect 143724 3748 143776 3800
rect 172980 3748 173032 3800
rect 180064 3748 180116 3800
rect 180156 3748 180208 3800
rect 222108 3748 222160 3800
rect 222844 3748 222896 3800
rect 226432 3748 226484 3800
rect 228916 3748 228968 3800
rect 19524 3680 19576 3732
rect 143540 3680 143592 3732
rect 155132 3680 155184 3732
rect 173900 3680 173952 3732
rect 176752 3680 176804 3732
rect 223764 3680 223816 3732
rect 226524 3680 226576 3732
rect 14832 3612 14884 3664
rect 140964 3612 141016 3664
rect 186228 3612 186280 3664
rect 222200 3612 222252 3664
rect 227720 3612 227772 3664
rect 229008 3612 229060 3664
rect 16028 3544 16080 3596
rect 142344 3544 142396 3596
rect 169392 3544 169444 3596
rect 220820 3544 220872 3596
rect 288256 3748 288308 3800
rect 299112 3748 299164 3800
rect 302884 3748 302936 3800
rect 230112 3680 230164 3732
rect 251180 3680 251232 3732
rect 291016 3680 291068 3732
rect 302608 3680 302660 3732
rect 250444 3612 250496 3664
rect 284208 3612 284260 3664
rect 290740 3612 290792 3664
rect 292396 3612 292448 3664
rect 306196 3680 306248 3732
rect 309600 3748 309652 3800
rect 321652 3748 321704 3800
rect 333888 3748 333940 3800
rect 385868 3748 385920 3800
rect 414664 3748 414716 3800
rect 542912 3748 542964 3800
rect 325240 3680 325292 3732
rect 342904 3680 342956 3732
rect 400220 3680 400272 3732
rect 420184 3680 420236 3732
rect 553584 3680 553636 3732
rect 305644 3612 305696 3664
rect 328828 3612 328880 3664
rect 345664 3612 345716 3664
rect 407304 3612 407356 3664
rect 407764 3612 407816 3664
rect 410892 3612 410944 3664
rect 423588 3612 423640 3664
rect 560760 3612 560812 3664
rect 250076 3544 250128 3596
rect 279792 3544 279844 3596
rect 283656 3544 283708 3596
rect 286876 3544 286928 3596
rect 296720 3544 296772 3596
rect 298008 3544 298060 3596
rect 318064 3544 318116 3596
rect 318708 3544 318760 3596
rect 357348 3544 357400 3596
rect 358084 3544 358136 3596
rect 364524 3544 364576 3596
rect 364984 3544 365036 3596
rect 428740 3544 428792 3596
rect 429844 3544 429896 3596
rect 567844 3544 567896 3596
rect 8852 3476 8904 3528
rect 9588 3476 9640 3528
rect 10048 3476 10100 3528
rect 138020 3476 138072 3528
rect 146852 3476 146904 3528
rect 162124 3476 162176 3528
rect 165896 3476 165948 3528
rect 219440 3476 219492 3528
rect 222108 3476 222160 3528
rect 222844 3476 222896 3528
rect 222936 3476 222988 3528
rect 248512 3476 248564 3528
rect 257436 3476 257488 3528
rect 257988 3476 258040 3528
rect 259828 3476 259880 3528
rect 260748 3476 260800 3528
rect 262220 3476 262272 3528
rect 263508 3476 263560 3528
rect 265808 3476 265860 3528
rect 266268 3476 266320 3528
rect 268108 3476 268160 3528
rect 269028 3476 269080 3528
rect 271696 3476 271748 3528
rect 272524 3476 272576 3528
rect 281448 3476 281500 3528
rect 284760 3476 284812 3528
rect 285404 3476 285456 3528
rect 294328 3476 294380 3528
rect 296628 3476 296680 3528
rect 11244 3408 11296 3460
rect 139584 3408 139636 3460
rect 149244 3408 149296 3460
rect 160008 3408 160060 3460
rect 162308 3408 162360 3460
rect 216956 3408 217008 3460
rect 218152 3408 218204 3460
rect 245844 3408 245896 3460
rect 267004 3408 267056 3460
rect 267648 3408 267700 3460
rect 270500 3408 270552 3460
rect 271788 3408 271840 3460
rect 285496 3408 285548 3460
rect 291936 3408 291988 3460
rect 292488 3408 292540 3460
rect 307392 3408 307444 3460
rect 315304 3476 315356 3528
rect 343088 3476 343140 3528
rect 349804 3476 349856 3528
rect 414480 3476 414532 3528
rect 439504 3476 439556 3528
rect 582196 3476 582248 3528
rect 313372 3408 313424 3460
rect 27896 3340 27948 3392
rect 28908 3340 28960 3392
rect 60004 3340 60056 3392
rect 60648 3340 60700 3392
rect 71872 3340 71924 3392
rect 72976 3340 73028 3392
rect 73804 3340 73856 3392
rect 74264 3340 74316 3392
rect 86132 3340 86184 3392
rect 86868 3340 86920 3392
rect 93308 3340 93360 3392
rect 174268 3340 174320 3392
rect 183744 3340 183796 3392
rect 202880 3340 202932 3392
rect 206284 3340 206336 3392
rect 232320 3340 232372 3392
rect 250352 3340 250404 3392
rect 251088 3340 251140 3392
rect 282828 3340 282880 3392
rect 287152 3340 287204 3392
rect 289636 3340 289688 3392
rect 300308 3340 300360 3392
rect 300768 3340 300820 3392
rect 309600 3340 309652 3392
rect 100484 3272 100536 3324
rect 184296 3272 184348 3324
rect 193220 3272 193272 3324
rect 194508 3272 194560 3324
rect 194600 3272 194652 3324
rect 202972 3272 203024 3324
rect 207480 3272 207532 3324
rect 225236 3272 225288 3324
rect 225328 3272 225380 3324
rect 226248 3272 226300 3324
rect 282736 3272 282788 3324
rect 103980 3204 104032 3256
rect 186320 3204 186372 3256
rect 200396 3204 200448 3256
rect 224224 3204 224276 3256
rect 261024 3204 261076 3256
rect 262128 3204 262180 3256
rect 113548 3136 113600 3188
rect 114468 3136 114520 3188
rect 115940 3136 115992 3188
rect 117136 3136 117188 3188
rect 107568 3068 107620 3120
rect 167644 3136 167696 3188
rect 180064 3136 180116 3188
rect 186136 3136 186188 3188
rect 192024 3136 192076 3188
rect 213184 3136 213236 3188
rect 220544 3136 220596 3188
rect 79048 3000 79100 3052
rect 79968 3000 80020 3052
rect 114744 3000 114796 3052
rect 169024 3068 169076 3120
rect 190828 3068 190880 3120
rect 204260 3068 204312 3120
rect 214656 3068 214708 3120
rect 233884 3068 233936 3120
rect 241980 3136 242032 3188
rect 242808 3136 242860 3188
rect 281356 3136 281408 3188
rect 285956 3136 286008 3188
rect 288348 3272 288400 3324
rect 297916 3272 297968 3324
rect 309048 3204 309100 3256
rect 339500 3408 339552 3460
rect 352472 3408 352524 3460
rect 421564 3408 421616 3460
rect 431224 3408 431276 3460
rect 575020 3408 575072 3460
rect 334624 3340 334676 3392
rect 375196 3340 375248 3392
rect 375288 3340 375340 3392
rect 467932 3340 467984 3392
rect 493324 3340 493376 3392
rect 564348 3340 564400 3392
rect 331956 3272 332008 3324
rect 360936 3272 360988 3324
rect 369124 3272 369176 3324
rect 453672 3272 453724 3324
rect 489552 3272 489604 3324
rect 557172 3272 557224 3324
rect 319444 3204 319496 3256
rect 346676 3204 346728 3256
rect 377404 3204 377456 3256
rect 460848 3204 460900 3256
rect 482192 3204 482244 3256
rect 546500 3204 546552 3256
rect 288348 3136 288400 3188
rect 322204 3136 322256 3188
rect 350264 3136 350316 3188
rect 380164 3136 380216 3188
rect 446588 3136 446640 3188
rect 451280 3136 451332 3188
rect 452476 3136 452528 3188
rect 486424 3136 486476 3188
rect 550088 3136 550140 3188
rect 242164 3068 242216 3120
rect 258632 3068 258684 3120
rect 259368 3068 259420 3120
rect 331864 3068 331916 3120
rect 353760 3068 353812 3120
rect 374644 3068 374696 3120
rect 432328 3068 432380 3120
rect 481272 3068 481324 3120
rect 539324 3068 539376 3120
rect 124220 3000 124272 3052
rect 125508 3000 125560 3052
rect 148048 3000 148100 3052
rect 191104 3000 191156 3052
rect 194416 3000 194468 3052
rect 204352 3000 204404 3052
rect 217048 3000 217100 3052
rect 217968 3000 218020 3052
rect 224132 3000 224184 3052
rect 243544 3000 243596 3052
rect 269304 3000 269356 3052
rect 271144 3000 271196 3052
rect 337384 3000 337436 3052
rect 382372 3000 382424 3052
rect 410524 3000 410576 3052
rect 439412 3000 439464 3052
rect 478144 3000 478196 3052
rect 532240 3000 532292 3052
rect 159916 2932 159968 2984
rect 193312 2932 193364 2984
rect 221740 2932 221792 2984
rect 168196 2864 168248 2916
rect 188068 2864 188120 2916
rect 201500 2864 201552 2916
rect 208308 2864 208360 2916
rect 187240 2796 187292 2848
rect 194600 2796 194652 2848
rect 205088 2796 205140 2848
rect 209228 2796 209280 2848
rect 225236 2932 225288 2984
rect 232596 2932 232648 2984
rect 475384 2932 475436 2984
rect 525064 2932 525116 2984
rect 474004 2864 474056 2916
rect 517888 2864 517940 2916
rect 235264 2796 235316 2848
rect 336924 2796 336976 2848
rect 339684 2796 339736 2848
rect 343916 2796 343968 2848
rect 502340 2796 502392 2848
rect 503628 2796 503680 2848
rect 337016 2728 337068 2780
rect 340144 2728 340196 2780
rect 344008 2728 344060 2780
rect 400956 756 401008 808
rect 403716 756 403768 808
rect 92112 552 92164 604
rect 92388 552 92440 604
rect 178960 552 179012 604
rect 179328 552 179380 604
rect 238392 552 238444 604
rect 238668 552 238720 604
rect 275284 552 275336 604
rect 275376 552 275428 604
rect 280344 552 280396 604
rect 281264 552 281316 604
rect 305000 552 305052 604
rect 305184 552 305236 604
rect 307944 552 307996 604
rect 308588 552 308640 604
rect 323124 552 323176 604
rect 324044 552 324096 604
rect 325884 552 325936 604
rect 326436 552 326488 604
rect 332876 552 332928 604
rect 333612 552 333664 604
rect 337016 552 337068 604
rect 337108 552 337160 604
rect 340144 552 340196 604
rect 340696 552 340748 604
rect 344008 552 344060 604
rect 344284 552 344336 604
rect 416964 552 417016 604
rect 417976 552 418028 604
rect 425152 552 425204 604
rect 425336 552 425388 604
rect 441620 552 441672 604
rect 441804 552 441856 604
rect 444380 552 444432 604
rect 445392 552 445444 604
rect 448520 552 448572 604
rect 448980 552 449032 604
rect 455420 552 455472 604
rect 456064 552 456116 604
rect 456800 552 456852 604
rect 457260 552 457312 604
rect 499580 552 499632 604
rect 500132 552 500184 604
rect 506480 552 506532 604
rect 507216 552 507268 604
rect 510620 552 510672 604
rect 510804 552 510856 604
rect 513380 552 513432 604
rect 514392 552 514444 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 703474 8156 703520
rect 8036 703446 8156 703474
rect 8036 698290 8064 703446
rect 24320 699718 24348 703520
rect 40512 700466 40540 703520
rect 40500 700460 40552 700466
rect 40500 700402 40552 700408
rect 72988 699718 73016 703520
rect 89180 699718 89208 703520
rect 105464 700670 105492 703520
rect 133880 701004 133932 701010
rect 133880 700946 133932 700952
rect 133604 700936 133656 700942
rect 133604 700878 133656 700884
rect 133236 700868 133288 700874
rect 133236 700810 133288 700816
rect 132224 700800 132276 700806
rect 132224 700742 132276 700748
rect 131120 700732 131172 700738
rect 131120 700674 131172 700680
rect 105452 700664 105504 700670
rect 105452 700606 105504 700612
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 72424 699712 72476 699718
rect 72424 699654 72476 699660
rect 72976 699712 73028 699718
rect 72976 699654 73028 699660
rect 89168 699712 89220 699718
rect 89168 699654 89220 699660
rect 89628 699712 89680 699718
rect 89628 699654 89680 699660
rect 8024 698284 8076 698290
rect 8024 698226 8076 698232
rect 8208 698284 8260 698290
rect 8208 698226 8260 698232
rect 8220 695502 8248 698226
rect 7932 695496 7984 695502
rect 7932 695438 7984 695444
rect 8208 695496 8260 695502
rect 8208 695438 8260 695444
rect 7944 685914 7972 695438
rect 7932 685908 7984 685914
rect 7932 685850 7984 685856
rect 8116 685908 8168 685914
rect 8116 685850 8168 685856
rect 3790 682272 3846 682281
rect 3790 682207 3846 682216
rect 3804 681766 3832 682207
rect 3792 681760 3844 681766
rect 3792 681702 3844 681708
rect 8128 679046 8156 685850
rect 8116 679040 8168 679046
rect 8116 678982 8168 678988
rect 8024 678972 8076 678978
rect 8024 678914 8076 678920
rect 8036 673538 8064 678914
rect 8024 673532 8076 673538
rect 8024 673474 8076 673480
rect 8208 673532 8260 673538
rect 8208 673474 8260 673480
rect 3422 667992 3478 668001
rect 3422 667927 3478 667936
rect 3054 624880 3110 624889
rect 3054 624815 3110 624824
rect 3068 623830 3096 624815
rect 3056 623824 3108 623830
rect 3056 623766 3108 623772
rect 3146 481128 3202 481137
rect 3146 481063 3148 481072
rect 3200 481063 3202 481072
rect 3148 481034 3200 481040
rect 3238 452432 3294 452441
rect 3238 452367 3294 452376
rect 3252 451382 3280 452367
rect 3240 451376 3292 451382
rect 3240 451318 3292 451324
rect 3330 438016 3386 438025
rect 3330 437951 3386 437960
rect 3238 423736 3294 423745
rect 3238 423671 3294 423680
rect 3054 395040 3110 395049
rect 3054 394975 3110 394984
rect 2962 366208 3018 366217
rect 2962 366143 2964 366152
rect 3016 366143 3018 366152
rect 2964 366114 3016 366120
rect 2962 337512 3018 337521
rect 2962 337447 3018 337456
rect 2976 336802 3004 337447
rect 2964 336796 3016 336802
rect 2964 336738 3016 336744
rect 2962 323096 3018 323105
rect 2962 323031 3018 323040
rect 2976 322998 3004 323031
rect 2964 322992 3016 322998
rect 2964 322934 3016 322940
rect 2962 308816 3018 308825
rect 2962 308751 3018 308760
rect 2976 307834 3004 308751
rect 2964 307828 3016 307834
rect 2964 307770 3016 307776
rect 2962 294400 3018 294409
rect 2962 294335 3018 294344
rect 2976 294030 3004 294335
rect 2964 294024 3016 294030
rect 2964 293966 3016 293972
rect 2962 280120 3018 280129
rect 2962 280055 3018 280064
rect 2870 265704 2926 265713
rect 2870 265639 2926 265648
rect 2884 264994 2912 265639
rect 2872 264988 2924 264994
rect 2872 264930 2924 264936
rect 2870 251288 2926 251297
rect 2870 251223 2872 251232
rect 2924 251223 2926 251232
rect 2872 251194 2924 251200
rect 2870 237008 2926 237017
rect 2870 236943 2926 236952
rect 2778 222592 2834 222601
rect 2778 222527 2780 222536
rect 2832 222527 2834 222536
rect 2780 222498 2832 222504
rect 2780 210452 2832 210458
rect 2780 210394 2832 210400
rect 2792 201074 2820 210394
rect 2780 201068 2832 201074
rect 2780 201010 2832 201016
rect 2780 199844 2832 199850
rect 2780 199786 2832 199792
rect 2792 165073 2820 199786
rect 2778 165064 2834 165073
rect 2778 164999 2834 165008
rect 2884 154562 2912 236943
rect 2872 154556 2924 154562
rect 2872 154498 2924 154504
rect 2976 153202 3004 280055
rect 3068 210458 3096 394975
rect 3146 380624 3202 380633
rect 3146 380559 3202 380568
rect 3056 210452 3108 210458
rect 3056 210394 3108 210400
rect 3054 208176 3110 208185
rect 3054 208111 3110 208120
rect 3068 207058 3096 208111
rect 3056 207052 3108 207058
rect 3056 206994 3108 207000
rect 3054 193896 3110 193905
rect 3054 193831 3110 193840
rect 3068 155922 3096 193831
rect 3056 155916 3108 155922
rect 3056 155858 3108 155864
rect 2964 153196 3016 153202
rect 2964 153138 3016 153144
rect 3160 151774 3188 380559
rect 3252 190466 3280 423671
rect 3240 190460 3292 190466
rect 3240 190402 3292 190408
rect 3148 151768 3200 151774
rect 3148 151710 3200 151716
rect 3344 150414 3372 437951
rect 3332 150408 3384 150414
rect 3332 150350 3384 150356
rect 3436 146266 3464 667927
rect 8220 663762 8248 673474
rect 8036 663734 8248 663762
rect 8036 654158 8064 663734
rect 8024 654152 8076 654158
rect 8024 654094 8076 654100
rect 8208 654152 8260 654158
rect 8208 654094 8260 654100
rect 3514 653576 3570 653585
rect 3514 653511 3570 653520
rect 3528 186318 3556 653511
rect 8220 644450 8248 654094
rect 8036 644422 8248 644450
rect 8036 634846 8064 644422
rect 8024 634840 8076 634846
rect 8024 634782 8076 634788
rect 8208 634840 8260 634846
rect 8208 634782 8260 634788
rect 8220 625138 8248 634782
rect 8036 625110 8248 625138
rect 8036 615534 8064 625110
rect 8024 615528 8076 615534
rect 8024 615470 8076 615476
rect 8208 615528 8260 615534
rect 8208 615470 8260 615476
rect 3606 610464 3662 610473
rect 3606 610399 3662 610408
rect 3516 186312 3568 186318
rect 3516 186254 3568 186260
rect 3620 147626 3648 610399
rect 8220 605826 8248 615470
rect 8036 605798 8248 605826
rect 8036 596222 8064 605798
rect 8024 596216 8076 596222
rect 8208 596216 8260 596222
rect 8024 596158 8076 596164
rect 8128 596164 8208 596170
rect 8128 596158 8260 596164
rect 8128 596142 8248 596158
rect 3698 596048 3754 596057
rect 3698 595983 3754 595992
rect 3712 187678 3740 595983
rect 8128 591954 8156 596142
rect 8036 591926 8156 591954
rect 8036 582434 8064 591926
rect 7944 582406 8064 582434
rect 7944 579630 7972 582406
rect 7656 579624 7708 579630
rect 7656 579566 7708 579572
rect 7932 579624 7984 579630
rect 7932 579566 7984 579572
rect 7668 569974 7696 579566
rect 7656 569968 7708 569974
rect 7656 569910 7708 569916
rect 7840 569968 7892 569974
rect 7840 569910 7892 569916
rect 3882 567352 3938 567361
rect 3882 567287 3938 567296
rect 3790 553072 3846 553081
rect 3790 553007 3846 553016
rect 3700 187672 3752 187678
rect 3700 187614 3752 187620
rect 3700 179512 3752 179518
rect 3698 179480 3700 179489
rect 3752 179480 3754 179489
rect 3698 179415 3754 179424
rect 3804 148714 3832 553007
rect 3896 201142 3924 567287
rect 7852 563106 7880 569910
rect 7840 563100 7892 563106
rect 7840 563042 7892 563048
rect 7932 562964 7984 562970
rect 7932 562906 7984 562912
rect 7944 553330 7972 562906
rect 7944 553302 8064 553330
rect 8036 550594 8064 553302
rect 8024 550588 8076 550594
rect 8024 550530 8076 550536
rect 8116 550588 8168 550594
rect 8116 550530 8168 550536
rect 8128 541006 8156 550530
rect 8116 541000 8168 541006
rect 8116 540942 8168 540948
rect 8208 541000 8260 541006
rect 8208 540942 8260 540948
rect 3974 538656 4030 538665
rect 3974 538591 4030 538600
rect 3988 538490 4016 538591
rect 3976 538484 4028 538490
rect 3976 538426 4028 538432
rect 4804 538484 4856 538490
rect 4804 538426 4856 538432
rect 4066 509960 4122 509969
rect 4066 509895 4122 509904
rect 3974 495544 4030 495553
rect 3974 495479 4030 495488
rect 3884 201136 3936 201142
rect 3884 201078 3936 201084
rect 3884 198756 3936 198762
rect 3884 198698 3936 198704
rect 3792 148708 3844 148714
rect 3792 148650 3844 148656
rect 3608 147620 3660 147626
rect 3608 147562 3660 147568
rect 3424 146260 3476 146266
rect 3424 146202 3476 146208
rect 2780 136400 2832 136406
rect 2778 136368 2780 136377
rect 2832 136368 2834 136377
rect 2778 136303 2834 136312
rect 3238 122088 3294 122097
rect 3238 122023 3294 122032
rect 3252 120630 3280 122023
rect 3240 120624 3292 120630
rect 3240 120566 3292 120572
rect 3240 108996 3292 109002
rect 3240 108938 3292 108944
rect 3252 107681 3280 108938
rect 3238 107672 3294 107681
rect 3238 107607 3294 107616
rect 3424 93832 3476 93838
rect 3424 93774 3476 93780
rect 3436 93265 3464 93774
rect 3422 93256 3478 93265
rect 3422 93191 3478 93200
rect 3148 80028 3200 80034
rect 3148 79970 3200 79976
rect 3160 78985 3188 79970
rect 3146 78976 3202 78985
rect 3146 78911 3202 78920
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 3424 35896 3476 35902
rect 3422 35864 3424 35873
rect 3476 35864 3478 35873
rect 3422 35799 3478 35808
rect 2780 21480 2832 21486
rect 2778 21448 2780 21457
rect 2832 21448 2834 21457
rect 2778 21383 2834 21392
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 572 7608 624 7614
rect 572 7550 624 7556
rect 584 480 612 7550
rect 1688 480 1716 7686
rect 2872 7676 2924 7682
rect 2872 7618 2924 7624
rect 2884 480 2912 7618
rect 3896 7177 3924 198698
rect 3988 149054 4016 495479
rect 4080 201210 4108 509895
rect 4068 201204 4120 201210
rect 4068 201146 4120 201152
rect 4068 197396 4120 197402
rect 4068 197338 4120 197344
rect 3976 149048 4028 149054
rect 3976 148990 4028 148996
rect 4080 50153 4108 197338
rect 4816 188902 4844 538426
rect 8220 534018 8248 540942
rect 8128 533990 8248 534018
rect 8128 531321 8156 533990
rect 8114 531312 8170 531321
rect 8114 531247 8170 531256
rect 8390 531312 8446 531321
rect 8390 531247 8446 531256
rect 8404 521694 8432 531247
rect 8208 521688 8260 521694
rect 8208 521630 8260 521636
rect 8392 521688 8444 521694
rect 8392 521630 8444 521636
rect 8220 514706 8248 521630
rect 8128 514678 8248 514706
rect 8128 512009 8156 514678
rect 8114 512000 8170 512009
rect 8114 511935 8170 511944
rect 8390 512000 8446 512009
rect 8390 511935 8446 511944
rect 8404 502382 8432 511935
rect 8208 502376 8260 502382
rect 8208 502318 8260 502324
rect 8392 502376 8444 502382
rect 8392 502318 8444 502324
rect 8220 495394 8248 502318
rect 8128 495366 8248 495394
rect 8128 485858 8156 495366
rect 8116 485852 8168 485858
rect 8116 485794 8168 485800
rect 8208 485784 8260 485790
rect 8208 485726 8260 485732
rect 8220 483002 8248 485726
rect 7932 482996 7984 483002
rect 7932 482938 7984 482944
rect 8208 482996 8260 483002
rect 8208 482938 8260 482944
rect 4896 481092 4948 481098
rect 4896 481034 4948 481040
rect 4908 189038 4936 481034
rect 7944 473385 7972 482938
rect 7930 473376 7986 473385
rect 7930 473311 7986 473320
rect 8114 473376 8170 473385
rect 8114 473311 8170 473320
rect 8128 466478 8156 473311
rect 8116 466472 8168 466478
rect 8116 466414 8168 466420
rect 8208 466404 8260 466410
rect 8208 466346 8260 466352
rect 8220 456770 8248 466346
rect 8036 456742 8248 456770
rect 8036 454034 8064 456742
rect 7840 454028 7892 454034
rect 7840 453970 7892 453976
rect 8024 454028 8076 454034
rect 8024 453970 8076 453976
rect 7852 444446 7880 453970
rect 7840 444440 7892 444446
rect 7840 444382 7892 444388
rect 7932 444440 7984 444446
rect 7932 444382 7984 444388
rect 7944 437458 7972 444382
rect 7944 437430 8156 437458
rect 8128 427854 8156 437430
rect 8116 427848 8168 427854
rect 8116 427790 8168 427796
rect 8208 427780 8260 427786
rect 8208 427722 8260 427728
rect 8220 425066 8248 427722
rect 7932 425060 7984 425066
rect 7932 425002 7984 425008
rect 8208 425060 8260 425066
rect 8208 425002 8260 425008
rect 7944 415478 7972 425002
rect 7932 415472 7984 415478
rect 7932 415414 7984 415420
rect 8116 415472 8168 415478
rect 8116 415414 8168 415420
rect 8128 408542 8156 415414
rect 8116 408536 8168 408542
rect 8116 408478 8168 408484
rect 8208 408400 8260 408406
rect 8208 408342 8260 408348
rect 8220 400926 8248 408342
rect 8208 400920 8260 400926
rect 8208 400862 8260 400868
rect 8392 400920 8444 400926
rect 8392 400862 8444 400868
rect 8404 396098 8432 400862
rect 8024 396092 8076 396098
rect 8024 396034 8076 396040
rect 8392 396092 8444 396098
rect 8392 396034 8444 396040
rect 8036 394738 8064 396034
rect 8024 394732 8076 394738
rect 8024 394674 8076 394680
rect 8116 394732 8168 394738
rect 8116 394674 8168 394680
rect 8128 389230 8156 394674
rect 8116 389224 8168 389230
rect 8116 389166 8168 389172
rect 8208 389088 8260 389094
rect 8208 389030 8260 389036
rect 8220 379574 8248 389030
rect 8208 379568 8260 379574
rect 8208 379510 8260 379516
rect 8024 379500 8076 379506
rect 8024 379442 8076 379448
rect 8036 375358 8064 379442
rect 7840 375352 7892 375358
rect 7840 375294 7892 375300
rect 8024 375352 8076 375358
rect 8024 375294 8076 375300
rect 4988 366172 5040 366178
rect 4988 366114 5040 366120
rect 5000 191826 5028 366114
rect 7852 365770 7880 375294
rect 7840 365764 7892 365770
rect 7840 365706 7892 365712
rect 8116 365764 8168 365770
rect 8116 365706 8168 365712
rect 8128 360262 8156 365706
rect 8116 360256 8168 360262
rect 8116 360198 8168 360204
rect 8208 360188 8260 360194
rect 8208 360130 8260 360136
rect 8220 354686 8248 360130
rect 8208 354680 8260 354686
rect 8208 354622 8260 354628
rect 8392 354680 8444 354686
rect 8392 354622 8444 354628
rect 8404 345098 8432 354622
rect 8208 345092 8260 345098
rect 8208 345034 8260 345040
rect 8392 345092 8444 345098
rect 8392 345034 8444 345040
rect 8220 335322 8248 345034
rect 8036 335294 8248 335322
rect 8036 325718 8064 335294
rect 8024 325712 8076 325718
rect 8024 325654 8076 325660
rect 8208 325712 8260 325718
rect 8208 325654 8260 325660
rect 5080 322992 5132 322998
rect 5080 322934 5132 322940
rect 4988 191820 5040 191826
rect 4988 191762 5040 191768
rect 4896 189032 4948 189038
rect 4896 188974 4948 188980
rect 4804 188896 4856 188902
rect 4804 188838 4856 188844
rect 4804 158772 4856 158778
rect 4804 158714 4856 158720
rect 4160 155984 4212 155990
rect 4160 155926 4212 155932
rect 4172 150793 4200 155926
rect 4158 150784 4214 150793
rect 4158 150719 4214 150728
rect 4066 50144 4122 50153
rect 4066 50079 4122 50088
rect 4816 21486 4844 158714
rect 5092 153134 5120 322934
rect 8220 316010 8248 325654
rect 8036 315982 8248 316010
rect 5172 307828 5224 307834
rect 5172 307770 5224 307776
rect 5184 193186 5212 307770
rect 8036 306406 8064 315982
rect 8024 306400 8076 306406
rect 8024 306342 8076 306348
rect 8208 306400 8260 306406
rect 8208 306342 8260 306348
rect 8220 296698 8248 306342
rect 8036 296670 8248 296698
rect 8036 287094 8064 296670
rect 8024 287088 8076 287094
rect 8024 287030 8076 287036
rect 8208 287088 8260 287094
rect 8208 287030 8260 287036
rect 8220 277386 8248 287030
rect 8036 277358 8248 277386
rect 8036 267782 8064 277358
rect 8024 267776 8076 267782
rect 8208 267776 8260 267782
rect 8024 267718 8076 267724
rect 8128 267724 8208 267730
rect 8128 267718 8260 267724
rect 8128 267702 8248 267718
rect 5264 264988 5316 264994
rect 5264 264930 5316 264936
rect 5172 193180 5224 193186
rect 5172 193122 5224 193128
rect 5276 193118 5304 264930
rect 8128 263514 8156 267702
rect 8036 263486 8156 263514
rect 8036 253994 8064 263486
rect 7944 253966 8064 253994
rect 7944 251190 7972 253966
rect 7748 251184 7800 251190
rect 7748 251126 7800 251132
rect 7932 251184 7984 251190
rect 7932 251126 7984 251132
rect 7760 241534 7788 251126
rect 7748 241528 7800 241534
rect 7748 241470 7800 241476
rect 8024 241528 8076 241534
rect 8024 241470 8076 241476
rect 8036 234734 8064 241470
rect 8024 234728 8076 234734
rect 8024 234670 8076 234676
rect 7932 234592 7984 234598
rect 7932 234534 7984 234540
rect 7944 231810 7972 234534
rect 7748 231804 7800 231810
rect 7748 231746 7800 231752
rect 7932 231804 7984 231810
rect 7932 231746 7984 231752
rect 6184 222556 6236 222562
rect 6184 222498 6236 222504
rect 5356 196036 5408 196042
rect 5356 195978 5408 195984
rect 5264 193112 5316 193118
rect 5264 193054 5316 193060
rect 5080 153128 5132 153134
rect 5080 153070 5132 153076
rect 5368 136406 5396 195978
rect 6196 194478 6224 222498
rect 7760 222222 7788 231746
rect 7748 222216 7800 222222
rect 7748 222158 7800 222164
rect 8024 222216 8076 222222
rect 8024 222158 8076 222164
rect 8036 215422 8064 222158
rect 8024 215416 8076 215422
rect 8024 215358 8076 215364
rect 7932 215280 7984 215286
rect 7932 215222 7984 215228
rect 7944 212514 7972 215222
rect 7944 212486 8064 212514
rect 8036 205630 8064 212486
rect 8024 205624 8076 205630
rect 8024 205566 8076 205572
rect 8116 205556 8168 205562
rect 8116 205498 8168 205504
rect 8128 201482 8156 205498
rect 8024 201476 8076 201482
rect 8024 201418 8076 201424
rect 8116 201476 8168 201482
rect 8116 201418 8168 201424
rect 6184 194472 6236 194478
rect 6184 194414 6236 194420
rect 8036 193225 8064 201418
rect 14464 196104 14516 196110
rect 14464 196046 14516 196052
rect 8944 194608 8996 194614
rect 8944 194550 8996 194556
rect 8022 193216 8078 193225
rect 8022 193151 8078 193160
rect 8298 193216 8354 193225
rect 8298 193151 8354 193160
rect 8312 184890 8340 193151
rect 8300 184884 8352 184890
rect 8300 184826 8352 184832
rect 8956 179518 8984 194550
rect 9678 189000 9734 189009
rect 9678 188935 9734 188944
rect 9692 188902 9720 188935
rect 9680 188896 9732 188902
rect 9680 188838 9732 188844
rect 8944 179512 8996 179518
rect 8944 179454 8996 179460
rect 6920 153128 6972 153134
rect 6918 153096 6920 153105
rect 6972 153096 6974 153105
rect 6918 153031 6974 153040
rect 5356 136400 5408 136406
rect 5356 136342 5408 136348
rect 9588 117972 9640 117978
rect 9588 117914 9640 117920
rect 4804 21480 4856 21486
rect 4804 21422 4856 21428
rect 6460 9036 6512 9042
rect 6460 8978 6512 8984
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 3882 7168 3938 7177
rect 3882 7103 3938 7112
rect 4068 6180 4120 6186
rect 4068 6122 4120 6128
rect 4080 480 4108 6122
rect 5276 480 5304 8910
rect 6472 480 6500 8978
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7668 480 7696 7754
rect 9600 3534 9628 117914
rect 14476 93838 14504 196046
rect 19246 189000 19302 189009
rect 19246 188935 19302 188944
rect 19260 188902 19288 188935
rect 19248 188896 19300 188902
rect 19248 188838 19300 188844
rect 22100 188896 22152 188902
rect 22192 188896 22244 188902
rect 22152 188844 22192 188850
rect 22100 188838 22244 188844
rect 22112 188822 22232 188838
rect 16486 153096 16542 153105
rect 16486 153031 16542 153040
rect 16500 152998 16528 153031
rect 16488 152992 16540 152998
rect 16488 152934 16540 152940
rect 22192 148776 22244 148782
rect 22020 148724 22192 148730
rect 22020 148718 22244 148724
rect 22020 148714 22232 148718
rect 22008 148708 22232 148714
rect 22060 148702 22232 148708
rect 22008 148650 22060 148656
rect 24780 144906 24808 699654
rect 70216 524476 70268 524482
rect 70216 524418 70268 524424
rect 70124 407788 70176 407794
rect 70124 407730 70176 407736
rect 70136 370297 70164 407730
rect 70122 370288 70178 370297
rect 70122 370223 70178 370232
rect 70122 355600 70178 355609
rect 70122 355535 70178 355544
rect 70136 341465 70164 355535
rect 70228 348265 70256 524418
rect 70308 500268 70360 500274
rect 70308 500210 70360 500216
rect 70320 377913 70348 500210
rect 71688 398880 71740 398886
rect 71688 398822 71740 398828
rect 71504 396772 71556 396778
rect 71504 396714 71556 396720
rect 71516 385257 71544 396714
rect 71596 395752 71648 395758
rect 71596 395694 71648 395700
rect 71502 385248 71558 385257
rect 71502 385183 71558 385192
rect 70306 377904 70362 377913
rect 70306 377839 70362 377848
rect 71042 377904 71098 377913
rect 71042 377839 71098 377848
rect 70306 370288 70362 370297
rect 70306 370223 70362 370232
rect 70214 348256 70270 348265
rect 70214 348191 70270 348200
rect 70122 341456 70178 341465
rect 70122 341391 70178 341400
rect 67638 188864 67694 188873
rect 67638 188799 67640 188808
rect 67692 188799 67694 188808
rect 67640 188770 67692 188776
rect 41512 188760 41564 188766
rect 41340 188708 41512 188714
rect 60740 188760 60792 188766
rect 41340 188702 41564 188708
rect 60660 188708 60740 188714
rect 60660 188702 60792 188708
rect 41340 188698 41552 188702
rect 60660 188698 60780 188702
rect 41328 188692 41552 188698
rect 41380 188686 41552 188692
rect 48320 188692 48372 188698
rect 41328 188634 41380 188640
rect 48320 188634 48372 188640
rect 57888 188692 57940 188698
rect 57888 188634 57940 188640
rect 60648 188692 60780 188698
rect 60700 188686 60780 188692
rect 60648 188634 60700 188640
rect 48332 188562 48360 188634
rect 57900 188562 57928 188634
rect 48320 188556 48372 188562
rect 48320 188498 48372 188504
rect 57888 188556 57940 188562
rect 57888 188498 57940 188504
rect 41512 148776 41564 148782
rect 41340 148724 41512 148730
rect 41340 148718 41564 148724
rect 50988 148776 51040 148782
rect 56600 148776 56652 148782
rect 51040 148724 51120 148730
rect 50988 148718 51120 148724
rect 41340 148714 41552 148718
rect 26240 148708 26292 148714
rect 26240 148650 26292 148656
rect 35808 148708 35860 148714
rect 35808 148650 35860 148656
rect 41328 148708 41552 148714
rect 41380 148702 41552 148708
rect 51000 148714 51120 148718
rect 56520 148724 56600 148730
rect 64880 148776 64932 148782
rect 56520 148718 56652 148724
rect 64878 148744 64880 148753
rect 64932 148744 64934 148753
rect 56520 148714 56640 148718
rect 51000 148708 51132 148714
rect 51000 148702 51080 148708
rect 41328 148650 41380 148656
rect 51080 148650 51132 148656
rect 56508 148708 56640 148714
rect 56560 148702 56640 148708
rect 64878 148679 64934 148688
rect 56508 148650 56560 148656
rect 26252 148578 26280 148650
rect 35820 148578 35848 148650
rect 26240 148572 26292 148578
rect 26240 148514 26292 148520
rect 35808 148572 35860 148578
rect 35808 148514 35860 148520
rect 24768 144900 24820 144906
rect 24768 144842 24820 144848
rect 70320 118658 70348 370223
rect 70400 148844 70452 148850
rect 70400 148786 70452 148792
rect 70412 148753 70440 148786
rect 70398 148744 70454 148753
rect 70398 148679 70454 148688
rect 69848 118652 69900 118658
rect 69848 118594 69900 118600
rect 70308 118652 70360 118658
rect 70308 118594 70360 118600
rect 56508 118312 56560 118318
rect 56508 118254 56560 118260
rect 31668 118244 31720 118250
rect 31668 118186 31720 118192
rect 28908 118176 28960 118182
rect 28908 118118 28960 118124
rect 23388 118108 23440 118114
rect 23388 118050 23440 118056
rect 14464 93832 14516 93838
rect 14464 93774 14516 93780
rect 13636 9104 13688 9110
rect 13636 9046 13688 9052
rect 12440 4820 12492 4826
rect 12440 4762 12492 4768
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 8864 480 8892 3470
rect 10060 480 10088 3470
rect 11244 3460 11296 3466
rect 11244 3402 11296 3408
rect 11256 480 11284 3402
rect 12452 480 12480 4762
rect 13648 480 13676 9046
rect 18328 6316 18380 6322
rect 18328 6258 18380 6264
rect 17224 4888 17276 4894
rect 17224 4830 17276 4836
rect 14832 3664 14884 3670
rect 14832 3606 14884 3612
rect 14844 480 14872 3606
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 16040 480 16068 3538
rect 17236 480 17264 4830
rect 18340 480 18368 6258
rect 21916 4956 21968 4962
rect 21916 4898 21968 4904
rect 20720 3800 20772 3806
rect 20720 3742 20772 3748
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19536 480 19564 3674
rect 20732 480 20760 3742
rect 21928 480 21956 4898
rect 23400 3482 23428 118050
rect 26700 5024 26752 5030
rect 26700 4966 26752 4972
rect 25504 4140 25556 4146
rect 25504 4082 25556 4088
rect 24308 3868 24360 3874
rect 24308 3810 24360 3816
rect 23124 3454 23428 3482
rect 23124 480 23152 3454
rect 24320 480 24348 3810
rect 25516 480 25544 4082
rect 26712 480 26740 4966
rect 28920 3398 28948 118118
rect 30288 5092 30340 5098
rect 30288 5034 30340 5040
rect 29092 3936 29144 3942
rect 29092 3878 29144 3884
rect 27896 3392 27948 3398
rect 27896 3334 27948 3340
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 27908 480 27936 3334
rect 29104 480 29132 3878
rect 30300 480 30328 5034
rect 31680 626 31708 118186
rect 38568 10396 38620 10402
rect 38568 10338 38620 10344
rect 33876 9172 33928 9178
rect 33876 9114 33928 9120
rect 32680 6248 32732 6254
rect 32680 6190 32732 6196
rect 31496 598 31708 626
rect 31496 480 31524 598
rect 32692 480 32720 6190
rect 33888 480 33916 9114
rect 34980 8288 35032 8294
rect 34980 8230 35032 8236
rect 34992 480 35020 8230
rect 37372 5160 37424 5166
rect 37372 5102 37424 5108
rect 36176 4004 36228 4010
rect 36176 3946 36228 3952
rect 36188 480 36216 3946
rect 37384 480 37412 5102
rect 38580 480 38608 10338
rect 42708 10328 42760 10334
rect 42708 10270 42760 10276
rect 40960 9240 41012 9246
rect 40960 9182 41012 9188
rect 39764 6384 39816 6390
rect 39764 6326 39816 6332
rect 39776 480 39804 6326
rect 40972 480 41000 9182
rect 42720 4078 42748 10270
rect 45744 9580 45796 9586
rect 45744 9522 45796 9528
rect 44548 6452 44600 6458
rect 44548 6394 44600 6400
rect 42156 4072 42208 4078
rect 42156 4014 42208 4020
rect 42708 4072 42760 4078
rect 42708 4014 42760 4020
rect 43352 4072 43404 4078
rect 43352 4014 43404 4020
rect 42168 480 42196 4014
rect 43364 480 43392 4014
rect 44560 480 44588 6394
rect 45756 480 45784 9522
rect 55220 9376 55272 9382
rect 55220 9318 55272 9324
rect 51632 9308 51684 9314
rect 51632 9250 51684 9256
rect 48136 7880 48188 7886
rect 48136 7822 48188 7828
rect 46940 6520 46992 6526
rect 46940 6462 46992 6468
rect 46952 480 46980 6462
rect 48148 480 48176 7822
rect 50528 6588 50580 6594
rect 50528 6530 50580 6536
rect 49332 4548 49384 4554
rect 49332 4490 49384 4496
rect 49344 480 49372 4490
rect 50540 480 50568 6530
rect 51644 480 51672 9250
rect 54024 6656 54076 6662
rect 54024 6598 54076 6604
rect 52828 4480 52880 4486
rect 52828 4422 52880 4428
rect 52840 480 52868 4422
rect 54036 480 54064 6598
rect 55232 480 55260 9318
rect 56520 4842 56548 118254
rect 60648 118040 60700 118046
rect 60648 117982 60700 117988
rect 58808 9444 58860 9450
rect 58808 9386 58860 9392
rect 57612 6724 57664 6730
rect 57612 6666 57664 6672
rect 56428 4814 56548 4842
rect 56428 480 56456 4814
rect 57624 480 57652 6666
rect 58820 480 58848 9386
rect 60660 3398 60688 117982
rect 69860 117978 69888 118594
rect 69848 117972 69900 117978
rect 69848 117914 69900 117920
rect 71056 117502 71084 377839
rect 71608 362953 71636 395694
rect 71594 362944 71650 362953
rect 71594 362879 71650 362888
rect 71594 348256 71650 348265
rect 71594 348191 71650 348200
rect 71608 118386 71636 348191
rect 71596 118380 71648 118386
rect 71596 118322 71648 118328
rect 71700 117774 71728 398822
rect 72332 395548 72384 395554
rect 72332 395490 72384 395496
rect 72344 393009 72372 395490
rect 72330 393000 72386 393009
rect 72330 392935 72386 392944
rect 72436 183530 72464 699654
rect 85396 578332 85448 578338
rect 85396 578274 85448 578280
rect 84106 545864 84162 545873
rect 84106 545799 84162 545808
rect 84014 541512 84070 541521
rect 84014 541447 84070 541456
rect 83922 537160 83978 537169
rect 83922 537095 83978 537104
rect 83830 528728 83886 528737
rect 83830 528663 83886 528672
rect 82818 524920 82874 524929
rect 82818 524855 82874 524864
rect 82832 524482 82860 524855
rect 82820 524476 82872 524482
rect 82820 524418 82872 524424
rect 83844 497554 83872 528663
rect 83832 497548 83884 497554
rect 83832 497490 83884 497496
rect 75828 398132 75880 398138
rect 75828 398074 75880 398080
rect 75840 396250 75868 398074
rect 80796 397792 80848 397798
rect 80796 397734 80848 397740
rect 80808 396250 80836 397734
rect 75532 396222 75868 396250
rect 80500 396222 80836 396250
rect 83936 396030 83964 537095
rect 83924 396024 83976 396030
rect 83924 395966 83976 395972
rect 83936 395706 83964 395966
rect 83752 395690 83964 395706
rect 84028 395690 84056 541447
rect 84120 395758 84148 545799
rect 85302 533080 85358 533089
rect 85302 533015 85358 533024
rect 85316 521286 85344 533015
rect 85408 525609 85436 578274
rect 85580 578264 85632 578270
rect 85580 578206 85632 578212
rect 85488 549908 85540 549914
rect 85488 549850 85540 549856
rect 85394 525600 85450 525609
rect 85394 525535 85450 525544
rect 85304 521280 85356 521286
rect 85304 521222 85356 521228
rect 85500 398886 85528 549850
rect 85592 537781 85620 578206
rect 89168 553920 89220 553926
rect 89168 553862 89220 553868
rect 89180 551820 89208 553862
rect 89640 552702 89668 699654
rect 129648 696992 129700 696998
rect 129648 696934 129700 696940
rect 129556 650072 129608 650078
rect 129556 650014 129608 650020
rect 126244 583704 126296 583710
rect 126244 583646 126296 583652
rect 124864 583364 124916 583370
rect 124864 583306 124916 583312
rect 122748 578740 122800 578746
rect 122748 578682 122800 578688
rect 115952 578610 116072 578626
rect 115204 578604 115256 578610
rect 115204 578546 115256 578552
rect 115940 578604 116072 578610
rect 115992 578598 116072 578604
rect 115940 578546 115992 578552
rect 110328 575544 110380 575550
rect 110328 575486 110380 575492
rect 110340 554810 110368 575486
rect 109408 554804 109460 554810
rect 109408 554746 109460 554752
rect 110328 554804 110380 554810
rect 110328 554746 110380 554752
rect 92112 553988 92164 553994
rect 92112 553930 92164 553936
rect 89628 552696 89680 552702
rect 89628 552638 89680 552644
rect 92124 551820 92152 553930
rect 95056 553784 95108 553790
rect 95056 553726 95108 553732
rect 95068 551820 95096 553726
rect 100760 553716 100812 553722
rect 100760 553658 100812 553664
rect 97816 553512 97868 553518
rect 97816 553454 97868 553460
rect 97828 551820 97856 553454
rect 100772 551820 100800 553658
rect 106464 553648 106516 553654
rect 106464 553590 106516 553596
rect 103704 553580 103756 553586
rect 103704 553522 103756 553528
rect 103716 551820 103744 553522
rect 106476 551820 106504 553590
rect 109420 551820 109448 554746
rect 115112 553852 115164 553858
rect 115112 553794 115164 553800
rect 112352 553444 112404 553450
rect 112352 553386 112404 553392
rect 112364 551820 112392 553386
rect 115124 551820 115152 553794
rect 86406 549944 86462 549953
rect 86406 549879 86408 549888
rect 86460 549879 86462 549888
rect 86408 549850 86460 549856
rect 85578 537772 85634 537781
rect 85578 537707 85634 537716
rect 86604 518702 86632 520132
rect 89364 518906 89392 520132
rect 89352 518900 89404 518906
rect 89352 518842 89404 518848
rect 86592 518696 86644 518702
rect 86592 518638 86644 518644
rect 92308 518226 92336 520132
rect 92296 518220 92348 518226
rect 92296 518162 92348 518168
rect 95252 500274 95280 520132
rect 98012 518430 98040 520132
rect 99300 518770 99420 518786
rect 99288 518764 99432 518770
rect 99340 518758 99380 518764
rect 99288 518706 99340 518712
rect 99380 518706 99432 518712
rect 98000 518424 98052 518430
rect 98000 518366 98052 518372
rect 100956 518294 100984 520132
rect 103532 520118 103914 520146
rect 100944 518288 100996 518294
rect 100944 518230 100996 518236
rect 96528 500948 96580 500954
rect 96528 500890 96580 500896
rect 96540 500274 96568 500890
rect 103532 500886 103560 520118
rect 106660 518362 106688 520132
rect 109604 518838 109632 520132
rect 111812 520118 112562 520146
rect 109592 518832 109644 518838
rect 109592 518774 109644 518780
rect 109040 518696 109092 518702
rect 109132 518696 109184 518702
rect 109092 518644 109132 518650
rect 109040 518638 109184 518644
rect 109052 518622 109172 518638
rect 106648 518356 106700 518362
rect 106648 518298 106700 518304
rect 103520 500880 103572 500886
rect 103520 500822 103572 500828
rect 104808 500880 104860 500886
rect 104808 500822 104860 500828
rect 95240 500268 95292 500274
rect 95240 500210 95292 500216
rect 96528 500268 96580 500274
rect 96528 500210 96580 500216
rect 104820 407794 104848 500822
rect 111708 497888 111760 497894
rect 111708 497830 111760 497836
rect 108948 497616 109000 497622
rect 108948 497558 109000 497564
rect 104808 407788 104860 407794
rect 104808 407730 104860 407736
rect 85488 398880 85540 398886
rect 85488 398822 85540 398828
rect 85500 398750 85528 398822
rect 85488 398744 85540 398750
rect 85488 398686 85540 398692
rect 90272 398744 90324 398750
rect 90272 398686 90324 398692
rect 85948 397588 86000 397594
rect 85948 397530 86000 397536
rect 85960 396250 85988 397530
rect 85652 396222 85988 396250
rect 90284 396250 90312 398686
rect 100668 398200 100720 398206
rect 100668 398142 100720 398148
rect 95884 397656 95936 397662
rect 95884 397598 95936 397604
rect 95896 396250 95924 397598
rect 100680 396250 100708 398142
rect 106004 397724 106056 397730
rect 106004 397666 106056 397672
rect 106016 396250 106044 397666
rect 90284 396222 90620 396250
rect 95588 396222 95924 396250
rect 100556 396222 100708 396250
rect 105708 396222 106044 396250
rect 84568 396024 84620 396030
rect 84568 395966 84620 395972
rect 84580 395758 84608 395966
rect 96620 395888 96672 395894
rect 96618 395856 96620 395865
rect 96672 395856 96674 395865
rect 96618 395791 96674 395800
rect 99286 395856 99342 395865
rect 99286 395791 99342 395800
rect 99300 395758 99328 395791
rect 108960 395758 108988 497558
rect 111720 398886 111748 497830
rect 111812 497486 111840 520118
rect 115216 518838 115244 578546
rect 116044 578377 116072 578598
rect 119344 578536 119396 578542
rect 119344 578478 119396 578484
rect 116030 578368 116086 578377
rect 116030 578303 116086 578312
rect 115940 554804 115992 554810
rect 115940 554746 115992 554752
rect 115296 553988 115348 553994
rect 115296 553930 115348 553936
rect 113824 518832 113876 518838
rect 113824 518774 113876 518780
rect 115204 518832 115256 518838
rect 115204 518774 115256 518780
rect 111800 497480 111852 497486
rect 111800 497422 111852 497428
rect 110972 398880 111024 398886
rect 110972 398822 111024 398828
rect 111708 398880 111760 398886
rect 111708 398822 111760 398828
rect 110984 396250 111012 398822
rect 113836 398818 113864 518774
rect 115308 497894 115336 553930
rect 115296 497888 115348 497894
rect 115296 497830 115348 497836
rect 113548 398812 113600 398818
rect 113548 398754 113600 398760
rect 113824 398812 113876 398818
rect 113824 398754 113876 398760
rect 113560 398206 113588 398754
rect 113548 398200 113600 398206
rect 113548 398142 113600 398148
rect 115952 398138 115980 554746
rect 116032 553444 116084 553450
rect 116032 553386 116084 553392
rect 116044 498098 116072 553386
rect 118054 546544 118110 546553
rect 118054 546479 118110 546488
rect 117778 537432 117834 537441
rect 117778 537367 117834 537376
rect 117792 536858 117820 537367
rect 117780 536852 117832 536858
rect 117780 536794 117832 536800
rect 117778 533352 117834 533361
rect 117778 533287 117834 533296
rect 117792 532778 117820 533287
rect 117780 532772 117832 532778
rect 117780 532714 117832 532720
rect 117964 529916 118016 529922
rect 117964 529858 118016 529864
rect 117976 529689 118004 529858
rect 117962 529680 118018 529689
rect 117962 529615 118018 529624
rect 117318 521112 117374 521121
rect 117318 521047 117374 521056
rect 117332 520946 117360 521047
rect 117320 520940 117372 520946
rect 117320 520882 117372 520888
rect 116032 498092 116084 498098
rect 116032 498034 116084 498040
rect 116044 497622 116072 498034
rect 116032 497616 116084 497622
rect 116032 497558 116084 497564
rect 115940 398132 115992 398138
rect 115940 398074 115992 398080
rect 115848 397520 115900 397526
rect 115848 397462 115900 397468
rect 115860 396250 115888 397462
rect 117976 396778 118004 529615
rect 118068 498846 118096 546479
rect 118606 542464 118662 542473
rect 118606 542399 118608 542408
rect 118660 542399 118662 542408
rect 118608 542370 118660 542376
rect 119356 529922 119384 578478
rect 120724 553784 120776 553790
rect 120724 553726 120776 553732
rect 119344 529916 119396 529922
rect 119344 529858 119396 529864
rect 118606 525192 118662 525201
rect 118606 525127 118662 525136
rect 118620 525094 118648 525127
rect 118608 525088 118660 525094
rect 118608 525030 118660 525036
rect 118056 498840 118108 498846
rect 118056 498782 118108 498788
rect 120736 498030 120764 553726
rect 122760 519738 122788 578682
rect 122484 519710 122788 519738
rect 122484 518770 122512 519710
rect 122564 518900 122616 518906
rect 122564 518842 122616 518848
rect 122840 518900 122892 518906
rect 122840 518842 122892 518848
rect 122576 518786 122604 518842
rect 122852 518786 122880 518842
rect 122472 518764 122524 518770
rect 122576 518758 122880 518786
rect 122472 518706 122524 518712
rect 120724 498024 120776 498030
rect 120724 497966 120776 497972
rect 121368 498024 121420 498030
rect 121368 497966 121420 497972
rect 121380 398954 121408 497966
rect 120908 398948 120960 398954
rect 120908 398890 120960 398896
rect 121368 398948 121420 398954
rect 121368 398890 121420 398896
rect 117964 396772 118016 396778
rect 117964 396714 118016 396720
rect 120920 396250 120948 398890
rect 124128 397792 124180 397798
rect 124128 397734 124180 397740
rect 124140 397458 124168 397734
rect 124876 397458 124904 583306
rect 125692 578944 125744 578950
rect 125692 578886 125744 578892
rect 125704 578542 125732 578886
rect 125692 578536 125744 578542
rect 125692 578478 125744 578484
rect 125508 578400 125560 578406
rect 125506 578368 125508 578377
rect 125560 578368 125562 578377
rect 125506 578303 125562 578312
rect 125600 578332 125652 578338
rect 125600 578274 125652 578280
rect 125784 578332 125836 578338
rect 125784 578274 125836 578280
rect 125612 578218 125640 578274
rect 125796 578218 125824 578274
rect 125612 578190 125824 578218
rect 125968 497480 126020 497486
rect 125968 497422 126020 497428
rect 125692 398948 125744 398954
rect 125692 398890 125744 398896
rect 125600 398268 125652 398274
rect 125600 398210 125652 398216
rect 124128 397452 124180 397458
rect 124128 397394 124180 397400
rect 124864 397452 124916 397458
rect 124864 397394 124916 397400
rect 125612 396250 125640 398210
rect 110676 396222 111012 396250
rect 115644 396222 115888 396250
rect 120612 396222 120948 396250
rect 125580 396222 125640 396250
rect 84108 395752 84160 395758
rect 84108 395694 84160 395700
rect 84568 395752 84620 395758
rect 84568 395694 84620 395700
rect 99288 395752 99340 395758
rect 99288 395694 99340 395700
rect 108948 395752 109000 395758
rect 108948 395694 109000 395700
rect 83740 395684 83964 395690
rect 83792 395678 83964 395684
rect 84016 395684 84068 395690
rect 83740 395626 83792 395632
rect 84016 395626 84068 395632
rect 114468 340264 114520 340270
rect 114468 340206 114520 340212
rect 110328 340196 110380 340202
rect 110328 340138 110380 340144
rect 72588 340054 72924 340082
rect 77556 340054 77892 340082
rect 82524 340054 82768 340082
rect 87492 340054 87828 340082
rect 92460 340054 92796 340082
rect 97612 340054 97948 340082
rect 102580 340054 102916 340082
rect 107548 340054 107608 340082
rect 72896 337550 72924 340054
rect 72884 337544 72936 337550
rect 72884 337486 72936 337492
rect 77864 337482 77892 340054
rect 77852 337476 77904 337482
rect 77852 337418 77904 337424
rect 82740 336734 82768 340054
rect 87800 337414 87828 340054
rect 92768 337754 92796 340054
rect 97920 338026 97948 340054
rect 97908 338020 97960 338026
rect 97908 337962 97960 337968
rect 92756 337748 92808 337754
rect 92756 337690 92808 337696
rect 93768 337748 93820 337754
rect 93768 337690 93820 337696
rect 87788 337408 87840 337414
rect 87788 337350 87840 337356
rect 82728 336728 82780 336734
rect 82728 336670 82780 336676
rect 77206 188864 77262 188873
rect 77206 188799 77262 188808
rect 77220 188766 77248 188799
rect 77208 188760 77260 188766
rect 77208 188702 77260 188708
rect 79968 188760 80020 188766
rect 80060 188760 80112 188766
rect 80020 188708 80060 188714
rect 79968 188702 80112 188708
rect 79980 188686 80100 188702
rect 72424 183524 72476 183530
rect 72424 183466 72476 183472
rect 79968 148776 80020 148782
rect 80060 148776 80112 148782
rect 80020 148724 80060 148730
rect 79968 148718 80112 148724
rect 79980 148702 80100 148718
rect 82740 118522 82768 336670
rect 93780 202162 93808 337690
rect 93768 202156 93820 202162
rect 93768 202098 93820 202104
rect 86958 188864 87014 188873
rect 86958 188799 86960 188808
rect 87012 188799 87014 188808
rect 96342 188864 96398 188873
rect 96342 188799 96398 188808
rect 86960 188770 87012 188776
rect 96356 188578 96384 188799
rect 96528 188692 96580 188698
rect 96528 188634 96580 188640
rect 96540 188578 96568 188634
rect 96356 188550 96568 188578
rect 82820 153128 82872 153134
rect 82912 153128 82964 153134
rect 82872 153076 82912 153082
rect 82820 153070 82964 153076
rect 82832 153054 82952 153070
rect 84198 148880 84254 148889
rect 84198 148815 84200 148824
rect 84252 148815 84254 148824
rect 93582 148880 93638 148889
rect 93582 148815 93638 148824
rect 84200 148786 84252 148792
rect 93596 148594 93624 148815
rect 93768 148708 93820 148714
rect 93768 148650 93820 148656
rect 93780 148594 93808 148650
rect 93596 148566 93808 148594
rect 97920 118590 97948 337962
rect 102888 337754 102916 340054
rect 107580 338094 107608 340054
rect 107568 338088 107620 338094
rect 107568 338030 107620 338036
rect 102876 337748 102928 337754
rect 102876 337690 102928 337696
rect 103428 337748 103480 337754
rect 103428 337690 103480 337696
rect 99288 337476 99340 337482
rect 99288 337418 99340 337424
rect 97908 118584 97960 118590
rect 97908 118526 97960 118532
rect 82728 118516 82780 118522
rect 82728 118458 82780 118464
rect 82740 118046 82768 118458
rect 88340 118380 88392 118386
rect 88340 118322 88392 118328
rect 88352 118046 88380 118322
rect 82728 118040 82780 118046
rect 82728 117982 82780 117988
rect 88340 118040 88392 118046
rect 88340 117982 88392 117988
rect 71688 117768 71740 117774
rect 71688 117710 71740 117716
rect 73804 117768 73856 117774
rect 73804 117710 73856 117716
rect 79968 117768 80020 117774
rect 80020 117716 80192 117722
rect 79968 117710 80192 117716
rect 67548 117496 67600 117502
rect 67548 117438 67600 117444
rect 71044 117496 71096 117502
rect 71044 117438 71096 117444
rect 64788 10464 64840 10470
rect 64788 10406 64840 10412
rect 62396 9512 62448 9518
rect 62396 9454 62448 9460
rect 61200 6792 61252 6798
rect 61200 6734 61252 6740
rect 60004 3392 60056 3398
rect 60004 3334 60056 3340
rect 60648 3392 60700 3398
rect 60648 3334 60700 3340
rect 60016 480 60044 3334
rect 61212 480 61240 6734
rect 62408 480 62436 9454
rect 63592 7268 63644 7274
rect 63592 7210 63644 7216
rect 63604 480 63632 7210
rect 64800 480 64828 10406
rect 65984 5228 66036 5234
rect 65984 5170 66036 5176
rect 65996 480 66024 5170
rect 67560 4842 67588 117438
rect 72976 10532 73028 10538
rect 72976 10474 73028 10480
rect 68284 7948 68336 7954
rect 68284 7890 68336 7896
rect 67192 4814 67588 4842
rect 67192 480 67220 4814
rect 68296 480 68324 7890
rect 69480 5296 69532 5302
rect 69480 5238 69532 5244
rect 69492 480 69520 5238
rect 70676 4412 70728 4418
rect 70676 4354 70728 4360
rect 70688 480 70716 4354
rect 72988 3398 73016 10474
rect 73068 5364 73120 5370
rect 73068 5306 73120 5312
rect 71872 3392 71924 3398
rect 71872 3334 71924 3340
rect 72976 3392 73028 3398
rect 72976 3334 73028 3340
rect 71884 480 71912 3334
rect 73080 480 73108 5306
rect 73816 3398 73844 117710
rect 79980 117706 80192 117710
rect 79980 117700 80204 117706
rect 79980 117694 80152 117700
rect 80152 117642 80204 117648
rect 86960 117700 87012 117706
rect 86960 117642 87012 117648
rect 86972 117570 87000 117642
rect 86960 117564 87012 117570
rect 86960 117506 87012 117512
rect 86868 10668 86920 10674
rect 86868 10610 86920 10616
rect 79968 10600 80020 10606
rect 79968 10542 80020 10548
rect 77852 8832 77904 8838
rect 77852 8774 77904 8780
rect 75460 8016 75512 8022
rect 75460 7958 75512 7964
rect 73804 3392 73856 3398
rect 73804 3334 73856 3340
rect 74264 3392 74316 3398
rect 74264 3334 74316 3340
rect 74276 480 74304 3334
rect 75472 480 75500 7958
rect 76656 5432 76708 5438
rect 76656 5374 76708 5380
rect 76668 480 76696 5374
rect 77864 480 77892 8774
rect 79980 3058 80008 10542
rect 84936 8764 84988 8770
rect 84936 8706 84988 8712
rect 82636 8084 82688 8090
rect 82636 8026 82688 8032
rect 81440 5840 81492 5846
rect 81440 5782 81492 5788
rect 80244 5500 80296 5506
rect 80244 5442 80296 5448
rect 79048 3052 79100 3058
rect 79048 2994 79100 3000
rect 79968 3052 80020 3058
rect 79968 2994 80020 3000
rect 79060 480 79088 2994
rect 80256 480 80284 5442
rect 81452 480 81480 5782
rect 82648 480 82676 8026
rect 84200 6248 84252 6254
rect 84200 6190 84252 6196
rect 84212 6050 84240 6190
rect 84200 6044 84252 6050
rect 84200 5986 84252 5992
rect 83832 4752 83884 4758
rect 83832 4694 83884 4700
rect 83844 480 83872 4694
rect 84948 480 84976 8706
rect 86880 3398 86908 10610
rect 87328 4616 87380 4622
rect 87328 4558 87380 4564
rect 86132 3392 86184 3398
rect 86132 3334 86184 3340
rect 86868 3392 86920 3398
rect 86868 3334 86920 3340
rect 86144 480 86172 3334
rect 87340 480 87368 4558
rect 88352 3482 88380 117982
rect 96528 117836 96580 117842
rect 96528 117778 96580 117784
rect 96540 117570 96568 117778
rect 96528 117564 96580 117570
rect 96528 117506 96580 117512
rect 97920 117366 97948 118526
rect 99300 117881 99328 337418
rect 103440 202230 103468 337690
rect 103428 202224 103480 202230
rect 103428 202166 103480 202172
rect 99392 188698 99512 188714
rect 99380 188692 99524 188698
rect 99432 188686 99472 188692
rect 99380 188634 99432 188640
rect 99472 188634 99524 188640
rect 99392 148714 99512 148730
rect 99380 148708 99524 148714
rect 99432 148702 99472 148708
rect 99380 148650 99432 148656
rect 99472 148650 99524 148656
rect 107580 118250 107608 338030
rect 110340 118386 110368 340138
rect 112516 340054 112852 340082
rect 112824 337958 112852 340054
rect 112812 337952 112864 337958
rect 112812 337894 112864 337900
rect 113088 337952 113140 337958
rect 113088 337894 113140 337900
rect 110328 118380 110380 118386
rect 110328 118322 110380 118328
rect 107568 118244 107620 118250
rect 107568 118186 107620 118192
rect 107580 117910 107608 118186
rect 110340 118114 110368 118322
rect 113100 118250 113128 337894
rect 113088 118244 113140 118250
rect 113088 118186 113140 118192
rect 110328 118108 110380 118114
rect 110328 118050 110380 118056
rect 107568 117904 107620 117910
rect 97998 117872 98054 117881
rect 99286 117872 99342 117881
rect 97998 117807 98054 117816
rect 99196 117836 99248 117842
rect 92388 117360 92440 117366
rect 92388 117302 92440 117308
rect 97908 117360 97960 117366
rect 97908 117302 97960 117308
rect 89720 8152 89772 8158
rect 89720 8094 89772 8100
rect 88352 3454 88564 3482
rect 88536 480 88564 3454
rect 89732 480 89760 8094
rect 90916 4684 90968 4690
rect 90916 4626 90968 4632
rect 90928 480 90956 4626
rect 92400 610 92428 117302
rect 94504 9648 94556 9654
rect 94504 9590 94556 9596
rect 93308 3392 93360 3398
rect 93308 3334 93360 3340
rect 92112 604 92164 610
rect 92112 546 92164 552
rect 92388 604 92440 610
rect 92388 546 92440 552
rect 92124 480 92152 546
rect 93320 480 93348 3334
rect 94516 480 94544 9590
rect 95700 8696 95752 8702
rect 95700 8638 95752 8644
rect 95712 480 95740 8638
rect 96896 8220 96948 8226
rect 96896 8162 96948 8168
rect 96908 480 96936 8162
rect 98012 7546 98040 117807
rect 107568 117846 107620 117852
rect 99286 117807 99342 117816
rect 99196 117778 99248 117784
rect 99208 117722 99236 117778
rect 99472 117768 99524 117774
rect 99208 117716 99472 117722
rect 99208 117710 99524 117716
rect 99208 117694 99512 117710
rect 113100 117366 113128 118186
rect 114480 118182 114508 340206
rect 117668 340054 118004 340082
rect 122636 340054 122696 340082
rect 117976 337618 118004 340054
rect 122668 337890 122696 340054
rect 122656 337884 122708 337890
rect 122656 337826 122708 337832
rect 117964 337612 118016 337618
rect 117964 337554 118016 337560
rect 117228 337408 117280 337414
rect 117228 337350 117280 337356
rect 115938 188864 115994 188873
rect 115938 188799 115940 188808
rect 115992 188799 115994 188808
rect 115940 188770 115992 188776
rect 116308 152992 116360 152998
rect 116308 152934 116360 152940
rect 116320 152862 116348 152934
rect 116308 152856 116360 152862
rect 116308 152798 116360 152804
rect 115952 148974 116072 149002
rect 115952 148918 115980 148974
rect 115940 148912 115992 148918
rect 115940 148854 115992 148860
rect 116044 148646 116072 148974
rect 116032 148640 116084 148646
rect 116032 148582 116084 148588
rect 114468 118176 114520 118182
rect 114468 118118 114520 118124
rect 114480 117434 114508 118118
rect 115204 118108 115256 118114
rect 115204 118050 115256 118056
rect 114468 117428 114520 117434
rect 114468 117370 114520 117376
rect 109684 117360 109736 117366
rect 109684 117302 109736 117308
rect 113088 117360 113140 117366
rect 113088 117302 113140 117308
rect 98092 8900 98144 8906
rect 98092 8842 98144 8848
rect 98000 7540 98052 7546
rect 98000 7482 98052 7488
rect 98104 480 98132 8842
rect 99288 7540 99340 7546
rect 99288 7482 99340 7488
rect 99300 480 99328 7482
rect 101588 6860 101640 6866
rect 101588 6802 101640 6808
rect 100484 3324 100536 3330
rect 100484 3266 100536 3272
rect 100496 480 100524 3266
rect 101600 480 101628 6802
rect 103428 6248 103480 6254
rect 103428 6190 103480 6196
rect 102784 6112 102836 6118
rect 102784 6054 102836 6060
rect 102796 480 102824 6054
rect 103440 6050 103468 6190
rect 103428 6044 103480 6050
rect 103428 5986 103480 5992
rect 105176 6044 105228 6050
rect 105176 5986 105228 5992
rect 103980 3256 104032 3262
rect 103980 3198 104032 3204
rect 103992 480 104020 3198
rect 105188 480 105216 5986
rect 106372 5976 106424 5982
rect 106372 5918 106424 5924
rect 106384 480 106412 5918
rect 108764 5908 108816 5914
rect 108764 5850 108816 5856
rect 107568 3120 107620 3126
rect 107568 3062 107620 3068
rect 107580 480 107608 3062
rect 108776 480 108804 5850
rect 109696 5846 109724 117302
rect 114468 10736 114520 10742
rect 114468 10678 114520 10684
rect 111156 7540 111208 7546
rect 111156 7482 111208 7488
rect 109960 7336 110012 7342
rect 109960 7278 110012 7284
rect 109684 5840 109736 5846
rect 109684 5782 109736 5788
rect 109972 480 110000 7278
rect 111168 480 111196 7482
rect 113180 6248 113232 6254
rect 113180 6190 113232 6196
rect 112352 5840 112404 5846
rect 112352 5782 112404 5788
rect 112364 480 112392 5782
rect 113192 5642 113220 6190
rect 113180 5636 113232 5642
rect 113180 5578 113232 5584
rect 114480 3194 114508 10678
rect 115216 8294 115244 118050
rect 117240 117745 117268 337350
rect 122668 321586 122696 337826
rect 122576 321570 122696 321586
rect 122564 321564 122696 321570
rect 122616 321558 122696 321564
rect 122748 321564 122800 321570
rect 122564 321506 122616 321512
rect 122748 321506 122800 321512
rect 122576 321475 122604 321506
rect 122760 318782 122788 321506
rect 122472 318776 122524 318782
rect 122472 318718 122524 318724
rect 122748 318776 122800 318782
rect 122748 318718 122800 318724
rect 122484 309194 122512 318718
rect 122472 309188 122524 309194
rect 122472 309130 122524 309136
rect 122656 309188 122708 309194
rect 122656 309130 122708 309136
rect 122668 302240 122696 309130
rect 122576 302212 122696 302240
rect 122576 302138 122604 302212
rect 122576 302110 122696 302138
rect 122668 292584 122696 302110
rect 122668 292556 122788 292584
rect 122760 292482 122788 292556
rect 122668 292454 122788 292482
rect 122668 282962 122696 292454
rect 122576 282934 122696 282962
rect 122576 282826 122604 282934
rect 122576 282798 122696 282826
rect 122668 273306 122696 282798
rect 122668 273278 122788 273306
rect 122760 273170 122788 273278
rect 122668 273142 122788 273170
rect 122668 263650 122696 273142
rect 122576 263622 122696 263650
rect 122576 263514 122604 263622
rect 122576 263486 122696 263514
rect 122668 253994 122696 263486
rect 122668 253966 122788 253994
rect 122760 253858 122788 253966
rect 122668 253830 122788 253858
rect 122668 244338 122696 253830
rect 122576 244310 122696 244338
rect 122576 244202 122604 244310
rect 122576 244174 122696 244202
rect 122668 234682 122696 244174
rect 122668 234654 122788 234682
rect 122760 234546 122788 234654
rect 122668 234518 122788 234546
rect 122668 225026 122696 234518
rect 122576 224998 122696 225026
rect 122576 224942 122604 224998
rect 122564 224936 122616 224942
rect 122564 224878 122616 224884
rect 122748 224936 122800 224942
rect 122748 224878 122800 224884
rect 122760 215422 122788 224878
rect 122748 215416 122800 215422
rect 122748 215358 122800 215364
rect 122656 215280 122708 215286
rect 122656 215222 122708 215228
rect 122668 212537 122696 215222
rect 122654 212528 122710 212537
rect 122654 212463 122710 212472
rect 122838 212528 122894 212537
rect 122838 212463 122894 212472
rect 122852 205442 122880 212463
rect 122668 205414 122880 205442
rect 122668 202881 122696 205414
rect 122654 202872 122710 202881
rect 122654 202807 122710 202816
rect 122930 202872 122986 202881
rect 122930 202807 122986 202816
rect 122944 195906 122972 202807
rect 122748 195900 122800 195906
rect 122748 195842 122800 195848
rect 122932 195900 122984 195906
rect 122932 195842 122984 195848
rect 122760 186402 122788 195842
rect 125506 188864 125562 188873
rect 125506 188799 125562 188808
rect 125520 188766 125548 188799
rect 125508 188760 125560 188766
rect 125508 188702 125560 188708
rect 122576 186374 122788 186402
rect 122576 186266 122604 186374
rect 122576 186238 122696 186266
rect 122668 183546 122696 186238
rect 122668 183518 122788 183546
rect 122760 176730 122788 183518
rect 122748 176724 122800 176730
rect 122748 176666 122800 176672
rect 122656 176588 122708 176594
rect 122656 176530 122708 176536
rect 122668 167090 122696 176530
rect 122576 167062 122696 167090
rect 122576 161498 122604 167062
rect 122564 161492 122616 161498
rect 122564 161434 122616 161440
rect 122748 161492 122800 161498
rect 122748 161434 122800 161440
rect 122760 147558 122788 161434
rect 122564 147552 122616 147558
rect 122564 147494 122616 147500
rect 122748 147552 122800 147558
rect 122748 147494 122800 147500
rect 122576 138038 122604 147494
rect 122564 138032 122616 138038
rect 122564 137974 122616 137980
rect 122656 137896 122708 137902
rect 122656 137838 122708 137844
rect 120724 118448 120776 118454
rect 120724 118390 120776 118396
rect 117226 117736 117282 117745
rect 117226 117671 117282 117680
rect 117240 117337 117268 117671
rect 115938 117328 115994 117337
rect 115938 117263 115994 117272
rect 117226 117328 117282 117337
rect 117226 117263 117282 117272
rect 115204 8288 115256 8294
rect 115204 8230 115256 8236
rect 115952 3194 115980 117263
rect 120632 8628 120684 8634
rect 120632 8570 120684 8576
rect 118240 8288 118292 8294
rect 118240 8230 118292 8236
rect 116032 5772 116084 5778
rect 116032 5714 116084 5720
rect 113548 3188 113600 3194
rect 113548 3130 113600 3136
rect 114468 3188 114520 3194
rect 114468 3130 114520 3136
rect 115940 3188 115992 3194
rect 115940 3130 115992 3136
rect 113560 480 113588 3130
rect 114744 3052 114796 3058
rect 114744 2994 114796 3000
rect 114756 480 114784 2994
rect 116044 2938 116072 5714
rect 117136 3188 117188 3194
rect 117136 3130 117188 3136
rect 115952 2910 116072 2938
rect 115952 480 115980 2910
rect 117148 480 117176 3130
rect 118252 480 118280 8230
rect 119436 5704 119488 5710
rect 119436 5646 119488 5652
rect 119448 480 119476 5646
rect 120644 480 120672 8570
rect 120736 4418 120764 118390
rect 122668 117842 122696 137838
rect 125704 118454 125732 398890
rect 125784 397452 125836 397458
rect 125784 397394 125836 397400
rect 125692 118448 125744 118454
rect 125796 118425 125824 397394
rect 125876 395752 125928 395758
rect 125876 395694 125928 395700
rect 125692 118390 125744 118396
rect 125782 118416 125838 118425
rect 125782 118351 125838 118360
rect 125796 118130 125824 118351
rect 125888 118318 125916 395694
rect 125980 336734 126008 497422
rect 126060 398880 126112 398886
rect 126060 398822 126112 398828
rect 126072 340882 126100 398822
rect 126256 397662 126284 583646
rect 129004 583432 129056 583438
rect 129004 583374 129056 583380
rect 129016 553858 129044 583374
rect 129096 578604 129148 578610
rect 129096 578546 129148 578552
rect 128452 553852 128504 553858
rect 128452 553794 128504 553800
rect 129004 553852 129056 553858
rect 129004 553794 129056 553800
rect 128464 553382 128492 553794
rect 128452 553376 128504 553382
rect 128452 553318 128504 553324
rect 128636 553376 128688 553382
rect 128636 553318 128688 553324
rect 128648 543862 128676 553318
rect 129004 552696 129056 552702
rect 129004 552638 129056 552644
rect 128636 543856 128688 543862
rect 128636 543798 128688 543804
rect 128544 543720 128596 543726
rect 128544 543662 128596 543668
rect 128556 540954 128584 543662
rect 128464 540926 128584 540954
rect 128464 534138 128492 540926
rect 128452 534132 128504 534138
rect 128452 534074 128504 534080
rect 128544 534064 128596 534070
rect 128544 534006 128596 534012
rect 128556 531350 128584 534006
rect 128452 531344 128504 531350
rect 128452 531286 128504 531292
rect 128544 531344 128596 531350
rect 128544 531286 128596 531292
rect 128360 525088 128412 525094
rect 128360 525030 128412 525036
rect 128372 524226 128400 525030
rect 128464 524482 128492 531286
rect 128452 524476 128504 524482
rect 128452 524418 128504 524424
rect 128636 524340 128688 524346
rect 128636 524282 128688 524288
rect 128372 524198 128584 524226
rect 128452 521620 128504 521626
rect 128452 521562 128504 521568
rect 128464 520946 128492 521562
rect 128452 520940 128504 520946
rect 128452 520882 128504 520888
rect 128360 518968 128412 518974
rect 128360 518910 128412 518916
rect 127716 518832 127768 518838
rect 127716 518774 127768 518780
rect 127624 518424 127676 518430
rect 127624 518366 127676 518372
rect 127072 518220 127124 518226
rect 127072 518162 127124 518168
rect 126980 398812 127032 398818
rect 126980 398754 127032 398760
rect 126244 397656 126296 397662
rect 126244 397598 126296 397604
rect 126060 340876 126112 340882
rect 126060 340818 126112 340824
rect 126072 340270 126100 340818
rect 126060 340264 126112 340270
rect 126060 340206 126112 340212
rect 125968 336728 126020 336734
rect 125968 336670 126020 336676
rect 125876 118312 125928 118318
rect 126256 118289 126284 397598
rect 126336 396772 126388 396778
rect 126336 396714 126388 396720
rect 126348 385014 126376 396714
rect 126888 395684 126940 395690
rect 126888 395626 126940 395632
rect 126900 391950 126928 395626
rect 126888 391944 126940 391950
rect 126888 391886 126940 391892
rect 126900 386374 126928 391886
rect 126888 386368 126940 386374
rect 126888 386310 126940 386316
rect 126336 385008 126388 385014
rect 126336 384950 126388 384956
rect 126992 118697 127020 398754
rect 127084 338026 127112 518162
rect 127636 497622 127664 518366
rect 127624 497616 127676 497622
rect 127624 497558 127676 497564
rect 127164 497548 127216 497554
rect 127164 497490 127216 497496
rect 127072 338020 127124 338026
rect 127072 337962 127124 337968
rect 127176 337958 127204 497490
rect 127256 398132 127308 398138
rect 127256 398074 127308 398080
rect 127268 340814 127296 398074
rect 127624 397520 127676 397526
rect 127624 397462 127676 397468
rect 127256 340808 127308 340814
rect 127256 340750 127308 340756
rect 127268 340202 127296 340750
rect 127256 340196 127308 340202
rect 127256 340138 127308 340144
rect 127164 337952 127216 337958
rect 127164 337894 127216 337900
rect 127636 201618 127664 397462
rect 127728 340746 127756 518774
rect 128372 509250 128400 518910
rect 128360 509244 128412 509250
rect 128360 509186 128412 509192
rect 128360 499588 128412 499594
rect 128360 499530 128412 499536
rect 128268 497956 128320 497962
rect 128268 497898 128320 497904
rect 128280 497622 128308 497898
rect 128268 497616 128320 497622
rect 128268 497558 128320 497564
rect 127808 407176 127860 407182
rect 127808 407118 127860 407124
rect 127820 398818 127848 407118
rect 127808 398812 127860 398818
rect 127808 398754 127860 398760
rect 128280 398274 128308 497558
rect 128372 489870 128400 499530
rect 128360 489864 128412 489870
rect 128360 489806 128412 489812
rect 128360 480344 128412 480350
rect 128360 480286 128412 480292
rect 128372 431934 128400 480286
rect 128360 431928 128412 431934
rect 128360 431870 128412 431876
rect 128360 422408 128412 422414
rect 128360 422350 128412 422356
rect 128268 398268 128320 398274
rect 128268 398210 128320 398216
rect 128268 398132 128320 398138
rect 128268 398074 128320 398080
rect 128280 397594 128308 398074
rect 128268 397588 128320 397594
rect 128268 397530 128320 397536
rect 127716 340740 127768 340746
rect 127716 340682 127768 340688
rect 127728 337890 127756 340682
rect 127716 337884 127768 337890
rect 127716 337826 127768 337832
rect 128176 337612 128228 337618
rect 128176 337554 128228 337560
rect 128084 260840 128136 260846
rect 128084 260782 128136 260788
rect 128096 251297 128124 260782
rect 128082 251288 128138 251297
rect 128082 251223 128138 251232
rect 127624 201612 127676 201618
rect 127624 201554 127676 201560
rect 126978 118688 127034 118697
rect 126978 118623 127034 118632
rect 126888 118312 126940 118318
rect 125876 118254 125928 118260
rect 126242 118280 126298 118289
rect 126888 118254 126940 118260
rect 126242 118215 126298 118224
rect 125520 118102 125824 118130
rect 122840 117972 122892 117978
rect 122840 117914 122892 117920
rect 122104 117836 122156 117842
rect 122104 117778 122156 117784
rect 122656 117836 122708 117842
rect 122656 117778 122708 117784
rect 121828 7472 121880 7478
rect 121828 7414 121880 7420
rect 120724 4412 120776 4418
rect 120724 4354 120776 4360
rect 120816 4412 120868 4418
rect 120816 4354 120868 4360
rect 120828 4146 120856 4354
rect 120816 4140 120868 4146
rect 120816 4082 120868 4088
rect 121840 480 121868 7414
rect 122116 4486 122144 117778
rect 122852 117774 122880 117914
rect 122840 117768 122892 117774
rect 122840 117710 122892 117716
rect 122748 6248 122800 6254
rect 122748 6190 122800 6196
rect 122760 5642 122788 6190
rect 122748 5636 122800 5642
rect 122748 5578 122800 5584
rect 123024 5636 123076 5642
rect 123024 5578 123076 5584
rect 122104 4480 122156 4486
rect 122104 4422 122156 4428
rect 123036 480 123064 5578
rect 125416 4140 125468 4146
rect 125416 4082 125468 4088
rect 124220 3052 124272 3058
rect 124220 2994 124272 3000
rect 124232 480 124260 2994
rect 125428 480 125456 4082
rect 125520 3058 125548 118102
rect 126256 8498 126284 118215
rect 126900 117774 126928 118254
rect 126992 118114 127020 118623
rect 128188 118114 128216 337554
rect 128280 118726 128308 397530
rect 128372 393310 128400 422350
rect 128360 393304 128412 393310
rect 128360 393246 128412 393252
rect 128360 383716 128412 383722
rect 128360 383658 128412 383664
rect 128372 373998 128400 383658
rect 128360 373992 128412 373998
rect 128360 373934 128412 373940
rect 128464 373289 128492 520882
rect 128556 387977 128584 524198
rect 128648 518974 128676 524282
rect 128636 518968 128688 518974
rect 128636 518910 128688 518916
rect 128636 509244 128688 509250
rect 128636 509186 128688 509192
rect 128648 499594 128676 509186
rect 128636 499588 128688 499594
rect 128636 499530 128688 499536
rect 128636 489864 128688 489870
rect 128636 489806 128688 489812
rect 128648 480350 128676 489806
rect 128636 480344 128688 480350
rect 128636 480286 128688 480292
rect 128636 431928 128688 431934
rect 128636 431870 128688 431876
rect 128648 422414 128676 431870
rect 128636 422408 128688 422414
rect 128636 422350 128688 422356
rect 128636 393304 128688 393310
rect 128636 393246 128688 393252
rect 128542 387968 128598 387977
rect 128542 387903 128598 387912
rect 128648 383722 128676 393246
rect 128636 383716 128688 383722
rect 128636 383658 128688 383664
rect 128820 374060 128872 374066
rect 128820 374002 128872 374008
rect 128544 373992 128596 373998
rect 128544 373934 128596 373940
rect 128450 373280 128506 373289
rect 128450 373215 128506 373224
rect 128464 372745 128492 373215
rect 128450 372736 128506 372745
rect 128450 372671 128506 372680
rect 128556 369850 128584 373934
rect 128544 369844 128596 369850
rect 128544 369786 128596 369792
rect 128636 369776 128688 369782
rect 128636 369718 128688 369724
rect 128648 358737 128676 369718
rect 128832 360262 128860 374002
rect 128910 365936 128966 365945
rect 128910 365871 128966 365880
rect 128924 365702 128952 365871
rect 128912 365696 128964 365702
rect 128912 365638 128964 365644
rect 128820 360256 128872 360262
rect 128820 360198 128872 360204
rect 128634 358728 128690 358737
rect 128690 358686 128768 358714
rect 128634 358663 128690 358672
rect 128740 347954 128768 358686
rect 128728 347948 128780 347954
rect 128728 347890 128780 347896
rect 128636 347812 128688 347818
rect 128636 347754 128688 347760
rect 128728 347812 128780 347818
rect 128728 347754 128780 347760
rect 128648 342938 128676 347754
rect 128740 345574 128768 347754
rect 128728 345568 128780 345574
rect 128728 345510 128780 345516
rect 128818 343632 128874 343641
rect 128818 343567 128874 343576
rect 128464 342910 128676 342938
rect 128464 338178 128492 342910
rect 128832 342514 128860 343567
rect 128820 342508 128872 342514
rect 128820 342450 128872 342456
rect 128464 338150 128584 338178
rect 128556 335345 128584 338150
rect 128728 336048 128780 336054
rect 128728 335990 128780 335996
rect 128358 335336 128414 335345
rect 128358 335271 128414 335280
rect 128542 335336 128598 335345
rect 128542 335271 128598 335280
rect 128372 325718 128400 335271
rect 128740 327078 128768 335990
rect 128728 327072 128780 327078
rect 128728 327014 128780 327020
rect 128360 325712 128412 325718
rect 128360 325654 128412 325660
rect 128452 325712 128504 325718
rect 128452 325654 128504 325660
rect 128464 311794 128492 325654
rect 128464 311766 128676 311794
rect 128648 302274 128676 311766
rect 128728 311636 128780 311642
rect 128728 311578 128780 311584
rect 128740 307086 128768 311578
rect 128728 307080 128780 307086
rect 128728 307022 128780 307028
rect 128648 302246 128860 302274
rect 128832 299538 128860 302246
rect 128636 299532 128688 299538
rect 128636 299474 128688 299480
rect 128820 299532 128872 299538
rect 128820 299474 128872 299480
rect 128648 290494 128676 299474
rect 128728 297424 128780 297430
rect 128728 297366 128780 297372
rect 128452 290488 128504 290494
rect 128452 290430 128504 290436
rect 128636 290488 128688 290494
rect 128636 290430 128688 290436
rect 128464 282826 128492 290430
rect 128740 287774 128768 297366
rect 128728 287768 128780 287774
rect 128728 287710 128780 287716
rect 128464 282798 128676 282826
rect 128648 280158 128676 282798
rect 128452 280152 128504 280158
rect 128452 280094 128504 280100
rect 128636 280152 128688 280158
rect 128636 280094 128688 280100
rect 128464 270570 128492 280094
rect 128728 274304 128780 274310
rect 128728 274246 128780 274252
rect 128452 270564 128504 270570
rect 128452 270506 128504 270512
rect 128636 270564 128688 270570
rect 128636 270506 128688 270512
rect 128648 263514 128676 270506
rect 128740 268462 128768 274246
rect 128728 268456 128780 268462
rect 128728 268398 128780 268404
rect 128556 263486 128676 263514
rect 128556 260846 128584 263486
rect 128544 260840 128596 260846
rect 128544 260782 128596 260788
rect 128728 258800 128780 258806
rect 128728 258742 128780 258748
rect 128450 251288 128506 251297
rect 128450 251223 128506 251232
rect 128464 244202 128492 251223
rect 128740 249150 128768 258742
rect 128728 249144 128780 249150
rect 128728 249086 128780 249092
rect 128464 244174 128584 244202
rect 128556 241482 128584 244174
rect 128556 241454 128860 241482
rect 128728 239488 128780 239494
rect 128728 239430 128780 239436
rect 128636 231872 128688 231878
rect 128636 231814 128688 231820
rect 128648 224890 128676 231814
rect 128740 229770 128768 239430
rect 128832 231878 128860 241454
rect 128820 231872 128872 231878
rect 128820 231814 128872 231820
rect 128728 229764 128780 229770
rect 128728 229706 128780 229712
rect 128556 224862 128676 224890
rect 128556 222170 128584 224862
rect 128464 222142 128584 222170
rect 128464 215422 128492 222142
rect 128728 220108 128780 220114
rect 128728 220050 128780 220056
rect 128452 215416 128504 215422
rect 128452 215358 128504 215364
rect 128452 215280 128504 215286
rect 128452 215222 128504 215228
rect 128464 212537 128492 215222
rect 128450 212528 128506 212537
rect 128450 212463 128506 212472
rect 128634 212528 128690 212537
rect 128634 212463 128690 212472
rect 128648 202910 128676 212463
rect 128740 210458 128768 220050
rect 128728 210452 128780 210458
rect 128728 210394 128780 210400
rect 128452 202904 128504 202910
rect 128452 202846 128504 202852
rect 128636 202904 128688 202910
rect 128636 202846 128688 202852
rect 128464 198098 128492 202846
rect 128372 198070 128492 198098
rect 128372 195906 128400 198070
rect 128360 195900 128412 195906
rect 128360 195842 128412 195848
rect 128544 195900 128596 195906
rect 128544 195842 128596 195848
rect 128556 193225 128584 195842
rect 128728 195628 128780 195634
rect 128728 195570 128780 195576
rect 128358 193216 128414 193225
rect 128358 193151 128414 193160
rect 128542 193216 128598 193225
rect 128542 193151 128598 193160
rect 128372 183598 128400 193151
rect 128740 191146 128768 195570
rect 128728 191140 128780 191146
rect 128728 191082 128780 191088
rect 128360 183592 128412 183598
rect 128360 183534 128412 183540
rect 128544 183592 128596 183598
rect 128544 183534 128596 183540
rect 128556 176730 128584 183534
rect 128728 177404 128780 177410
rect 128728 177346 128780 177352
rect 128544 176724 128596 176730
rect 128544 176666 128596 176672
rect 128636 176588 128688 176594
rect 128636 176530 128688 176536
rect 128648 173890 128676 176530
rect 128740 175642 128768 177346
rect 128728 175636 128780 175642
rect 128728 175578 128780 175584
rect 128556 173862 128676 173890
rect 128556 169114 128584 173862
rect 128360 169108 128412 169114
rect 128360 169050 128412 169056
rect 128544 169108 128596 169114
rect 128544 169050 128596 169056
rect 128372 164257 128400 169050
rect 128358 164248 128414 164257
rect 128358 164183 128414 164192
rect 128542 164248 128598 164257
rect 128542 164183 128598 164192
rect 128556 154873 128584 164183
rect 128728 162172 128780 162178
rect 128728 162114 128780 162120
rect 128542 154864 128598 154873
rect 128542 154799 128598 154808
rect 128542 154592 128598 154601
rect 128542 154527 128598 154536
rect 128556 135266 128584 154527
rect 128740 149870 128768 162114
rect 128728 149864 128780 149870
rect 128728 149806 128780 149812
rect 128820 143540 128872 143546
rect 128820 143482 128872 143488
rect 128556 135250 128676 135266
rect 128832 135250 128860 143482
rect 128556 135244 128688 135250
rect 128556 135238 128636 135244
rect 128636 135186 128688 135192
rect 128728 135244 128780 135250
rect 128728 135186 128780 135192
rect 128820 135244 128872 135250
rect 128820 135186 128872 135192
rect 128648 135155 128676 135186
rect 128740 128382 128768 135186
rect 128820 130416 128872 130422
rect 128820 130358 128872 130364
rect 128728 128376 128780 128382
rect 128728 128318 128780 128324
rect 128636 128308 128688 128314
rect 128636 128250 128688 128256
rect 128648 125610 128676 128250
rect 128832 125633 128860 130358
rect 128818 125624 128874 125633
rect 128648 125594 128768 125610
rect 128648 125588 128780 125594
rect 128648 125582 128728 125588
rect 128818 125559 128820 125568
rect 128728 125530 128780 125536
rect 128872 125559 128874 125568
rect 128820 125530 128872 125536
rect 128268 118720 128320 118726
rect 128268 118662 128320 118668
rect 126980 118108 127032 118114
rect 126980 118050 127032 118056
rect 128176 118108 128228 118114
rect 128176 118050 128228 118056
rect 126888 117768 126940 117774
rect 126888 117710 126940 117716
rect 128188 117706 128216 118050
rect 127624 117700 127676 117706
rect 127624 117642 127676 117648
rect 128176 117700 128228 117706
rect 128176 117642 128228 117648
rect 126244 8492 126296 8498
rect 126244 8434 126296 8440
rect 126612 7404 126664 7410
rect 126612 7346 126664 7352
rect 125508 3052 125560 3058
rect 125508 2994 125560 3000
rect 126624 480 126652 7346
rect 127636 7342 127664 117642
rect 128832 117570 128860 125530
rect 128924 118318 128952 365638
rect 129016 143585 129044 552638
rect 129108 521626 129136 578546
rect 129280 578400 129332 578406
rect 129280 578342 129332 578348
rect 129188 553716 129240 553722
rect 129188 553658 129240 553664
rect 129096 521620 129148 521626
rect 129096 521562 129148 521568
rect 129200 496874 129228 553658
rect 129292 525094 129320 578342
rect 129464 563100 129516 563106
rect 129464 563042 129516 563048
rect 129280 525088 129332 525094
rect 129280 525030 129332 525036
rect 129372 500472 129424 500478
rect 129372 500414 129424 500420
rect 129188 496868 129240 496874
rect 129188 496810 129240 496816
rect 129094 387968 129150 387977
rect 129094 387903 129150 387912
rect 129108 374134 129136 387903
rect 129200 380633 129228 496810
rect 129186 380624 129242 380633
rect 129186 380559 129242 380568
rect 129096 374128 129148 374134
rect 129096 374070 129148 374076
rect 129096 360256 129148 360262
rect 129096 360198 129148 360204
rect 129108 347818 129136 360198
rect 129096 347812 129148 347818
rect 129096 347754 129148 347760
rect 129096 345568 129148 345574
rect 129096 345510 129148 345516
rect 129108 336054 129136 345510
rect 129096 336048 129148 336054
rect 129096 335990 129148 335996
rect 129096 327072 129148 327078
rect 129096 327014 129148 327020
rect 129108 311642 129136 327014
rect 129096 311636 129148 311642
rect 129096 311578 129148 311584
rect 129096 307080 129148 307086
rect 129096 307022 129148 307028
rect 129108 297430 129136 307022
rect 129096 297424 129148 297430
rect 129096 297366 129148 297372
rect 129096 287768 129148 287774
rect 129096 287710 129148 287716
rect 129108 274310 129136 287710
rect 129096 274304 129148 274310
rect 129096 274246 129148 274252
rect 129096 268456 129148 268462
rect 129096 268398 129148 268404
rect 129108 258806 129136 268398
rect 129096 258800 129148 258806
rect 129096 258742 129148 258748
rect 129096 249144 129148 249150
rect 129096 249086 129148 249092
rect 129108 239494 129136 249086
rect 129096 239488 129148 239494
rect 129096 239430 129148 239436
rect 129096 229764 129148 229770
rect 129096 229706 129148 229712
rect 129108 220114 129136 229706
rect 129096 220108 129148 220114
rect 129096 220050 129148 220056
rect 129096 210452 129148 210458
rect 129096 210394 129148 210400
rect 129108 195634 129136 210394
rect 129096 195628 129148 195634
rect 129096 195570 129148 195576
rect 129096 191140 129148 191146
rect 129096 191082 129148 191088
rect 129108 177410 129136 191082
rect 129096 177404 129148 177410
rect 129096 177346 129148 177352
rect 129096 175636 129148 175642
rect 129096 175578 129148 175584
rect 129108 162178 129136 175578
rect 129096 162172 129148 162178
rect 129096 162114 129148 162120
rect 129096 149864 129148 149870
rect 129096 149806 129148 149812
rect 129002 143576 129058 143585
rect 129108 143546 129136 149806
rect 129002 143511 129058 143520
rect 129096 143540 129148 143546
rect 129096 143482 129148 143488
rect 129096 135244 129148 135250
rect 129096 135186 129148 135192
rect 129108 130422 129136 135186
rect 129096 130416 129148 130422
rect 129096 130358 129148 130364
rect 129094 125624 129150 125633
rect 129200 125594 129228 380559
rect 129278 372736 129334 372745
rect 129278 372671 129334 372680
rect 129094 125559 129096 125568
rect 129148 125559 129150 125568
rect 129188 125588 129240 125594
rect 129096 125530 129148 125536
rect 129188 125530 129240 125536
rect 129096 125452 129148 125458
rect 129096 125394 129148 125400
rect 129188 125452 129240 125458
rect 129188 125394 129240 125400
rect 128912 118312 128964 118318
rect 128912 118254 128964 118260
rect 129108 117706 129136 125394
rect 129200 118153 129228 125394
rect 129292 118182 129320 372671
rect 129384 118794 129412 500414
rect 129476 118930 129504 563042
rect 129568 175166 129596 650014
rect 129660 175234 129688 696934
rect 130936 603152 130988 603158
rect 130936 603094 130988 603100
rect 130384 579012 130436 579018
rect 130384 578954 130436 578960
rect 129740 518900 129792 518906
rect 129740 518842 129792 518848
rect 129752 518566 129780 518842
rect 130396 518566 130424 578954
rect 129740 518560 129792 518566
rect 129740 518502 129792 518508
rect 130384 518560 130436 518566
rect 130384 518502 130436 518508
rect 129752 350985 129780 518502
rect 130844 500404 130896 500410
rect 130844 500346 130896 500352
rect 130660 500336 130712 500342
rect 130660 500278 130712 500284
rect 130568 462392 130620 462398
rect 130568 462334 130620 462340
rect 130108 397724 130160 397730
rect 130108 397666 130160 397672
rect 129738 350976 129794 350985
rect 129738 350911 129794 350920
rect 129752 350606 129780 350911
rect 129740 350600 129792 350606
rect 129740 350542 129792 350548
rect 130016 321632 130068 321638
rect 130016 321574 130068 321580
rect 129648 175228 129700 175234
rect 129648 175170 129700 175176
rect 129556 175160 129608 175166
rect 129556 175102 129608 175108
rect 130028 166870 130056 321574
rect 130120 202502 130148 397666
rect 130384 386368 130436 386374
rect 130384 386310 130436 386316
rect 130292 385008 130344 385014
rect 130292 384950 130344 384956
rect 130304 346526 130332 384950
rect 130292 346520 130344 346526
rect 130292 346462 130344 346468
rect 130200 340468 130252 340474
rect 130200 340410 130252 340416
rect 130108 202496 130160 202502
rect 130108 202438 130160 202444
rect 130016 166864 130068 166870
rect 130016 166806 130068 166812
rect 130212 119406 130240 340410
rect 130292 337544 130344 337550
rect 130292 337486 130344 337492
rect 130200 119400 130252 119406
rect 130200 119342 130252 119348
rect 129464 118924 129516 118930
rect 129464 118866 129516 118872
rect 129372 118788 129424 118794
rect 129372 118730 129424 118736
rect 129280 118176 129332 118182
rect 129186 118144 129242 118153
rect 129280 118118 129332 118124
rect 129186 118079 129242 118088
rect 129096 117700 129148 117706
rect 129096 117642 129148 117648
rect 128820 117564 128872 117570
rect 128820 117506 128872 117512
rect 128832 115977 128860 117506
rect 128818 115968 128874 115977
rect 128728 115932 128780 115938
rect 128818 115903 128874 115912
rect 129002 115968 129058 115977
rect 129002 115903 129004 115912
rect 128728 115874 128780 115880
rect 129056 115903 129058 115912
rect 129004 115874 129056 115880
rect 128740 106321 128768 115874
rect 128726 106312 128782 106321
rect 128726 106247 128782 106256
rect 128910 106312 128966 106321
rect 128910 106247 128966 106256
rect 128924 99090 128952 106247
rect 128924 99062 129136 99090
rect 129108 89706 129136 99062
rect 128924 89678 129136 89706
rect 128924 79914 128952 89678
rect 128924 79886 129044 79914
rect 129016 77246 129044 79886
rect 128912 77240 128964 77246
rect 128912 77182 128964 77188
rect 129004 77240 129056 77246
rect 129004 77182 129056 77188
rect 128924 67833 128952 77182
rect 128910 67824 128966 67833
rect 128910 67759 128966 67768
rect 129094 67688 129150 67697
rect 129094 67623 129150 67632
rect 129108 67590 129136 67623
rect 128820 67584 128872 67590
rect 128820 67526 128872 67532
rect 129096 67584 129148 67590
rect 129096 67526 129148 67532
rect 128832 60722 128860 67526
rect 128820 60716 128872 60722
rect 128820 60658 128872 60664
rect 129096 60716 129148 60722
rect 129096 60658 129148 60664
rect 129108 58018 129136 60658
rect 129016 57990 129136 58018
rect 129016 53258 129044 57990
rect 129016 53230 129136 53258
rect 129108 48346 129136 53230
rect 129096 48340 129148 48346
rect 129096 48282 129148 48288
rect 129004 48272 129056 48278
rect 129004 48214 129056 48220
rect 129016 47002 129044 48214
rect 129016 46974 129136 47002
rect 129108 46918 129136 46974
rect 129096 46912 129148 46918
rect 129096 46854 129148 46860
rect 129096 46776 129148 46782
rect 129096 46718 129148 46724
rect 129108 33862 129136 46718
rect 128820 33856 128872 33862
rect 128820 33798 128872 33804
rect 129096 33856 129148 33862
rect 129096 33798 129148 33804
rect 128832 31634 128860 33798
rect 128832 31606 128952 31634
rect 128924 22114 128952 31606
rect 128924 22086 129136 22114
rect 129108 19310 129136 22086
rect 128728 19304 128780 19310
rect 128728 19246 128780 19252
rect 129096 19304 129148 19310
rect 129096 19246 129148 19252
rect 128740 9722 128768 19246
rect 128728 9716 128780 9722
rect 128728 9658 128780 9664
rect 128912 9716 128964 9722
rect 128912 9658 128964 9664
rect 127624 7336 127676 7342
rect 127624 7278 127676 7284
rect 127808 7336 127860 7342
rect 127808 7278 127860 7284
rect 127820 480 127848 7278
rect 128924 7274 128952 9658
rect 129004 8832 129056 8838
rect 129004 8774 129056 8780
rect 128912 7268 128964 7274
rect 128912 7210 128964 7216
rect 128360 6248 128412 6254
rect 128360 6190 128412 6196
rect 128372 5574 128400 6190
rect 128360 5568 128412 5574
rect 128360 5510 128412 5516
rect 129016 480 129044 8774
rect 129200 8770 129228 118079
rect 129188 8764 129240 8770
rect 129188 8706 129240 8712
rect 129292 8702 129320 118118
rect 129372 117700 129424 117706
rect 129372 117642 129424 117648
rect 129280 8696 129332 8702
rect 129280 8638 129332 8644
rect 129384 8566 129412 117642
rect 130304 117230 130332 337486
rect 130396 118017 130424 386310
rect 130476 350600 130528 350606
rect 130476 350542 130528 350548
rect 130488 340678 130516 350542
rect 130476 340672 130528 340678
rect 130476 340614 130528 340620
rect 130382 118008 130438 118017
rect 130382 117943 130438 117952
rect 130488 117638 130516 340614
rect 130580 169833 130608 462334
rect 130672 172009 130700 500278
rect 130752 500268 130804 500274
rect 130752 500210 130804 500216
rect 130658 172000 130714 172009
rect 130658 171935 130714 171944
rect 130764 170921 130792 500210
rect 130750 170912 130806 170921
rect 130750 170847 130806 170856
rect 130566 169824 130622 169833
rect 130566 169759 130622 169768
rect 130856 119134 130884 500346
rect 130948 172961 130976 603094
rect 131028 583296 131080 583302
rect 131028 583238 131080 583244
rect 130934 172952 130990 172961
rect 130934 172887 130990 172896
rect 130934 156632 130990 156641
rect 130934 156567 130990 156576
rect 130948 148238 130976 156567
rect 130936 148232 130988 148238
rect 130936 148174 130988 148180
rect 130936 146396 130988 146402
rect 130936 146338 130988 146344
rect 130948 144378 130976 146338
rect 131040 144498 131068 583238
rect 131132 146402 131160 700674
rect 132040 700120 132092 700126
rect 132040 700062 132092 700068
rect 131948 638988 132000 638994
rect 131948 638930 132000 638936
rect 131856 498228 131908 498234
rect 131856 498170 131908 498176
rect 131764 310548 131816 310554
rect 131764 310490 131816 310496
rect 131580 274712 131632 274718
rect 131580 274654 131632 274660
rect 131304 200932 131356 200938
rect 131304 200874 131356 200880
rect 131210 199336 131266 199345
rect 131210 199271 131266 199280
rect 131224 198762 131252 199271
rect 131212 198756 131264 198762
rect 131212 198698 131264 198704
rect 131210 198248 131266 198257
rect 131210 198183 131266 198192
rect 131224 197402 131252 198183
rect 131212 197396 131264 197402
rect 131212 197338 131264 197344
rect 131316 197282 131344 200874
rect 131396 200864 131448 200870
rect 131396 200806 131448 200812
rect 131224 197254 131344 197282
rect 131224 196194 131252 197254
rect 131302 197160 131358 197169
rect 131302 197095 131358 197104
rect 131316 196382 131344 197095
rect 131304 196376 131356 196382
rect 131304 196318 131356 196324
rect 131224 196166 131344 196194
rect 131210 196072 131266 196081
rect 131210 196007 131212 196016
rect 131264 196007 131266 196016
rect 131212 195978 131264 195984
rect 131210 195120 131266 195129
rect 131210 195055 131266 195064
rect 131224 194614 131252 195055
rect 131212 194608 131264 194614
rect 131212 194550 131264 194556
rect 131212 194472 131264 194478
rect 131212 194414 131264 194420
rect 131224 194041 131252 194414
rect 131210 194032 131266 194041
rect 131210 193967 131266 193976
rect 131212 193112 131264 193118
rect 131212 193054 131264 193060
rect 131224 192953 131252 193054
rect 131210 192944 131266 192953
rect 131210 192879 131266 192888
rect 131212 192840 131264 192846
rect 131212 192782 131264 192788
rect 131224 192001 131252 192782
rect 131210 191992 131266 192001
rect 131210 191927 131266 191936
rect 131212 191820 131264 191826
rect 131212 191762 131264 191768
rect 131224 190913 131252 191762
rect 131210 190904 131266 190913
rect 131210 190839 131266 190848
rect 131212 190460 131264 190466
rect 131212 190402 131264 190408
rect 131224 189825 131252 190402
rect 131210 189816 131266 189825
rect 131210 189751 131266 189760
rect 131212 189032 131264 189038
rect 131212 188974 131264 188980
rect 131224 188737 131252 188974
rect 131210 188728 131266 188737
rect 131210 188663 131266 188672
rect 131212 188624 131264 188630
rect 131212 188566 131264 188572
rect 131224 187785 131252 188566
rect 131210 187776 131266 187785
rect 131210 187711 131266 187720
rect 131212 187672 131264 187678
rect 131212 187614 131264 187620
rect 131224 186697 131252 187614
rect 131210 186688 131266 186697
rect 131210 186623 131266 186632
rect 131212 186312 131264 186318
rect 131212 186254 131264 186260
rect 131224 185609 131252 186254
rect 131210 185600 131266 185609
rect 131210 185535 131266 185544
rect 131212 184884 131264 184890
rect 131212 184826 131264 184832
rect 131224 184521 131252 184826
rect 131210 184512 131266 184521
rect 131210 184447 131266 184456
rect 131210 183560 131266 183569
rect 131210 183495 131212 183504
rect 131264 183495 131266 183504
rect 131212 183466 131264 183472
rect 131212 175228 131264 175234
rect 131212 175170 131264 175176
rect 131224 175137 131252 175170
rect 131210 175128 131266 175137
rect 131210 175063 131266 175072
rect 131210 159352 131266 159361
rect 131210 159287 131266 159296
rect 131224 158778 131252 159287
rect 131212 158772 131264 158778
rect 131212 158714 131264 158720
rect 131210 156224 131266 156233
rect 131210 156159 131266 156168
rect 131224 155990 131252 156159
rect 131212 155984 131264 155990
rect 131212 155926 131264 155932
rect 131212 155848 131264 155854
rect 131212 155790 131264 155796
rect 131224 155145 131252 155790
rect 131210 155136 131266 155145
rect 131210 155071 131266 155080
rect 131212 154556 131264 154562
rect 131212 154498 131264 154504
rect 131224 154057 131252 154498
rect 131210 154048 131266 154057
rect 131210 153983 131266 153992
rect 131212 153196 131264 153202
rect 131212 153138 131264 153144
rect 131224 152969 131252 153138
rect 131210 152960 131266 152969
rect 131210 152895 131266 152904
rect 131212 152856 131264 152862
rect 131212 152798 131264 152804
rect 131224 152017 131252 152798
rect 131210 152008 131266 152017
rect 131210 151943 131266 151952
rect 131212 151768 131264 151774
rect 131212 151710 131264 151716
rect 131224 150929 131252 151710
rect 131210 150920 131266 150929
rect 131210 150855 131266 150864
rect 131212 150408 131264 150414
rect 131212 150350 131264 150356
rect 131224 149841 131252 150350
rect 131210 149832 131266 149841
rect 131210 149767 131266 149776
rect 131212 149048 131264 149054
rect 131212 148990 131264 148996
rect 131224 148753 131252 148990
rect 131210 148744 131266 148753
rect 131210 148679 131266 148688
rect 131212 148640 131264 148646
rect 131212 148582 131264 148588
rect 131224 148345 131252 148582
rect 131210 148336 131266 148345
rect 131210 148271 131266 148280
rect 131212 148232 131264 148238
rect 131212 148174 131264 148180
rect 131120 146396 131172 146402
rect 131120 146338 131172 146344
rect 131120 146260 131172 146266
rect 131120 146202 131172 146208
rect 131132 145625 131160 146202
rect 131118 145616 131174 145625
rect 131118 145551 131174 145560
rect 131120 144900 131172 144906
rect 131120 144842 131172 144848
rect 131132 144537 131160 144842
rect 131118 144528 131174 144537
rect 131028 144492 131080 144498
rect 131118 144463 131174 144472
rect 131028 144434 131080 144440
rect 130948 144350 131160 144378
rect 131028 144152 131080 144158
rect 131028 144094 131080 144100
rect 130844 119128 130896 119134
rect 130844 119070 130896 119076
rect 131040 118862 131068 144094
rect 131132 138281 131160 144350
rect 131118 138272 131174 138281
rect 131118 138207 131174 138216
rect 131028 118856 131080 118862
rect 131028 118798 131080 118804
rect 130476 117632 130528 117638
rect 130476 117574 130528 117580
rect 130292 117224 130344 117230
rect 130292 117166 130344 117172
rect 129372 8560 129424 8566
rect 129372 8502 129424 8508
rect 130200 7200 130252 7206
rect 130200 7142 130252 7148
rect 130212 480 130240 7142
rect 130488 4554 130516 117574
rect 131224 109002 131252 148174
rect 131316 132025 131344 196166
rect 131302 132016 131358 132025
rect 131302 131951 131358 131960
rect 131408 128761 131436 200806
rect 131488 200796 131540 200802
rect 131488 200738 131540 200744
rect 131394 128752 131450 128761
rect 131394 128687 131450 128696
rect 131500 127809 131528 200738
rect 131592 165617 131620 274654
rect 131672 263628 131724 263634
rect 131672 263570 131724 263576
rect 131578 165608 131634 165617
rect 131578 165543 131634 165552
rect 131578 158264 131634 158273
rect 131578 158199 131634 158208
rect 131486 127800 131542 127809
rect 131486 127735 131542 127744
rect 131212 108996 131264 109002
rect 131212 108938 131264 108944
rect 131592 64870 131620 158199
rect 131684 125633 131712 263570
rect 131776 126721 131804 310490
rect 131868 130937 131896 498170
rect 131960 134065 131988 638930
rect 132052 180441 132080 700062
rect 132132 685908 132184 685914
rect 132132 685850 132184 685856
rect 132038 180432 132094 180441
rect 132038 180367 132094 180376
rect 132040 175160 132092 175166
rect 132040 175102 132092 175108
rect 132052 174049 132080 175102
rect 132038 174040 132094 174049
rect 132038 173975 132094 173984
rect 132040 166864 132092 166870
rect 132040 166806 132092 166812
rect 132052 166705 132080 166806
rect 132038 166696 132094 166705
rect 132038 166631 132094 166640
rect 132038 160440 132094 160449
rect 132038 160375 132094 160384
rect 131946 134056 132002 134065
rect 131946 133991 132002 134000
rect 131854 130928 131910 130937
rect 131854 130863 131910 130872
rect 131762 126712 131818 126721
rect 131762 126647 131818 126656
rect 131670 125624 131726 125633
rect 131670 125559 131726 125568
rect 131580 64864 131632 64870
rect 131580 64806 131632 64812
rect 132052 41410 132080 160375
rect 132144 135153 132172 685850
rect 132236 147801 132264 700742
rect 132592 700392 132644 700398
rect 132592 700334 132644 700340
rect 132500 700324 132552 700330
rect 132500 700266 132552 700272
rect 132316 700188 132368 700194
rect 132316 700130 132368 700136
rect 132222 147792 132278 147801
rect 132222 147727 132278 147736
rect 132328 147626 132356 700130
rect 132408 318776 132460 318782
rect 132408 318718 132460 318724
rect 132420 309194 132448 318718
rect 132408 309188 132460 309194
rect 132408 309130 132460 309136
rect 132408 201000 132460 201006
rect 132408 200942 132460 200948
rect 132420 167793 132448 200942
rect 132406 167784 132462 167793
rect 132406 167719 132462 167728
rect 132406 162480 132462 162489
rect 132406 162415 132462 162424
rect 132224 147620 132276 147626
rect 132224 147562 132276 147568
rect 132316 147620 132368 147626
rect 132316 147562 132368 147568
rect 132236 146713 132264 147562
rect 132314 147520 132370 147529
rect 132314 147455 132370 147464
rect 132222 146704 132278 146713
rect 132222 146639 132278 146648
rect 132224 146600 132276 146606
rect 132224 146542 132276 146548
rect 132236 140457 132264 146542
rect 132328 142497 132356 147455
rect 132314 142488 132370 142497
rect 132314 142423 132370 142432
rect 132222 140448 132278 140457
rect 132222 140383 132278 140392
rect 132130 135144 132186 135153
rect 132130 135079 132186 135088
rect 132314 121408 132370 121417
rect 132314 121343 132370 121352
rect 132130 120456 132186 120465
rect 132130 120391 132186 120400
rect 132040 41404 132092 41410
rect 132040 41346 132092 41352
rect 132144 30326 132172 120391
rect 132328 77246 132356 121343
rect 132420 120698 132448 162415
rect 132512 136241 132540 700266
rect 132604 181286 132632 700334
rect 133144 700052 133196 700058
rect 133144 699994 133196 700000
rect 133052 699712 133104 699718
rect 133052 699654 133104 699660
rect 132960 415472 133012 415478
rect 132960 415414 133012 415420
rect 132776 346520 132828 346526
rect 132776 346462 132828 346468
rect 132788 340610 132816 346462
rect 132776 340604 132828 340610
rect 132776 340546 132828 340552
rect 132788 321586 132816 340546
rect 132696 321570 132816 321586
rect 132684 321564 132816 321570
rect 132736 321558 132816 321564
rect 132868 321564 132920 321570
rect 132684 321506 132736 321512
rect 132868 321506 132920 321512
rect 132696 321475 132724 321506
rect 132880 318782 132908 321506
rect 132868 318776 132920 318782
rect 132868 318718 132920 318724
rect 132776 309188 132828 309194
rect 132776 309130 132828 309136
rect 132788 302274 132816 309130
rect 132696 302246 132816 302274
rect 132696 302138 132724 302246
rect 132696 302110 132816 302138
rect 132788 292618 132816 302110
rect 132788 292590 132908 292618
rect 132880 282946 132908 292590
rect 132684 282940 132736 282946
rect 132684 282882 132736 282888
rect 132868 282940 132920 282946
rect 132868 282882 132920 282888
rect 132696 282826 132724 282882
rect 132696 282798 132816 282826
rect 132788 263650 132816 282798
rect 132696 263622 132816 263650
rect 132696 263514 132724 263622
rect 132696 263486 132816 263514
rect 132788 253994 132816 263486
rect 132788 253966 132908 253994
rect 132880 241505 132908 253966
rect 132866 241496 132922 241505
rect 132866 241431 132922 241440
rect 132684 227792 132736 227798
rect 132684 227734 132736 227740
rect 132592 181280 132644 181286
rect 132592 181222 132644 181228
rect 132696 164529 132724 227734
rect 132776 216708 132828 216714
rect 132776 216650 132828 216656
rect 132682 164520 132738 164529
rect 132682 164455 132738 164464
rect 132498 136232 132554 136241
rect 132498 136167 132554 136176
rect 132788 124545 132816 216650
rect 132868 210452 132920 210458
rect 132868 210394 132920 210400
rect 132880 196081 132908 210394
rect 132866 196072 132922 196081
rect 132866 196007 132922 196016
rect 132866 195936 132922 195945
rect 132866 195871 132922 195880
rect 132880 185230 132908 195871
rect 132868 185224 132920 185230
rect 132868 185166 132920 185172
rect 132868 185020 132920 185026
rect 132868 184962 132920 184968
rect 132880 182481 132908 184962
rect 132866 182472 132922 182481
rect 132866 182407 132922 182416
rect 132866 182336 132922 182345
rect 132866 182271 132922 182280
rect 132880 178265 132908 182271
rect 132866 178256 132922 178265
rect 132866 178191 132922 178200
rect 132972 168745 133000 415414
rect 133064 185026 133092 699654
rect 133156 185314 133184 699994
rect 133248 185473 133276 700810
rect 133420 700596 133472 700602
rect 133420 700538 133472 700544
rect 133328 700256 133380 700262
rect 133328 700198 133380 700204
rect 133234 185464 133290 185473
rect 133234 185399 133290 185408
rect 133156 185286 133276 185314
rect 133144 185224 133196 185230
rect 133144 185166 133196 185172
rect 133052 185020 133104 185026
rect 133052 184962 133104 184968
rect 133050 184920 133106 184929
rect 133050 184855 133106 184864
rect 132958 168736 133014 168745
rect 133064 168706 133092 184855
rect 132958 168671 133014 168680
rect 133052 168700 133104 168706
rect 133052 168642 133104 168648
rect 133052 168496 133104 168502
rect 133052 168438 133104 168444
rect 132958 164248 133014 164257
rect 132958 164183 133014 164192
rect 132972 154737 133000 164183
rect 132958 154728 133014 154737
rect 132958 154663 133014 154672
rect 132958 154592 133014 154601
rect 132880 154550 132958 154578
rect 132880 149682 132908 154550
rect 132958 154527 133014 154536
rect 132880 149654 133000 149682
rect 132972 144888 133000 149654
rect 132880 144860 133000 144888
rect 132880 135250 132908 144860
rect 132868 135244 132920 135250
rect 132868 135186 132920 135192
rect 132960 135176 133012 135182
rect 132960 135118 133012 135124
rect 132774 124536 132830 124545
rect 132774 124471 132830 124480
rect 132408 120692 132460 120698
rect 132408 120634 132460 120640
rect 132972 118561 133000 135118
rect 132958 118552 133014 118561
rect 132958 118487 133014 118496
rect 132972 117178 133000 118487
rect 133064 117609 133092 168438
rect 133156 164257 133184 185166
rect 133248 181393 133276 185286
rect 133234 181384 133290 181393
rect 133234 181319 133290 181328
rect 133236 181280 133288 181286
rect 133236 181222 133288 181228
rect 133248 176225 133276 181222
rect 133340 179353 133368 700198
rect 133326 179344 133382 179353
rect 133326 179279 133382 179288
rect 133432 177177 133460 700538
rect 133510 241496 133566 241505
rect 133510 241431 133566 241440
rect 133524 210458 133552 241431
rect 133512 210452 133564 210458
rect 133512 210394 133564 210400
rect 133512 200116 133564 200122
rect 133512 200058 133564 200064
rect 133524 189922 133552 200058
rect 133512 189916 133564 189922
rect 133512 189858 133564 189864
rect 133512 189780 133564 189786
rect 133512 189722 133564 189728
rect 133418 177168 133474 177177
rect 133418 177103 133474 177112
rect 133234 176216 133290 176225
rect 133234 176151 133290 176160
rect 133142 164248 133198 164257
rect 133142 164183 133198 164192
rect 133524 163577 133552 189722
rect 133510 163568 133566 163577
rect 133510 163503 133566 163512
rect 133510 161392 133566 161401
rect 133510 161327 133566 161336
rect 133234 118144 133290 118153
rect 133144 118108 133196 118114
rect 133234 118079 133236 118088
rect 133144 118050 133196 118056
rect 133288 118079 133290 118088
rect 133236 118050 133288 118056
rect 133050 117600 133106 117609
rect 133050 117535 133106 117544
rect 133156 117366 133184 118050
rect 133144 117360 133196 117366
rect 133144 117302 133196 117308
rect 132972 117150 133184 117178
rect 133156 99482 133184 117150
rect 133144 99476 133196 99482
rect 133144 99418 133196 99424
rect 133144 99340 133196 99346
rect 133144 99282 133196 99288
rect 133156 96642 133184 99282
rect 133156 96614 133276 96642
rect 132316 77240 132368 77246
rect 132316 77182 132368 77188
rect 133248 67658 133276 96614
rect 133524 88330 133552 161327
rect 133616 139369 133644 700878
rect 133696 700528 133748 700534
rect 133696 700470 133748 700476
rect 133602 139360 133658 139369
rect 133602 139295 133658 139304
rect 133708 137193 133736 700470
rect 133788 200184 133840 200190
rect 133788 200126 133840 200132
rect 133800 189786 133828 200126
rect 133788 189780 133840 189786
rect 133788 189722 133840 189728
rect 133788 189644 133840 189650
rect 133788 189586 133840 189592
rect 133694 137184 133750 137193
rect 133694 137119 133750 137128
rect 133800 117298 133828 189586
rect 133892 141409 133920 700946
rect 137848 699718 137876 703520
rect 154132 700806 154160 703520
rect 170324 700806 170352 703520
rect 154120 700800 154172 700806
rect 154120 700742 154172 700748
rect 170312 700800 170364 700806
rect 170312 700742 170364 700748
rect 202800 700058 202828 703520
rect 218992 701010 219020 703520
rect 235184 701010 235212 703520
rect 218980 701004 219032 701010
rect 218980 700946 219032 700952
rect 235172 701004 235224 701010
rect 235172 700946 235224 700952
rect 267660 700126 267688 703520
rect 283852 700194 283880 703520
rect 300136 700194 300164 703520
rect 332520 700262 332548 703520
rect 348804 700942 348832 703520
rect 364996 700942 365024 703520
rect 348792 700936 348844 700942
rect 348792 700878 348844 700884
rect 364984 700936 365036 700942
rect 364984 700878 365036 700884
rect 397472 700874 397500 703520
rect 397460 700868 397512 700874
rect 397460 700810 397512 700816
rect 413664 700738 413692 703520
rect 413652 700732 413704 700738
rect 413652 700674 413704 700680
rect 332508 700256 332560 700262
rect 332508 700198 332560 700204
rect 283840 700188 283892 700194
rect 283840 700130 283892 700136
rect 300124 700188 300176 700194
rect 300124 700130 300176 700136
rect 267648 700120 267700 700126
rect 267648 700062 267700 700068
rect 202788 700052 202840 700058
rect 202788 699994 202840 700000
rect 429856 699718 429884 703520
rect 434076 701004 434128 701010
rect 434076 700946 434128 700952
rect 433984 700936 434036 700942
rect 433984 700878 434036 700884
rect 137836 699712 137888 699718
rect 137836 699654 137888 699660
rect 429844 699712 429896 699718
rect 429844 699654 429896 699660
rect 433892 699712 433944 699718
rect 433892 699654 433944 699660
rect 133972 592068 134024 592074
rect 133972 592010 134024 592016
rect 133878 141400 133934 141409
rect 133878 141335 133934 141344
rect 133984 133521 134012 592010
rect 302792 583704 302844 583710
rect 302792 583646 302844 583652
rect 270408 583636 270460 583642
rect 270408 583578 270460 583584
rect 199384 583500 199436 583506
rect 199384 583442 199436 583448
rect 157340 579080 157392 579086
rect 157340 579022 157392 579028
rect 162400 579080 162452 579086
rect 162400 579022 162452 579028
rect 176660 579080 176712 579086
rect 176660 579022 176712 579028
rect 181720 579080 181772 579086
rect 181720 579022 181772 579028
rect 195980 579080 196032 579086
rect 195980 579022 196032 579028
rect 152556 579012 152608 579018
rect 152556 578954 152608 578960
rect 137836 578944 137888 578950
rect 137836 578886 137888 578892
rect 147588 578944 147640 578950
rect 147588 578886 147640 578892
rect 152280 578944 152332 578950
rect 152280 578886 152332 578892
rect 152372 578944 152424 578950
rect 152372 578886 152424 578892
rect 137848 578490 137876 578886
rect 138664 578808 138716 578814
rect 138664 578750 138716 578756
rect 138112 578672 138164 578678
rect 138112 578614 138164 578620
rect 137928 578536 137980 578542
rect 137848 578484 137928 578490
rect 137848 578478 137980 578484
rect 138020 578536 138072 578542
rect 138124 578524 138152 578614
rect 138072 578496 138152 578524
rect 138020 578478 138072 578484
rect 137848 578462 137968 578478
rect 138676 578474 138704 578750
rect 147600 578746 147628 578886
rect 147588 578740 147640 578746
rect 147588 578682 147640 578688
rect 152292 578678 152320 578886
rect 139584 578672 139636 578678
rect 139584 578614 139636 578620
rect 152280 578672 152332 578678
rect 152280 578614 152332 578620
rect 139596 578474 139624 578614
rect 152384 578474 152412 578886
rect 152568 578814 152596 578954
rect 157248 578944 157300 578950
rect 157248 578886 157300 578892
rect 152464 578808 152516 578814
rect 152464 578750 152516 578756
rect 152556 578808 152608 578814
rect 152556 578750 152608 578756
rect 152476 578474 152504 578750
rect 157260 578542 157288 578886
rect 157352 578542 157380 579022
rect 162308 578808 162360 578814
rect 162308 578750 162360 578756
rect 157248 578536 157300 578542
rect 157248 578478 157300 578484
rect 157340 578536 157392 578542
rect 157340 578478 157392 578484
rect 162320 578474 162348 578750
rect 162412 578474 162440 579022
rect 171876 579012 171928 579018
rect 171876 578954 171928 578960
rect 171600 578944 171652 578950
rect 171600 578886 171652 578892
rect 171692 578944 171744 578950
rect 171692 578886 171744 578892
rect 171612 578678 171640 578886
rect 171600 578672 171652 578678
rect 171600 578614 171652 578620
rect 171704 578474 171732 578886
rect 171888 578814 171916 578954
rect 176568 578944 176620 578950
rect 176568 578886 176620 578892
rect 171784 578808 171836 578814
rect 171784 578750 171836 578756
rect 171876 578808 171928 578814
rect 171876 578750 171928 578756
rect 171796 578474 171824 578750
rect 176580 578542 176608 578886
rect 176672 578542 176700 579022
rect 181628 578808 181680 578814
rect 181628 578750 181680 578756
rect 176568 578536 176620 578542
rect 176568 578478 176620 578484
rect 176660 578536 176712 578542
rect 176660 578478 176712 578484
rect 181640 578474 181668 578750
rect 181732 578474 181760 579022
rect 191196 579012 191248 579018
rect 191196 578954 191248 578960
rect 190920 578944 190972 578950
rect 190920 578886 190972 578892
rect 191012 578944 191064 578950
rect 191012 578886 191064 578892
rect 190932 578678 190960 578886
rect 190920 578672 190972 578678
rect 190920 578614 190972 578620
rect 191024 578474 191052 578886
rect 191208 578814 191236 578954
rect 195888 578944 195940 578950
rect 195888 578886 195940 578892
rect 191104 578808 191156 578814
rect 191104 578750 191156 578756
rect 191196 578808 191248 578814
rect 191196 578750 191248 578756
rect 191116 578474 191144 578750
rect 195900 578542 195928 578886
rect 195992 578542 196020 579022
rect 195888 578536 195940 578542
rect 195888 578478 195940 578484
rect 195980 578536 196032 578542
rect 195980 578478 196032 578484
rect 138664 578468 138716 578474
rect 138664 578410 138716 578416
rect 139584 578468 139636 578474
rect 139584 578410 139636 578416
rect 152372 578468 152424 578474
rect 152372 578410 152424 578416
rect 152464 578468 152516 578474
rect 152464 578410 152516 578416
rect 162308 578468 162360 578474
rect 162308 578410 162360 578416
rect 162400 578468 162452 578474
rect 162400 578410 162452 578416
rect 171692 578468 171744 578474
rect 171692 578410 171744 578416
rect 171784 578468 171836 578474
rect 171784 578410 171836 578416
rect 181628 578468 181680 578474
rect 181628 578410 181680 578416
rect 181720 578468 181772 578474
rect 181720 578410 181772 578416
rect 191012 578468 191064 578474
rect 191012 578410 191064 578416
rect 191104 578468 191156 578474
rect 191104 578410 191156 578416
rect 195796 562080 195848 562086
rect 195796 562022 195848 562028
rect 195704 562012 195756 562018
rect 195704 561954 195756 561960
rect 156604 553920 156656 553926
rect 156604 553862 156656 553868
rect 137284 553648 137336 553654
rect 137284 553590 137336 553596
rect 134064 451308 134116 451314
rect 134064 451250 134116 451256
rect 133970 133512 134026 133521
rect 133970 133447 134026 133456
rect 134076 130393 134104 451250
rect 135260 342916 135312 342922
rect 135260 342858 135312 342864
rect 135272 342514 135300 342858
rect 135260 342508 135312 342514
rect 135260 342450 135312 342456
rect 134338 341456 134394 341465
rect 134338 341391 134394 341400
rect 134156 201612 134208 201618
rect 134156 201554 134208 201560
rect 134168 200002 134196 201554
rect 134352 200161 134380 341391
rect 134432 202496 134484 202502
rect 134432 202438 134484 202444
rect 134338 200152 134394 200161
rect 134338 200087 134394 200096
rect 134444 200002 134472 202438
rect 134708 202156 134760 202162
rect 134708 202098 134760 202104
rect 134720 200002 134748 202098
rect 135272 200122 135300 342450
rect 137296 202366 137324 553590
rect 141424 553580 141476 553586
rect 141424 553522 141476 553528
rect 140044 536852 140096 536858
rect 140044 536794 140096 536800
rect 138020 398268 138072 398274
rect 138020 398210 138072 398216
rect 138032 340474 138060 398210
rect 138020 340468 138072 340474
rect 138020 340410 138072 340416
rect 137284 202360 137336 202366
rect 137284 202302 137336 202308
rect 140056 202298 140084 536794
rect 140044 202292 140096 202298
rect 140044 202234 140096 202240
rect 141436 202162 141464 553522
rect 151084 553512 151136 553518
rect 151084 553454 151136 553460
rect 144184 518356 144236 518362
rect 144184 518298 144236 518304
rect 144196 202230 144224 518298
rect 151096 202434 151124 553454
rect 155224 542428 155276 542434
rect 155224 542370 155276 542376
rect 153844 532772 153896 532778
rect 153844 532714 153896 532720
rect 152464 518288 152516 518294
rect 152464 518230 152516 518236
rect 152476 202502 152504 518230
rect 153856 202570 153884 532714
rect 155236 497826 155264 542370
rect 155224 497820 155276 497826
rect 155224 497762 155276 497768
rect 155236 496942 155264 497762
rect 155224 496936 155276 496942
rect 155224 496878 155276 496884
rect 155868 496936 155920 496942
rect 155868 496878 155920 496884
rect 155880 407658 155908 496878
rect 155224 407652 155276 407658
rect 155224 407594 155276 407600
rect 155868 407652 155920 407658
rect 155868 407594 155920 407600
rect 155236 398138 155264 407594
rect 155880 407250 155908 407594
rect 155868 407244 155920 407250
rect 155868 407186 155920 407192
rect 155224 398132 155276 398138
rect 155224 398074 155276 398080
rect 154578 340504 154634 340513
rect 154578 340439 154580 340448
rect 154632 340439 154634 340448
rect 154580 340410 154632 340416
rect 156616 202638 156644 553862
rect 195060 520940 195112 520946
rect 195060 520882 195112 520888
rect 191104 506524 191156 506530
rect 191104 506466 191156 506472
rect 188344 407856 188396 407862
rect 188344 407798 188396 407804
rect 168656 395616 168708 395622
rect 168656 395558 168708 395564
rect 157338 340504 157394 340513
rect 157338 340439 157394 340448
rect 157352 340406 157380 340439
rect 157340 340400 157392 340406
rect 157340 340342 157392 340348
rect 156604 202632 156656 202638
rect 156604 202574 156656 202580
rect 153844 202564 153896 202570
rect 153844 202506 153896 202512
rect 152464 202496 152516 202502
rect 152464 202438 152516 202444
rect 151084 202428 151136 202434
rect 151084 202370 151136 202376
rect 168380 202360 168432 202366
rect 168380 202302 168432 202308
rect 142528 202224 142580 202230
rect 142528 202166 142580 202172
rect 144184 202224 144236 202230
rect 144184 202166 144236 202172
rect 141424 202156 141476 202162
rect 141424 202098 141476 202104
rect 135260 200116 135312 200122
rect 135260 200058 135312 200064
rect 142540 200002 142568 202166
rect 168392 200002 168420 202302
rect 168668 200002 168696 395558
rect 179512 395548 179564 395554
rect 179512 395490 179564 395496
rect 173912 340598 174032 340626
rect 173912 340542 173940 340598
rect 173900 340536 173952 340542
rect 173900 340478 173952 340484
rect 174004 340338 174032 340598
rect 173992 340332 174044 340338
rect 173992 340274 174044 340280
rect 169116 202632 169168 202638
rect 169116 202574 169168 202580
rect 169128 200002 169156 202574
rect 178040 202564 178092 202570
rect 178040 202506 178092 202512
rect 176936 202496 176988 202502
rect 176936 202438 176988 202444
rect 176948 200002 176976 202438
rect 178052 200002 178080 202506
rect 178684 202292 178736 202298
rect 178684 202234 178736 202240
rect 178696 200002 178724 202234
rect 179524 200002 179552 395490
rect 188356 356046 188384 407798
rect 185584 356040 185636 356046
rect 185584 355982 185636 355988
rect 188344 356040 188396 356046
rect 188344 355982 188396 355988
rect 185596 341465 185624 355982
rect 191116 342922 191144 506466
rect 191104 342916 191156 342922
rect 191104 342858 191156 342864
rect 185582 341456 185638 341465
rect 185582 341391 185638 341400
rect 183468 340468 183520 340474
rect 183468 340410 183520 340416
rect 183480 340338 183508 340410
rect 193220 340400 193272 340406
rect 193218 340368 193220 340377
rect 193272 340368 193274 340377
rect 183468 340332 183520 340338
rect 193218 340303 193274 340312
rect 183468 340274 183520 340280
rect 195072 338774 195100 520882
rect 195520 410100 195572 410106
rect 195520 410042 195572 410048
rect 195428 409556 195480 409562
rect 195428 409498 195480 409504
rect 195152 409488 195204 409494
rect 195152 409430 195204 409436
rect 195060 338768 195112 338774
rect 195060 338710 195112 338716
rect 195164 205086 195192 409430
rect 195336 409284 195388 409290
rect 195336 409226 195388 409232
rect 195244 409148 195296 409154
rect 195244 409090 195296 409096
rect 195152 205080 195204 205086
rect 195152 205022 195204 205028
rect 195256 205018 195284 409090
rect 195244 205012 195296 205018
rect 195244 204954 195296 204960
rect 195348 202774 195376 409226
rect 195336 202768 195388 202774
rect 195336 202710 195388 202716
rect 182180 202428 182232 202434
rect 182180 202370 182232 202376
rect 181260 202224 181312 202230
rect 181260 202166 181312 202172
rect 180340 202156 180392 202162
rect 180340 202098 180392 202104
rect 180352 200002 180380 202098
rect 181272 200002 181300 202166
rect 182192 200002 182220 202370
rect 195440 202026 195468 409498
rect 195532 202502 195560 410042
rect 195612 410032 195664 410038
rect 195612 409974 195664 409980
rect 195520 202496 195572 202502
rect 195520 202438 195572 202444
rect 195624 202366 195652 409974
rect 195716 202745 195744 561954
rect 195702 202736 195758 202745
rect 195702 202671 195758 202680
rect 195808 202609 195836 562022
rect 197268 561944 197320 561950
rect 197268 561886 197320 561892
rect 195888 561876 195940 561882
rect 195888 561818 195940 561824
rect 195794 202600 195850 202609
rect 195794 202535 195850 202544
rect 195612 202360 195664 202366
rect 195612 202302 195664 202308
rect 195428 202020 195480 202026
rect 195428 201962 195480 201968
rect 195900 201958 195928 561818
rect 197176 561808 197228 561814
rect 197176 561750 197228 561756
rect 197084 560244 197136 560250
rect 197084 560186 197136 560192
rect 196440 521008 196492 521014
rect 196440 520950 196492 520956
rect 196348 518288 196400 518294
rect 196348 518230 196400 518236
rect 196360 339046 196388 518230
rect 196348 339040 196400 339046
rect 196348 338982 196400 338988
rect 196452 338842 196480 520950
rect 196992 409896 197044 409902
rect 196992 409838 197044 409844
rect 196808 409692 196860 409698
rect 196808 409634 196860 409640
rect 196624 409420 196676 409426
rect 196624 409362 196676 409368
rect 196532 409216 196584 409222
rect 196532 409158 196584 409164
rect 196440 338836 196492 338842
rect 196440 338778 196492 338784
rect 196544 204950 196572 409158
rect 196636 205154 196664 409362
rect 196716 409352 196768 409358
rect 196716 409294 196768 409300
rect 196624 205148 196676 205154
rect 196624 205090 196676 205096
rect 196532 204944 196584 204950
rect 196532 204886 196584 204892
rect 196728 202842 196756 409294
rect 196716 202836 196768 202842
rect 196716 202778 196768 202784
rect 195888 201952 195940 201958
rect 195888 201894 195940 201900
rect 196820 201822 196848 409634
rect 196900 409624 196952 409630
rect 196900 409566 196952 409572
rect 196912 202094 196940 409566
rect 197004 202570 197032 409838
rect 196992 202564 197044 202570
rect 196992 202506 197044 202512
rect 197096 202337 197124 560186
rect 197188 202473 197216 561750
rect 197280 202881 197308 561886
rect 198646 556744 198702 556753
rect 198646 556679 198702 556688
rect 198554 552120 198610 552129
rect 198554 552055 198610 552064
rect 198462 543824 198518 543833
rect 198462 543759 198518 543768
rect 198370 538520 198426 538529
rect 198370 538455 198426 538464
rect 198278 524648 198334 524657
rect 198278 524583 198334 524592
rect 197728 406564 197780 406570
rect 197728 406506 197780 406512
rect 197740 365702 197768 406506
rect 198186 399664 198242 399673
rect 198186 399599 198242 399608
rect 198094 391232 198150 391241
rect 198094 391167 198150 391176
rect 198002 387152 198058 387161
rect 198002 387087 198058 387096
rect 197910 378720 197966 378729
rect 197910 378655 197966 378664
rect 197818 370288 197874 370297
rect 197818 370223 197874 370232
rect 197728 365696 197780 365702
rect 197728 365638 197780 365644
rect 197726 361856 197782 361865
rect 197726 361791 197782 361800
rect 197634 357504 197690 357513
rect 197634 357439 197690 357448
rect 197542 353424 197598 353433
rect 197542 353359 197598 353368
rect 197450 349072 197506 349081
rect 197450 349007 197506 349016
rect 197464 204134 197492 349007
rect 197452 204128 197504 204134
rect 197452 204070 197504 204076
rect 197556 203726 197584 353359
rect 197648 204202 197676 357439
rect 197636 204196 197688 204202
rect 197636 204138 197688 204144
rect 197740 203930 197768 361791
rect 197728 203924 197780 203930
rect 197728 203866 197780 203872
rect 197544 203720 197596 203726
rect 197544 203662 197596 203668
rect 197832 203658 197860 370223
rect 197924 203862 197952 378655
rect 197912 203856 197964 203862
rect 197912 203798 197964 203804
rect 197820 203652 197872 203658
rect 197820 203594 197872 203600
rect 198016 203590 198044 387087
rect 198004 203584 198056 203590
rect 198004 203526 198056 203532
rect 198108 203522 198136 391167
rect 198200 203794 198228 399599
rect 198188 203788 198240 203794
rect 198188 203730 198240 203736
rect 198096 203516 198148 203522
rect 198096 203458 198148 203464
rect 197266 202872 197322 202881
rect 197266 202807 197322 202816
rect 198292 202638 198320 524583
rect 198384 203386 198412 538455
rect 198372 203380 198424 203386
rect 198372 203322 198424 203328
rect 198280 202632 198332 202638
rect 198280 202574 198332 202580
rect 197174 202464 197230 202473
rect 197174 202399 197230 202408
rect 197082 202328 197138 202337
rect 197082 202263 197138 202272
rect 196900 202088 196952 202094
rect 196900 202030 196952 202036
rect 196808 201816 196860 201822
rect 196808 201758 196860 201764
rect 198476 201618 198504 543759
rect 198568 201686 198596 552055
rect 198660 202065 198688 556679
rect 199396 549914 199424 583442
rect 201040 579080 201092 579086
rect 201040 579022 201092 579028
rect 215300 579080 215352 579086
rect 215300 579022 215352 579028
rect 220360 579080 220412 579086
rect 220360 579022 220412 579028
rect 234620 579080 234672 579086
rect 234620 579022 234672 579028
rect 239680 579080 239732 579086
rect 239680 579022 239732 579028
rect 253940 579080 253992 579086
rect 253940 579022 253992 579028
rect 259000 579080 259052 579086
rect 259000 579022 259052 579028
rect 200948 578808 201000 578814
rect 200948 578750 201000 578756
rect 200960 578474 200988 578750
rect 201052 578474 201080 579022
rect 210516 579012 210568 579018
rect 210516 578954 210568 578960
rect 210240 578944 210292 578950
rect 210240 578886 210292 578892
rect 210332 578944 210384 578950
rect 210332 578886 210384 578892
rect 210252 578678 210280 578886
rect 210240 578672 210292 578678
rect 210240 578614 210292 578620
rect 210344 578474 210372 578886
rect 210528 578814 210556 578954
rect 215208 578944 215260 578950
rect 215208 578886 215260 578892
rect 210424 578808 210476 578814
rect 210424 578750 210476 578756
rect 210516 578808 210568 578814
rect 210516 578750 210568 578756
rect 210436 578474 210464 578750
rect 215220 578542 215248 578886
rect 215312 578542 215340 579022
rect 220268 578808 220320 578814
rect 220268 578750 220320 578756
rect 215208 578536 215260 578542
rect 215208 578478 215260 578484
rect 215300 578536 215352 578542
rect 215300 578478 215352 578484
rect 220280 578474 220308 578750
rect 220372 578474 220400 579022
rect 229836 579012 229888 579018
rect 229836 578954 229888 578960
rect 229560 578944 229612 578950
rect 229560 578886 229612 578892
rect 229652 578944 229704 578950
rect 229652 578886 229704 578892
rect 229572 578678 229600 578886
rect 229560 578672 229612 578678
rect 229560 578614 229612 578620
rect 229664 578474 229692 578886
rect 229848 578814 229876 578954
rect 234528 578944 234580 578950
rect 234528 578886 234580 578892
rect 229744 578808 229796 578814
rect 229744 578750 229796 578756
rect 229836 578808 229888 578814
rect 229836 578750 229888 578756
rect 229756 578474 229784 578750
rect 234540 578542 234568 578886
rect 234632 578542 234660 579022
rect 239588 578808 239640 578814
rect 239588 578750 239640 578756
rect 234528 578536 234580 578542
rect 234528 578478 234580 578484
rect 234620 578536 234672 578542
rect 234620 578478 234672 578484
rect 239600 578474 239628 578750
rect 239692 578474 239720 579022
rect 249156 579012 249208 579018
rect 249156 578954 249208 578960
rect 248880 578944 248932 578950
rect 248880 578886 248932 578892
rect 248972 578944 249024 578950
rect 248972 578886 249024 578892
rect 248892 578678 248920 578886
rect 248880 578672 248932 578678
rect 248880 578614 248932 578620
rect 248984 578474 249012 578886
rect 249168 578814 249196 578954
rect 253848 578944 253900 578950
rect 253848 578886 253900 578892
rect 249064 578808 249116 578814
rect 249064 578750 249116 578756
rect 249156 578808 249208 578814
rect 249156 578750 249208 578756
rect 249076 578474 249104 578750
rect 253860 578542 253888 578886
rect 253952 578542 253980 579022
rect 258908 578808 258960 578814
rect 258908 578750 258960 578756
rect 253848 578536 253900 578542
rect 253848 578478 253900 578484
rect 253940 578536 253992 578542
rect 253940 578478 253992 578484
rect 258920 578474 258948 578750
rect 259012 578474 259040 579022
rect 268476 579012 268528 579018
rect 268476 578954 268528 578960
rect 268108 578944 268160 578950
rect 268108 578886 268160 578892
rect 268292 578944 268344 578950
rect 268292 578886 268344 578892
rect 268120 578678 268148 578886
rect 268108 578672 268160 578678
rect 268108 578614 268160 578620
rect 268304 578474 268332 578886
rect 268488 578814 268516 578954
rect 268384 578808 268436 578814
rect 268384 578750 268436 578756
rect 268476 578808 268528 578814
rect 268476 578750 268528 578756
rect 268396 578474 268424 578750
rect 200948 578468 201000 578474
rect 200948 578410 201000 578416
rect 201040 578468 201092 578474
rect 201040 578410 201092 578416
rect 210332 578468 210384 578474
rect 210332 578410 210384 578416
rect 210424 578468 210476 578474
rect 210424 578410 210476 578416
rect 220268 578468 220320 578474
rect 220268 578410 220320 578416
rect 220360 578468 220412 578474
rect 220360 578410 220412 578416
rect 229652 578468 229704 578474
rect 229652 578410 229704 578416
rect 229744 578468 229796 578474
rect 229744 578410 229796 578416
rect 239588 578468 239640 578474
rect 239588 578410 239640 578416
rect 239680 578468 239732 578474
rect 239680 578410 239732 578416
rect 248972 578468 249024 578474
rect 248972 578410 249024 578416
rect 249064 578468 249116 578474
rect 249064 578410 249116 578416
rect 258908 578468 258960 578474
rect 258908 578410 258960 578416
rect 259000 578468 259052 578474
rect 259000 578410 259052 578416
rect 268292 578468 268344 578474
rect 268292 578410 268344 578416
rect 268384 578468 268436 578474
rect 268384 578410 268436 578416
rect 200120 562148 200172 562154
rect 200120 562090 200172 562096
rect 209688 562148 209740 562154
rect 209688 562090 209740 562096
rect 200132 561814 200160 562090
rect 205548 562012 205600 562018
rect 205548 561954 205600 561960
rect 200120 561808 200172 561814
rect 200120 561750 200172 561756
rect 202052 560244 202104 560250
rect 202052 560186 202104 560192
rect 202064 559994 202092 560186
rect 202064 559966 202446 559994
rect 205560 559980 205588 561954
rect 208676 561944 208728 561950
rect 208676 561886 208728 561892
rect 208688 559980 208716 561886
rect 209700 561746 209728 562090
rect 214748 562080 214800 562086
rect 214748 562022 214800 562028
rect 211620 561876 211672 561882
rect 211620 561818 211672 561824
rect 209688 561740 209740 561746
rect 209688 561682 209740 561688
rect 211632 559980 211660 561818
rect 214760 559980 214788 562022
rect 217876 561740 217928 561746
rect 217876 561682 217928 561688
rect 217888 559980 217916 561682
rect 222198 556200 222254 556209
rect 222198 556135 222254 556144
rect 199384 549908 199436 549914
rect 199384 549850 199436 549856
rect 198922 547904 198978 547913
rect 198922 547839 198978 547848
rect 198738 534168 198794 534177
rect 198738 534103 198794 534112
rect 198646 202056 198702 202065
rect 198646 201991 198702 202000
rect 198752 201754 198780 534103
rect 198830 529272 198886 529281
rect 198830 529207 198886 529216
rect 198740 201748 198792 201754
rect 198740 201690 198792 201696
rect 198556 201680 198608 201686
rect 198556 201622 198608 201628
rect 198464 201612 198516 201618
rect 198464 201554 198516 201560
rect 198844 201550 198872 529207
rect 198936 291854 198964 547839
rect 219438 529000 219494 529009
rect 219438 528935 219494 528944
rect 199752 521144 199804 521150
rect 199752 521086 199804 521092
rect 199384 406496 199436 406502
rect 199384 406438 199436 406444
rect 199014 403744 199070 403753
rect 199014 403679 199070 403688
rect 198924 291848 198976 291854
rect 198924 291790 198976 291796
rect 199028 202201 199056 403679
rect 199106 395312 199162 395321
rect 199106 395247 199162 395256
rect 199120 202230 199148 395247
rect 199396 391950 199424 406438
rect 199384 391944 199436 391950
rect 199384 391886 199436 391892
rect 199198 382800 199254 382809
rect 199198 382735 199254 382744
rect 199212 203998 199240 382735
rect 199290 374368 199346 374377
rect 199290 374303 199346 374312
rect 199200 203992 199252 203998
rect 199200 203934 199252 203940
rect 199108 202224 199160 202230
rect 199014 202192 199070 202201
rect 199108 202166 199160 202172
rect 199304 202162 199332 374303
rect 199382 365936 199438 365945
rect 199382 365871 199438 365880
rect 199396 204066 199424 365871
rect 199474 344992 199530 345001
rect 199474 344927 199530 344936
rect 199488 204270 199516 344927
rect 199660 342780 199712 342786
rect 199660 342722 199712 342728
rect 199476 204264 199528 204270
rect 199476 204206 199528 204212
rect 199384 204060 199436 204066
rect 199384 204002 199436 204008
rect 199014 202127 199070 202136
rect 199292 202156 199344 202162
rect 199292 202098 199344 202104
rect 199672 201890 199700 342722
rect 199764 338978 199792 521086
rect 199844 521076 199896 521082
rect 199844 521018 199896 521024
rect 199752 338972 199804 338978
rect 199752 338914 199804 338920
rect 199856 338910 199884 521018
rect 200224 520118 200606 520146
rect 202892 520118 203550 520146
rect 200028 410168 200080 410174
rect 200028 410110 200080 410116
rect 199936 409964 199988 409970
rect 199936 409906 199988 409912
rect 199844 338904 199896 338910
rect 199844 338846 199896 338852
rect 199948 202434 199976 409906
rect 200040 202706 200068 410110
rect 200224 342786 200252 520118
rect 200580 409896 200632 409902
rect 200580 409838 200632 409844
rect 200592 408748 200620 409838
rect 202892 409698 202920 520118
rect 206664 517546 206692 520132
rect 205640 517540 205692 517546
rect 205640 517482 205692 517488
rect 206652 517540 206704 517546
rect 206652 517482 206704 517488
rect 203340 410576 203392 410582
rect 203340 410518 203392 410524
rect 202880 409692 202932 409698
rect 202880 409634 202932 409640
rect 203352 408748 203380 410518
rect 205652 409630 205680 517482
rect 206284 410644 206336 410650
rect 206284 410586 206336 410592
rect 205640 409624 205692 409630
rect 205640 409566 205692 409572
rect 206296 408748 206324 410586
rect 209044 409964 209096 409970
rect 209044 409906 209096 409912
rect 209056 408748 209084 409906
rect 209792 409562 209820 520132
rect 212552 520118 212934 520146
rect 215312 520118 216062 520146
rect 211988 410712 212040 410718
rect 211988 410654 212040 410660
rect 209780 409556 209832 409562
rect 209780 409498 209832 409504
rect 212000 408748 212028 410654
rect 212552 409494 212580 520118
rect 214748 410032 214800 410038
rect 214748 409974 214800 409980
rect 212540 409488 212592 409494
rect 212540 409430 212592 409436
rect 214760 408748 214788 409974
rect 215312 409426 215340 520118
rect 218992 518294 219020 520132
rect 218980 518288 219032 518294
rect 218980 518230 219032 518236
rect 217692 410168 217744 410174
rect 217692 410110 217744 410116
rect 215300 409420 215352 409426
rect 215300 409362 215352 409368
rect 217704 408748 217732 410110
rect 219452 409358 219480 528935
rect 219530 524512 219586 524521
rect 219530 524447 219586 524456
rect 219440 409352 219492 409358
rect 219440 409294 219492 409300
rect 219544 409290 219572 524447
rect 220452 410100 220504 410106
rect 220452 410042 220504 410048
rect 219532 409284 219584 409290
rect 219532 409226 219584 409232
rect 220464 408748 220492 410042
rect 222212 409222 222240 556135
rect 222290 552120 222346 552129
rect 222290 552055 222346 552064
rect 222200 409216 222252 409222
rect 222200 409158 222252 409164
rect 222304 409154 222332 552055
rect 222382 546952 222438 546961
rect 222382 546887 222438 546896
rect 222396 521150 222424 546887
rect 222474 542600 222530 542609
rect 222474 542535 222530 542544
rect 222384 521144 222436 521150
rect 222384 521086 222436 521092
rect 222488 521014 222516 542535
rect 222566 538384 222622 538393
rect 222566 538319 222622 538328
rect 222580 521082 222608 538319
rect 222658 533352 222714 533361
rect 222658 533287 222714 533296
rect 222568 521076 222620 521082
rect 222568 521018 222620 521024
rect 222476 521008 222528 521014
rect 222476 520950 222528 520956
rect 222672 520946 222700 533287
rect 222660 520940 222712 520946
rect 222660 520882 222712 520888
rect 261300 451376 261352 451382
rect 261300 451318 261352 451324
rect 261312 447098 261340 451318
rect 261300 447092 261352 447098
rect 261300 447034 261352 447040
rect 265992 447092 266044 447098
rect 265992 447034 266044 447040
rect 266004 444378 266032 447034
rect 265992 444372 266044 444378
rect 265992 444314 266044 444320
rect 266084 444372 266136 444378
rect 266084 444314 266136 444320
rect 266096 437510 266124 444314
rect 266084 437504 266136 437510
rect 266084 437446 266136 437452
rect 265992 437436 266044 437442
rect 265992 437378 266044 437384
rect 266004 434738 266032 437378
rect 266004 434710 266124 434738
rect 266096 429894 266124 434710
rect 265808 429888 265860 429894
rect 265808 429830 265860 429836
rect 266084 429888 266136 429894
rect 266084 429830 266136 429836
rect 265820 425202 265848 429830
rect 265808 425196 265860 425202
rect 265808 425138 265860 425144
rect 265992 425196 266044 425202
rect 265992 425138 266044 425144
rect 266004 425066 266032 425138
rect 265992 425060 266044 425066
rect 265992 425002 266044 425008
rect 266176 425060 266228 425066
rect 266176 425002 266228 425008
rect 266188 415449 266216 425002
rect 265990 415440 266046 415449
rect 265912 415398 265990 415426
rect 265912 411194 265940 415398
rect 265990 415375 266046 415384
rect 266174 415440 266230 415449
rect 266174 415375 266230 415384
rect 265716 411188 265768 411194
rect 265716 411130 265768 411136
rect 265900 411188 265952 411194
rect 265900 411130 265952 411136
rect 254584 411120 254636 411126
rect 254584 411062 254636 411068
rect 226156 410916 226208 410922
rect 226156 410858 226208 410864
rect 223396 410848 223448 410854
rect 223396 410790 223448 410796
rect 222292 409148 222344 409154
rect 222292 409090 222344 409096
rect 223408 408748 223436 410790
rect 226168 408748 226196 410858
rect 246028 410780 246080 410786
rect 246028 410722 246080 410728
rect 240324 410508 240376 410514
rect 240324 410450 240376 410456
rect 237564 410440 237616 410446
rect 237564 410382 237616 410388
rect 234620 410372 234672 410378
rect 234620 410314 234672 410320
rect 231860 410304 231912 410310
rect 231860 410246 231912 410252
rect 228916 410236 228968 410242
rect 228916 410178 228968 410184
rect 228928 408748 228956 410178
rect 231872 408748 231900 410246
rect 234632 408748 234660 410314
rect 237576 408748 237604 410382
rect 240336 408748 240364 410450
rect 243268 409964 243320 409970
rect 243268 409906 243320 409912
rect 243280 408748 243308 409906
rect 246040 408748 246068 410722
rect 254596 410582 254624 411062
rect 254676 411052 254728 411058
rect 254676 410994 254728 411000
rect 254584 410576 254636 410582
rect 254584 410518 254636 410524
rect 251732 410168 251784 410174
rect 251732 410110 251784 410116
rect 248972 410032 249024 410038
rect 248972 409974 249024 409980
rect 248984 408748 249012 409974
rect 251744 408748 251772 410110
rect 254688 408748 254716 410994
rect 258724 410984 258776 410990
rect 258724 410926 258776 410932
rect 258736 410718 258764 410926
rect 258724 410712 258776 410718
rect 258724 410654 258776 410660
rect 258816 410712 258868 410718
rect 258816 410654 258868 410660
rect 257252 410576 257304 410582
rect 257252 410518 257304 410524
rect 257264 410378 257292 410518
rect 258828 410446 258856 410654
rect 258816 410440 258868 410446
rect 258816 410382 258868 410388
rect 260380 410440 260432 410446
rect 260380 410382 260432 410388
rect 257252 410372 257304 410378
rect 257252 410314 257304 410320
rect 257344 410372 257396 410378
rect 257344 410314 257396 410320
rect 257356 410174 257384 410314
rect 257344 410168 257396 410174
rect 257344 410110 257396 410116
rect 257436 410168 257488 410174
rect 257436 410110 257488 410116
rect 257448 408748 257476 410110
rect 260392 408748 260420 410382
rect 263140 409964 263192 409970
rect 263140 409906 263192 409912
rect 263152 408748 263180 409906
rect 265728 408406 265756 411130
rect 269580 411120 269632 411126
rect 269580 411062 269632 411068
rect 266360 411052 266412 411058
rect 266360 410994 266412 411000
rect 265900 409896 265952 409902
rect 265900 409838 265952 409844
rect 265912 408748 265940 409838
rect 265716 408400 265768 408406
rect 265716 408342 265768 408348
rect 266084 408400 266136 408406
rect 266084 408342 266136 408348
rect 266096 398834 266124 408342
rect 266096 398806 266216 398834
rect 266188 392630 266216 398806
rect 266176 392624 266228 392630
rect 266176 392566 266228 392572
rect 200212 342780 200264 342786
rect 200212 342722 200264 342728
rect 240140 340536 240192 340542
rect 240138 340504 240140 340513
rect 240192 340504 240194 340513
rect 202788 340468 202840 340474
rect 202788 340410 202840 340416
rect 215208 340468 215260 340474
rect 215208 340410 215260 340416
rect 240048 340468 240100 340474
rect 240138 340439 240194 340448
rect 249706 340504 249762 340513
rect 249706 340439 249708 340448
rect 240048 340410 240100 340416
rect 249760 340439 249762 340448
rect 259458 340504 259514 340513
rect 259458 340439 259460 340448
rect 249708 340410 249760 340416
rect 259512 340439 259514 340448
rect 259460 340410 259512 340416
rect 202800 340377 202828 340410
rect 202786 340368 202842 340377
rect 215220 340354 215248 340410
rect 224960 340400 225012 340406
rect 215220 340338 215432 340354
rect 224880 340348 224960 340354
rect 230480 340400 230532 340406
rect 224880 340342 225012 340348
rect 230478 340368 230480 340377
rect 240060 340377 240088 340410
rect 230532 340368 230534 340377
rect 224880 340338 225000 340342
rect 215220 340332 215444 340338
rect 215220 340326 215392 340332
rect 202786 340303 202842 340312
rect 215392 340274 215444 340280
rect 224868 340332 225000 340338
rect 224920 340326 225000 340332
rect 230478 340303 230534 340312
rect 240046 340368 240102 340377
rect 240046 340303 240102 340312
rect 224868 340274 224920 340280
rect 200592 336870 200620 340068
rect 203352 337754 203380 340068
rect 203340 337748 203392 337754
rect 203340 337690 203392 337696
rect 206112 337686 206140 340068
rect 209070 340054 209728 340082
rect 207664 337748 207716 337754
rect 207664 337690 207716 337696
rect 206100 337680 206152 337686
rect 206100 337622 206152 337628
rect 200580 336864 200632 336870
rect 200580 336806 200632 336812
rect 201408 336864 201460 336870
rect 201408 336806 201460 336812
rect 200028 202700 200080 202706
rect 200028 202642 200080 202648
rect 199936 202428 199988 202434
rect 199936 202370 199988 202376
rect 201420 202298 201448 336806
rect 207676 202638 207704 337690
rect 209700 203454 209728 340054
rect 209780 339040 209832 339046
rect 209780 338982 209832 338988
rect 209792 215234 209820 338982
rect 211816 337822 211844 340068
rect 213920 338972 213972 338978
rect 213920 338914 213972 338920
rect 211804 337816 211856 337822
rect 211804 337758 211856 337764
rect 213932 222154 213960 338914
rect 214760 337754 214788 340068
rect 217534 340054 218008 340082
rect 215300 338904 215352 338910
rect 215300 338846 215352 338852
rect 214748 337748 214800 337754
rect 214748 337690 214800 337696
rect 213920 222148 213972 222154
rect 213920 222090 213972 222096
rect 214196 222148 214248 222154
rect 214196 222090 214248 222096
rect 209792 215206 209912 215234
rect 209884 205714 209912 215206
rect 214208 212566 214236 222090
rect 214196 212560 214248 212566
rect 214196 212502 214248 212508
rect 214380 212560 214432 212566
rect 214380 212502 214432 212508
rect 209884 205686 210004 205714
rect 209688 203448 209740 203454
rect 209688 203390 209740 203396
rect 202880 202632 202932 202638
rect 202880 202574 202932 202580
rect 207664 202632 207716 202638
rect 207664 202574 207716 202580
rect 201408 202292 201460 202298
rect 201408 202234 201460 202240
rect 199660 201884 199712 201890
rect 199660 201826 199712 201832
rect 198832 201544 198884 201550
rect 198832 201486 198884 201492
rect 202892 200002 202920 202574
rect 134168 199974 134228 200002
rect 134444 199974 134596 200002
rect 134720 199974 135056 200002
rect 142540 199974 142876 200002
rect 168392 199974 168544 200002
rect 168668 199974 169004 200002
rect 169128 199974 169372 200002
rect 176948 199974 177192 200002
rect 178052 199974 178112 200002
rect 178696 199974 178940 200002
rect 179524 199974 179860 200002
rect 180352 199974 180688 200002
rect 181272 199974 181608 200002
rect 182192 199974 182436 200002
rect 202860 199974 202920 200002
rect 209976 200002 210004 205686
rect 213458 202056 213514 202065
rect 213458 201991 213514 202000
rect 212540 201680 212592 201686
rect 212540 201622 212592 201628
rect 211160 201612 211212 201618
rect 211160 201554 211212 201560
rect 211172 200002 211200 201554
rect 211712 201544 211764 201550
rect 211712 201486 211764 201492
rect 209976 199974 210312 200002
rect 211140 199974 211200 200002
rect 211724 200002 211752 201486
rect 212552 200002 212580 201622
rect 213472 200002 213500 201991
rect 214392 200002 214420 212502
rect 215312 200002 215340 338846
rect 217980 202094 218008 340054
rect 220464 337890 220492 340068
rect 222200 338836 222252 338842
rect 222200 338778 222252 338784
rect 220820 338768 220872 338774
rect 220820 338710 220872 338716
rect 220452 337884 220504 337890
rect 220452 337826 220504 337832
rect 220358 202872 220414 202881
rect 220832 202842 220860 338710
rect 220358 202807 220414 202816
rect 220820 202836 220872 202842
rect 216864 202088 216916 202094
rect 216864 202030 216916 202036
rect 217968 202088 218020 202094
rect 217968 202030 218020 202036
rect 216036 201748 216088 201754
rect 216036 201690 216088 201696
rect 216048 200002 216076 201690
rect 216876 200002 216904 202030
rect 218060 201952 218112 201958
rect 218060 201894 218112 201900
rect 218072 200002 218100 201894
rect 219532 201884 219584 201890
rect 219532 201826 219584 201832
rect 218612 201816 218664 201822
rect 218612 201758 218664 201764
rect 218624 200002 218652 201758
rect 219544 200002 219572 201826
rect 220372 200002 220400 202807
rect 220820 202778 220872 202784
rect 221280 202836 221332 202842
rect 221280 202778 221332 202784
rect 220636 202768 220688 202774
rect 220636 202710 220688 202716
rect 220648 201958 220676 202710
rect 220636 201952 220688 201958
rect 220636 201894 220688 201900
rect 221292 200002 221320 202778
rect 222212 200002 222240 338778
rect 223224 337346 223252 340068
rect 226168 337958 226196 340068
rect 226156 337952 226208 337958
rect 226156 337894 226208 337900
rect 223212 337340 223264 337346
rect 223212 337282 223264 337288
rect 228928 337278 228956 340068
rect 231872 338026 231900 340068
rect 231860 338020 231912 338026
rect 231860 337962 231912 337968
rect 228916 337272 228968 337278
rect 228916 337214 228968 337220
rect 234632 336870 234660 340068
rect 237288 338768 237340 338774
rect 237288 338710 237340 338716
rect 236000 337272 236052 337278
rect 236000 337214 236052 337220
rect 234620 336864 234672 336870
rect 234620 336806 234672 336812
rect 231860 291848 231912 291854
rect 231860 291790 231912 291796
rect 231872 215234 231900 291790
rect 231872 215206 231992 215234
rect 231964 205714 231992 215206
rect 231964 205686 232176 205714
rect 230572 205148 230624 205154
rect 230572 205090 230624 205096
rect 229560 205080 229612 205086
rect 229560 205022 229612 205028
rect 225144 203380 225196 203386
rect 225144 203322 225196 203328
rect 223854 202736 223910 202745
rect 223854 202671 223910 202680
rect 223028 202020 223080 202026
rect 223028 201962 223080 201968
rect 223040 200002 223068 201962
rect 223868 200002 223896 202671
rect 225156 200002 225184 203322
rect 226892 202768 226944 202774
rect 226892 202710 226944 202716
rect 226338 202600 226394 202609
rect 226338 202535 226394 202544
rect 226352 200002 226380 202535
rect 211724 199974 211968 200002
rect 212552 199974 212888 200002
rect 213472 199974 213716 200002
rect 214392 199974 214636 200002
rect 215312 199974 215464 200002
rect 216048 199974 216384 200002
rect 216876 199974 217212 200002
rect 218072 199974 218132 200002
rect 218624 199974 218960 200002
rect 219544 199974 219880 200002
rect 220372 199974 220708 200002
rect 221292 199974 221536 200002
rect 222212 199974 222456 200002
rect 223040 199974 223284 200002
rect 223868 199974 224204 200002
rect 225156 199974 225492 200002
rect 226320 199974 226380 200002
rect 226904 200002 226932 202710
rect 228638 202464 228694 202473
rect 228638 202399 228694 202408
rect 227812 201952 227864 201958
rect 227812 201894 227864 201900
rect 227824 200002 227852 201894
rect 228652 200002 228680 202399
rect 229572 200002 229600 205022
rect 230584 200002 230612 205090
rect 231216 205012 231268 205018
rect 231216 204954 231268 204960
rect 231228 200002 231256 204954
rect 232148 200002 232176 205686
rect 233240 204944 233292 204950
rect 233240 204886 233292 204892
rect 236012 204898 236040 337214
rect 233252 200002 233280 204886
rect 236012 204870 236500 204898
rect 236368 202768 236420 202774
rect 236368 202710 236420 202716
rect 233422 202328 233478 202337
rect 233422 202263 233478 202272
rect 233436 200002 233464 202263
rect 236380 200002 236408 202710
rect 226904 199974 227240 200002
rect 227824 199974 228068 200002
rect 228652 199974 228988 200002
rect 229572 199974 229816 200002
rect 230584 199974 230736 200002
rect 231228 199974 231564 200002
rect 232148 199974 232484 200002
rect 233252 199974 233312 200002
rect 233436 199974 233772 200002
rect 236348 199974 236408 200002
rect 236472 200002 236500 204870
rect 237300 200002 237328 338710
rect 237576 336870 237604 340068
rect 240152 340054 240350 340082
rect 239404 337884 239456 337890
rect 239404 337826 239456 337832
rect 239416 337346 239444 337826
rect 237656 337340 237708 337346
rect 237656 337282 237708 337288
rect 239404 337340 239456 337346
rect 239404 337282 239456 337288
rect 237472 336864 237524 336870
rect 237472 336806 237524 336812
rect 237564 336864 237616 336870
rect 237564 336806 237616 336812
rect 237484 204950 237512 336806
rect 237472 204944 237524 204950
rect 237472 204886 237524 204892
rect 237668 200002 237696 337282
rect 239404 336864 239456 336870
rect 239404 336806 239456 336812
rect 240048 336864 240100 336870
rect 240048 336806 240100 336812
rect 237748 204944 237800 204950
rect 237748 204886 237800 204892
rect 236472 199974 236808 200002
rect 237268 199974 237328 200002
rect 237636 199974 237696 200002
rect 237760 200002 237788 204886
rect 238760 203516 238812 203522
rect 238760 203458 238812 203464
rect 238208 202700 238260 202706
rect 238208 202642 238260 202648
rect 238220 200002 238248 202642
rect 237760 199974 238096 200002
rect 238220 199974 238556 200002
rect 238772 199918 238800 203458
rect 239416 202638 239444 336806
rect 239680 202836 239732 202842
rect 239680 202778 239732 202784
rect 239312 202632 239364 202638
rect 239312 202574 239364 202580
rect 239404 202632 239456 202638
rect 239404 202574 239456 202580
rect 239220 202088 239272 202094
rect 239220 202030 239272 202036
rect 239232 200002 239260 202030
rect 239324 201890 239352 202574
rect 239312 201884 239364 201890
rect 239312 201826 239364 201832
rect 239692 200002 239720 202778
rect 240060 202094 240088 336806
rect 240152 202842 240180 340054
rect 240784 337816 240836 337822
rect 240784 337758 240836 337764
rect 242164 337816 242216 337822
rect 242164 337758 242216 337764
rect 240140 202836 240192 202842
rect 240140 202778 240192 202784
rect 240508 202836 240560 202842
rect 240508 202778 240560 202784
rect 240048 202088 240100 202094
rect 240048 202030 240100 202036
rect 240520 200002 240548 202778
rect 240796 202706 240824 337758
rect 240968 203516 241020 203522
rect 240968 203458 241020 203464
rect 240784 202700 240836 202706
rect 240784 202642 240836 202648
rect 240980 200002 241008 203458
rect 242176 202842 242204 337758
rect 242808 337272 242860 337278
rect 242808 337214 242860 337220
rect 242820 202842 242848 337214
rect 243096 336870 243124 340068
rect 244832 338020 244884 338026
rect 244832 337962 244884 337968
rect 243084 336864 243136 336870
rect 243084 336806 243136 336812
rect 244844 328506 244872 337962
rect 246040 337822 246068 340068
rect 248512 337952 248564 337958
rect 248512 337894 248564 337900
rect 246028 337816 246080 337822
rect 246028 337758 246080 337764
rect 246304 337340 246356 337346
rect 246304 337282 246356 337288
rect 244832 328500 244884 328506
rect 244832 328442 244884 328448
rect 244740 204264 244792 204270
rect 244740 204206 244792 204212
rect 243176 203448 243228 203454
rect 243176 203390 243228 203396
rect 242164 202836 242216 202842
rect 242164 202778 242216 202784
rect 242256 202836 242308 202842
rect 242256 202778 242308 202784
rect 242808 202836 242860 202842
rect 242808 202778 242860 202784
rect 241520 202564 241572 202570
rect 241520 202506 241572 202512
rect 241060 202496 241112 202502
rect 241060 202438 241112 202444
rect 238924 199974 239260 200002
rect 239384 199974 239720 200002
rect 240304 199974 240548 200002
rect 240672 199974 241008 200002
rect 241072 200002 241100 202438
rect 241532 200002 241560 202506
rect 242268 200002 242296 202778
rect 242348 202700 242400 202706
rect 242348 202642 242400 202648
rect 241072 199974 241132 200002
rect 241532 199974 241592 200002
rect 242052 199974 242296 200002
rect 242360 200002 242388 202642
rect 243084 201952 243136 201958
rect 243084 201894 243136 201900
rect 243096 200002 243124 201894
rect 242360 199974 242420 200002
rect 242880 199974 243124 200002
rect 243188 200002 243216 203390
rect 243820 202632 243872 202638
rect 243820 202574 243872 202580
rect 243728 202496 243780 202502
rect 243728 202438 243780 202444
rect 243740 200002 243768 202438
rect 243188 199974 243340 200002
rect 243708 199974 243768 200002
rect 243832 200002 243860 202574
rect 244648 201680 244700 201686
rect 244648 201622 244700 201628
rect 244660 200002 244688 201622
rect 243832 199974 244168 200002
rect 244628 199974 244688 200002
rect 244752 200002 244780 204206
rect 245660 204196 245712 204202
rect 245660 204138 245712 204144
rect 245200 202360 245252 202366
rect 245200 202302 245252 202308
rect 245212 200002 245240 202302
rect 245672 200002 245700 204138
rect 246316 202026 246344 337282
rect 247684 336864 247736 336870
rect 247684 336806 247736 336812
rect 247500 202564 247552 202570
rect 247500 202506 247552 202512
rect 246488 202428 246540 202434
rect 246488 202370 246540 202376
rect 246304 202020 246356 202026
rect 246304 201962 246356 201968
rect 246028 201816 246080 201822
rect 246028 201758 246080 201764
rect 246040 200002 246068 201758
rect 246500 200002 246528 202370
rect 247512 200002 247540 202506
rect 247592 202360 247644 202366
rect 247592 202302 247644 202308
rect 244752 199974 245088 200002
rect 245212 199974 245456 200002
rect 245672 199974 245916 200002
rect 246040 199974 246376 200002
rect 246500 199974 246836 200002
rect 247204 199974 247540 200002
rect 247604 200002 247632 202302
rect 247696 201958 247724 336806
rect 247684 201952 247736 201958
rect 247684 201894 247736 201900
rect 247776 201884 247828 201890
rect 247776 201826 247828 201832
rect 247788 200002 247816 201826
rect 248524 200002 248552 337894
rect 248800 336870 248828 340068
rect 250996 338020 251048 338026
rect 250996 337962 251048 337968
rect 249064 337816 249116 337822
rect 249064 337758 249116 337764
rect 249076 337278 249104 337758
rect 249064 337272 249116 337278
rect 249064 337214 249116 337220
rect 248788 336864 248840 336870
rect 248788 336806 248840 336812
rect 248696 328500 248748 328506
rect 248696 328442 248748 328448
rect 248708 200258 248736 328442
rect 250536 204196 250588 204202
rect 250536 204138 250588 204144
rect 248972 202632 249024 202638
rect 248972 202574 249024 202580
rect 248696 200252 248748 200258
rect 248696 200194 248748 200200
rect 248984 200002 249012 202574
rect 250076 201748 250128 201754
rect 250076 201690 250128 201696
rect 249386 200252 249438 200258
rect 249386 200194 249438 200200
rect 247604 199974 247664 200002
rect 247788 199974 248124 200002
rect 248492 199974 248552 200002
rect 248952 199974 249012 200002
rect 249398 199988 249426 200194
rect 250088 200002 250116 201690
rect 250548 200002 250576 204138
rect 250904 202700 250956 202706
rect 250904 202642 250956 202648
rect 250916 200002 250944 202642
rect 251008 201754 251036 337962
rect 251744 337278 251772 340068
rect 253756 337952 253808 337958
rect 253756 337894 253808 337900
rect 251732 337272 251784 337278
rect 251732 337214 251784 337220
rect 251916 204128 251968 204134
rect 251916 204070 251968 204076
rect 253572 204128 253624 204134
rect 253572 204070 253624 204076
rect 251456 202836 251508 202842
rect 251456 202778 251508 202784
rect 250996 201748 251048 201754
rect 250996 201690 251048 201696
rect 251468 200002 251496 202778
rect 251824 202088 251876 202094
rect 251824 202030 251876 202036
rect 251836 200002 251864 202030
rect 249872 199974 250116 200002
rect 250240 199974 250576 200002
rect 250700 199974 250944 200002
rect 251160 199974 251496 200002
rect 251620 199974 251864 200002
rect 251928 200002 251956 204070
rect 252652 202496 252704 202502
rect 252650 202464 252652 202473
rect 252704 202464 252706 202473
rect 252650 202399 252706 202408
rect 253480 202360 253532 202366
rect 253478 202328 253480 202337
rect 253532 202328 253534 202337
rect 253478 202263 253534 202272
rect 253112 202020 253164 202026
rect 253112 201962 253164 201968
rect 252744 201476 252796 201482
rect 252744 201418 252796 201424
rect 252756 200002 252784 201418
rect 253124 200002 253152 201962
rect 253584 200002 253612 204070
rect 253768 202178 253796 337894
rect 254504 336870 254532 340068
rect 257448 337822 257476 340068
rect 257988 338836 258040 338842
rect 257988 338778 258040 338784
rect 257436 337816 257488 337822
rect 257436 337758 257488 337764
rect 255596 337680 255648 337686
rect 255596 337622 255648 337628
rect 254492 336864 254544 336870
rect 254492 336806 254544 336812
rect 255608 323626 255636 337622
rect 255608 323598 255820 323626
rect 255792 318850 255820 323598
rect 255780 318844 255832 318850
rect 255780 318786 255832 318792
rect 255872 318844 255924 318850
rect 255872 318786 255924 318792
rect 255884 309233 255912 318786
rect 258000 318782 258028 338778
rect 260208 338026 260236 340068
rect 262128 338632 262180 338638
rect 262128 338574 262180 338580
rect 260196 338020 260248 338026
rect 260196 337962 260248 337968
rect 258724 337748 258776 337754
rect 258724 337690 258776 337696
rect 258448 336864 258500 336870
rect 258448 336806 258500 336812
rect 258460 336734 258488 336806
rect 258172 336728 258224 336734
rect 258172 336670 258224 336676
rect 258448 336728 258500 336734
rect 258448 336670 258500 336676
rect 258184 327146 258212 336670
rect 258172 327140 258224 327146
rect 258172 327082 258224 327088
rect 258356 327140 258408 327146
rect 258356 327082 258408 327088
rect 258368 327049 258396 327082
rect 258170 327040 258226 327049
rect 258170 326975 258226 326984
rect 258354 327040 258410 327049
rect 258354 326975 258410 326984
rect 257712 318776 257764 318782
rect 257712 318718 257764 318724
rect 257988 318776 258040 318782
rect 257988 318718 258040 318724
rect 255594 309224 255650 309233
rect 255594 309159 255650 309168
rect 255870 309224 255926 309233
rect 257724 309194 257752 318718
rect 258184 317490 258212 326975
rect 258172 317484 258224 317490
rect 258172 317426 258224 317432
rect 258632 317484 258684 317490
rect 258632 317426 258684 317432
rect 258644 309233 258672 317426
rect 258354 309224 258410 309233
rect 255870 309159 255926 309168
rect 257712 309188 257764 309194
rect 255608 299470 255636 309159
rect 257712 309130 257764 309136
rect 257804 309188 257856 309194
rect 258354 309159 258410 309168
rect 258630 309224 258686 309233
rect 258630 309159 258686 309168
rect 257804 309130 257856 309136
rect 257816 302138 257844 309130
rect 257816 302110 257936 302138
rect 257908 299470 257936 302110
rect 258368 299470 258396 309159
rect 255504 299464 255556 299470
rect 255504 299406 255556 299412
rect 255596 299464 255648 299470
rect 255596 299406 255648 299412
rect 257712 299464 257764 299470
rect 257712 299406 257764 299412
rect 257896 299464 257948 299470
rect 257896 299406 257948 299412
rect 258264 299464 258316 299470
rect 258264 299406 258316 299412
rect 258356 299464 258408 299470
rect 258356 299406 258408 299412
rect 255516 289950 255544 299406
rect 255504 289944 255556 289950
rect 255504 289886 255556 289892
rect 257724 289882 257752 299406
rect 258276 289950 258304 299406
rect 258264 289944 258316 289950
rect 258264 289886 258316 289892
rect 255596 289876 255648 289882
rect 255596 289818 255648 289824
rect 257712 289876 257764 289882
rect 257712 289818 257764 289824
rect 257804 289876 257856 289882
rect 257804 289818 257856 289824
rect 258356 289876 258408 289882
rect 258356 289818 258408 289824
rect 255608 269090 255636 289818
rect 257816 282946 257844 289818
rect 257804 282940 257856 282946
rect 257804 282882 257856 282888
rect 257988 282940 258040 282946
rect 257988 282882 258040 282888
rect 255608 269062 255728 269090
rect 255700 260914 255728 269062
rect 255688 260908 255740 260914
rect 255688 260850 255740 260856
rect 255688 260772 255740 260778
rect 255688 260714 255740 260720
rect 255700 251002 255728 260714
rect 255424 250974 255728 251002
rect 255424 236706 255452 250974
rect 258000 241505 258028 282882
rect 258368 277386 258396 289818
rect 258276 277358 258396 277386
rect 258276 276010 258304 277358
rect 258264 276004 258316 276010
rect 258264 275946 258316 275952
rect 258356 276004 258408 276010
rect 258356 275946 258408 275952
rect 258368 258074 258396 275946
rect 258368 258046 258488 258074
rect 258460 249150 258488 258046
rect 258448 249144 258500 249150
rect 258448 249086 258500 249092
rect 258448 249008 258500 249014
rect 258448 248950 258500 248956
rect 257986 241496 258042 241505
rect 257986 241431 258042 241440
rect 258170 241496 258226 241505
rect 258170 241431 258226 241440
rect 255412 236700 255464 236706
rect 255412 236642 255464 236648
rect 255596 236700 255648 236706
rect 255596 236642 255648 236648
rect 255608 222222 255636 236642
rect 258184 231878 258212 241431
rect 258460 240174 258488 248950
rect 258264 240168 258316 240174
rect 258264 240110 258316 240116
rect 258448 240168 258500 240174
rect 258448 240110 258500 240116
rect 258276 238746 258304 240110
rect 258264 238740 258316 238746
rect 258264 238682 258316 238688
rect 258448 238740 258500 238746
rect 258448 238682 258500 238688
rect 257988 231872 258040 231878
rect 257988 231814 258040 231820
rect 258172 231872 258224 231878
rect 258172 231814 258224 231820
rect 258000 224890 258028 231814
rect 258460 229106 258488 238682
rect 258460 229078 258580 229106
rect 257908 224862 258028 224890
rect 255596 222216 255648 222222
rect 255596 222158 255648 222164
rect 255688 222216 255740 222222
rect 255688 222158 255740 222164
rect 257908 222170 257936 224862
rect 255700 212566 255728 222158
rect 257908 222142 258028 222170
rect 258000 212566 258028 222142
rect 258552 215422 258580 229078
rect 258540 215416 258592 215422
rect 258540 215358 258592 215364
rect 258448 215280 258500 215286
rect 258448 215222 258500 215228
rect 255596 212560 255648 212566
rect 255596 212502 255648 212508
rect 255688 212560 255740 212566
rect 255688 212502 255740 212508
rect 257804 212560 257856 212566
rect 257804 212502 257856 212508
rect 257988 212560 258040 212566
rect 257988 212502 258040 212508
rect 255608 211546 255636 212502
rect 255596 211540 255648 211546
rect 255596 211482 255648 211488
rect 256148 211540 256200 211546
rect 256148 211482 256200 211488
rect 255780 204264 255832 204270
rect 255780 204206 255832 204212
rect 254032 204060 254084 204066
rect 254032 204002 254084 204008
rect 253848 202564 253900 202570
rect 253848 202506 253900 202512
rect 253676 202150 253796 202178
rect 253676 202026 253704 202150
rect 253664 202020 253716 202026
rect 253664 201962 253716 201968
rect 253756 202020 253808 202026
rect 253756 201962 253808 201968
rect 253768 200002 253796 201962
rect 253860 201686 253888 202506
rect 253940 202428 253992 202434
rect 253940 202370 253992 202376
rect 253952 202337 253980 202370
rect 253938 202328 253994 202337
rect 253938 202263 253994 202272
rect 253848 201680 253900 201686
rect 253848 201622 253900 201628
rect 251928 199974 251988 200002
rect 252448 199974 252784 200002
rect 252908 199974 253152 200002
rect 253276 199974 253612 200002
rect 253736 199974 253796 200002
rect 254044 200002 254072 204002
rect 254124 202496 254176 202502
rect 254122 202464 254124 202473
rect 254176 202464 254178 202473
rect 254122 202399 254178 202408
rect 254860 201748 254912 201754
rect 254860 201690 254912 201696
rect 254872 200002 254900 201690
rect 254998 200252 255050 200258
rect 254998 200194 255050 200200
rect 254044 199974 254196 200002
rect 254656 199974 254900 200002
rect 255010 199988 255038 200194
rect 255792 200002 255820 204206
rect 255964 204060 256016 204066
rect 255964 204002 256016 204008
rect 255976 200002 256004 204002
rect 255484 199974 255820 200002
rect 255944 199974 256004 200002
rect 256160 200002 256188 211482
rect 257816 205714 257844 212502
rect 257816 205686 257936 205714
rect 257908 205578 257936 205686
rect 257724 205550 257936 205578
rect 257160 203924 257212 203930
rect 257160 203866 257212 203872
rect 256516 202224 256568 202230
rect 256516 202166 256568 202172
rect 256528 201822 256556 202166
rect 257068 201884 257120 201890
rect 257068 201826 257120 201832
rect 256516 201816 256568 201822
rect 256516 201758 256568 201764
rect 257080 200002 257108 201826
rect 256160 199974 256404 200002
rect 256772 199974 257108 200002
rect 257172 200002 257200 203866
rect 257724 202824 257752 205550
rect 258460 204082 258488 215222
rect 258460 204054 258672 204082
rect 258448 203992 258500 203998
rect 258448 203934 258500 203940
rect 257632 202796 257752 202824
rect 257632 200138 257660 202796
rect 258356 201680 258408 201686
rect 258356 201622 258408 201628
rect 257632 200110 257706 200138
rect 257172 199974 257232 200002
rect 257678 199988 257706 200110
rect 258368 200002 258396 201622
rect 258060 199974 258396 200002
rect 258460 200002 258488 203934
rect 258538 202328 258594 202337
rect 258538 202263 258540 202272
rect 258592 202263 258594 202272
rect 258540 202234 258592 202240
rect 258644 200138 258672 204054
rect 258736 202774 258764 337690
rect 260104 337272 260156 337278
rect 260104 337214 260156 337220
rect 259828 203924 259880 203930
rect 259828 203866 259880 203872
rect 258816 202904 258868 202910
rect 258816 202846 258868 202852
rect 258724 202768 258776 202774
rect 258724 202710 258776 202716
rect 258828 202026 258856 202846
rect 259000 202836 259052 202842
rect 259000 202778 259052 202784
rect 259012 202230 259040 202778
rect 259458 202328 259514 202337
rect 259458 202263 259514 202272
rect 259000 202224 259052 202230
rect 259000 202166 259052 202172
rect 258908 202156 258960 202162
rect 258908 202098 258960 202104
rect 258724 202020 258776 202026
rect 258724 201962 258776 201968
rect 258816 202020 258868 202026
rect 258816 201962 258868 201968
rect 258736 201618 258764 201962
rect 258724 201612 258776 201618
rect 258724 201554 258776 201560
rect 258920 200258 258948 202098
rect 258908 200252 258960 200258
rect 258908 200194 258960 200200
rect 258644 200110 258764 200138
rect 258736 200002 258764 200110
rect 259472 200002 259500 202263
rect 259840 200002 259868 203866
rect 260116 202842 260144 337214
rect 260380 203856 260432 203862
rect 260380 203798 260432 203804
rect 260104 202836 260156 202842
rect 260104 202778 260156 202784
rect 259920 201816 259972 201822
rect 259920 201758 259972 201764
rect 258460 199974 258520 200002
rect 258736 199974 258980 200002
rect 259440 199974 259500 200002
rect 259808 199974 259868 200002
rect 259932 200002 259960 201758
rect 260392 200002 260420 203798
rect 262140 202314 262168 338574
rect 263152 337958 263180 340068
rect 263140 337952 263192 337958
rect 263140 337894 263192 337900
rect 265912 336870 265940 340068
rect 265900 336864 265952 336870
rect 265900 336806 265952 336812
rect 262772 203788 262824 203794
rect 262772 203730 262824 203736
rect 261772 202286 262168 202314
rect 260840 201952 260892 201958
rect 260840 201894 260892 201900
rect 260852 200002 260880 201894
rect 261772 200002 261800 202286
rect 261942 202192 261998 202201
rect 261942 202127 261998 202136
rect 259932 199974 260268 200002
rect 260392 199974 260728 200002
rect 260852 199974 261188 200002
rect 261556 199974 261800 200002
rect 261956 200002 261984 202127
rect 262680 201748 262732 201754
rect 262680 201690 262732 201696
rect 262692 200002 262720 201690
rect 261956 199974 262016 200002
rect 262476 199974 262720 200002
rect 262784 200002 262812 203730
rect 262956 203720 263008 203726
rect 262956 203662 263008 203668
rect 262968 200002 262996 203662
rect 265440 203652 265492 203658
rect 265440 203594 265492 203600
rect 263600 202836 263652 202842
rect 263600 202778 263652 202784
rect 263612 200002 263640 202778
rect 263876 202768 263928 202774
rect 263876 202710 263928 202716
rect 264888 202768 264940 202774
rect 264888 202710 264940 202716
rect 263888 200002 263916 202710
rect 264900 200002 264928 202710
rect 265348 201952 265400 201958
rect 265348 201894 265400 201900
rect 265360 200002 265388 201894
rect 262784 199974 262844 200002
rect 262968 199974 263304 200002
rect 263612 199974 263764 200002
rect 263888 199974 264224 200002
rect 264592 199974 264928 200002
rect 265052 199974 265388 200002
rect 265452 200002 265480 203594
rect 266268 202836 266320 202842
rect 266268 202778 266320 202784
rect 266280 202502 266308 202778
rect 266268 202496 266320 202502
rect 266268 202438 266320 202444
rect 266084 202360 266136 202366
rect 266084 202302 266136 202308
rect 266176 202360 266228 202366
rect 266176 202302 266228 202308
rect 266096 201890 266124 202302
rect 265992 201884 266044 201890
rect 265992 201826 266044 201832
rect 266084 201884 266136 201890
rect 266084 201826 266136 201832
rect 266004 201754 266032 201826
rect 265900 201748 265952 201754
rect 265900 201690 265952 201696
rect 265992 201748 266044 201754
rect 265992 201690 266044 201696
rect 265912 201482 265940 201690
rect 265900 201476 265952 201482
rect 265900 201418 265952 201424
rect 266188 200002 266216 202302
rect 266372 201618 266400 410994
rect 267004 410984 267056 410990
rect 267004 410926 267056 410932
rect 266544 410848 266596 410854
rect 266544 410790 266596 410796
rect 266452 410508 266504 410514
rect 266452 410450 266504 410456
rect 266464 202026 266492 410450
rect 266452 202020 266504 202026
rect 266452 201962 266504 201968
rect 266556 201906 266584 410790
rect 266728 410712 266780 410718
rect 266728 410654 266780 410660
rect 266636 410032 266688 410038
rect 266636 409974 266688 409980
rect 266464 201878 266584 201906
rect 266648 201906 266676 409974
rect 266740 202230 266768 410654
rect 266818 399664 266874 399673
rect 266818 399599 266874 399608
rect 266728 202224 266780 202230
rect 266728 202166 266780 202172
rect 266832 201958 266860 399599
rect 266910 382800 266966 382809
rect 266910 382735 266966 382744
rect 266924 204270 266952 382735
rect 266912 204264 266964 204270
rect 266912 204206 266964 204212
rect 267016 201958 267044 410926
rect 269212 410576 269264 410582
rect 269212 410518 269264 410524
rect 267280 410440 267332 410446
rect 267280 410382 267332 410388
rect 267094 357504 267150 357513
rect 267094 357439 267150 357448
rect 266820 201952 266872 201958
rect 266648 201878 266768 201906
rect 266820 201894 266872 201900
rect 267004 201952 267056 201958
rect 267004 201894 267056 201900
rect 266464 201822 266492 201878
rect 266452 201816 266504 201822
rect 266452 201758 266504 201764
rect 266740 201686 266768 201878
rect 267108 201736 267136 357439
rect 267186 349072 267242 349081
rect 267186 349007 267242 349016
rect 267200 203930 267228 349007
rect 267292 338842 267320 410382
rect 267372 409964 267424 409970
rect 267372 409906 267424 409912
rect 267280 338836 267332 338842
rect 267280 338778 267332 338784
rect 267384 338774 267412 409906
rect 268752 409896 268804 409902
rect 268752 409838 268804 409844
rect 267738 403744 267794 403753
rect 267738 403679 267794 403688
rect 267372 338768 267424 338774
rect 267372 338710 267424 338716
rect 267188 203924 267240 203930
rect 267188 203866 267240 203872
rect 267188 203584 267240 203590
rect 267188 203526 267240 203532
rect 266832 201708 267136 201736
rect 266728 201680 266780 201686
rect 266728 201622 266780 201628
rect 266360 201612 266412 201618
rect 266360 201554 266412 201560
rect 266452 201544 266504 201550
rect 266636 201544 266688 201550
rect 266504 201492 266636 201498
rect 266452 201486 266688 201492
rect 266464 201470 266676 201486
rect 266832 200138 266860 201708
rect 267096 201612 267148 201618
rect 267096 201554 267148 201560
rect 266648 200110 266860 200138
rect 266648 200002 266676 200110
rect 267108 200002 267136 201554
rect 265452 199974 265512 200002
rect 265972 199974 266216 200002
rect 266340 199974 266676 200002
rect 266800 199974 267136 200002
rect 267200 200002 267228 203526
rect 267648 202496 267700 202502
rect 267648 202438 267700 202444
rect 267660 200002 267688 202438
rect 267752 202094 267780 403679
rect 267830 395312 267886 395321
rect 267830 395247 267886 395256
rect 267844 204202 267872 395247
rect 267922 391232 267978 391241
rect 267922 391167 267978 391176
rect 267832 204196 267884 204202
rect 267832 204138 267884 204144
rect 267936 202570 267964 391167
rect 268014 386880 268070 386889
rect 268014 386815 268070 386824
rect 267924 202564 267976 202570
rect 267924 202506 267976 202512
rect 268028 202434 268056 386815
rect 268106 378448 268162 378457
rect 268106 378383 268162 378392
rect 268120 202638 268148 378383
rect 268198 374368 268254 374377
rect 268198 374303 268254 374312
rect 268108 202632 268160 202638
rect 268108 202574 268160 202580
rect 268016 202428 268068 202434
rect 268016 202370 268068 202376
rect 267740 202088 267792 202094
rect 268212 202042 268240 374303
rect 268290 370016 268346 370025
rect 268290 369951 268346 369960
rect 268304 202162 268332 369951
rect 268382 365936 268438 365945
rect 268382 365871 268438 365880
rect 268396 204066 268424 365871
rect 268474 361584 268530 361593
rect 268474 361519 268530 361528
rect 268488 210458 268516 361519
rect 268566 353424 268622 353433
rect 268566 353359 268622 353368
rect 268476 210452 268528 210458
rect 268476 210394 268528 210400
rect 268384 204060 268436 204066
rect 268384 204002 268436 204008
rect 268580 203522 268608 353359
rect 268658 344992 268714 345001
rect 268658 344927 268714 344936
rect 268672 204134 268700 344927
rect 268764 338638 268792 409838
rect 268948 340598 269068 340626
rect 268948 340513 268976 340598
rect 269040 340542 269068 340598
rect 269028 340536 269080 340542
rect 268934 340504 268990 340513
rect 269028 340478 269080 340484
rect 269118 340504 269174 340513
rect 268934 340439 268990 340448
rect 269118 340439 269120 340448
rect 269172 340439 269174 340448
rect 269120 340410 269172 340416
rect 268752 338632 268804 338638
rect 268752 338574 268804 338580
rect 268844 210452 268896 210458
rect 268844 210394 268896 210400
rect 268660 204128 268712 204134
rect 268660 204070 268712 204076
rect 268568 203516 268620 203522
rect 268568 203458 268620 203464
rect 268292 202156 268344 202162
rect 268292 202098 268344 202104
rect 267740 202030 267792 202036
rect 268028 202014 268240 202042
rect 268028 201550 268056 202014
rect 268200 201952 268252 201958
rect 268200 201894 268252 201900
rect 268108 201748 268160 201754
rect 268108 201690 268160 201696
rect 268016 201544 268068 201550
rect 268016 201486 268068 201492
rect 268120 200002 268148 201690
rect 267200 199974 267260 200002
rect 267628 199974 267688 200002
rect 268088 199974 268148 200002
rect 268212 200002 268240 201894
rect 268856 200002 268884 210394
rect 269224 202706 269252 410518
rect 269304 410372 269356 410378
rect 269304 410314 269356 410320
rect 269212 202700 269264 202706
rect 269212 202642 269264 202648
rect 269316 202502 269344 410314
rect 269396 410168 269448 410174
rect 269396 410110 269448 410116
rect 269408 202842 269436 410110
rect 269488 410100 269540 410106
rect 269488 410042 269540 410048
rect 269396 202836 269448 202842
rect 269396 202778 269448 202784
rect 269500 202774 269528 410042
rect 269488 202768 269540 202774
rect 269488 202710 269540 202716
rect 269304 202496 269356 202502
rect 269304 202438 269356 202444
rect 269592 202366 269620 411062
rect 269672 336864 269724 336870
rect 269672 336806 269724 336812
rect 269580 202360 269632 202366
rect 269580 202302 269632 202308
rect 269684 200002 269712 336806
rect 269764 202292 269816 202298
rect 269764 202234 269816 202240
rect 268212 199974 268548 200002
rect 268856 199974 269008 200002
rect 269376 199974 269712 200002
rect 269776 200002 269804 202234
rect 270420 200002 270448 583578
rect 282828 583568 282880 583574
rect 282828 583510 282880 583516
rect 275928 583160 275980 583166
rect 275928 583102 275980 583108
rect 274548 582752 274600 582758
rect 274548 582694 274600 582700
rect 273168 578944 273220 578950
rect 273168 578886 273220 578892
rect 273180 578542 273208 578886
rect 273168 578536 273220 578542
rect 273168 578478 273220 578484
rect 271788 569968 271840 569974
rect 271788 569910 271840 569916
rect 271800 563145 271828 569910
rect 271786 563136 271842 563145
rect 271786 563071 271842 563080
rect 271694 563000 271750 563009
rect 271694 562935 271750 562944
rect 271708 560289 271736 562935
rect 271510 560280 271566 560289
rect 271510 560215 271566 560224
rect 271694 560280 271750 560289
rect 271694 560215 271750 560224
rect 271524 550662 271552 560215
rect 273168 556232 273220 556238
rect 273168 556174 273220 556180
rect 271512 550656 271564 550662
rect 271512 550598 271564 550604
rect 271788 550656 271840 550662
rect 271788 550598 271840 550604
rect 271800 545834 271828 550598
rect 271512 545828 271564 545834
rect 271512 545770 271564 545776
rect 271788 545828 271840 545834
rect 271788 545770 271840 545776
rect 271524 541006 271552 545770
rect 271512 541000 271564 541006
rect 271512 540942 271564 540948
rect 271604 541000 271656 541006
rect 271694 540968 271750 540977
rect 271656 540948 271694 540954
rect 271604 540942 271694 540948
rect 271616 540926 271694 540942
rect 271694 540903 271750 540912
rect 271970 540968 272026 540977
rect 271970 540903 272026 540912
rect 271984 531350 272012 540903
rect 271788 531344 271840 531350
rect 271788 531286 271840 531292
rect 271972 531344 272024 531350
rect 271972 531286 272024 531292
rect 271800 524550 271828 531286
rect 271788 524544 271840 524550
rect 271788 524486 271840 524492
rect 271788 524408 271840 524414
rect 271788 524350 271840 524356
rect 271800 514826 271828 524350
rect 271788 514820 271840 514826
rect 271788 514762 271840 514768
rect 271696 514752 271748 514758
rect 271696 514694 271748 514700
rect 271708 512038 271736 514694
rect 271696 512032 271748 512038
rect 271696 511974 271748 511980
rect 271788 512032 271840 512038
rect 271788 511974 271840 511980
rect 271800 507210 271828 511974
rect 271512 507204 271564 507210
rect 271512 507146 271564 507152
rect 271788 507204 271840 507210
rect 271788 507146 271840 507152
rect 271524 502382 271552 507146
rect 271512 502376 271564 502382
rect 271604 502376 271656 502382
rect 271512 502318 271564 502324
rect 271602 502344 271604 502353
rect 271656 502344 271658 502353
rect 271602 502279 271658 502288
rect 271786 492688 271842 492697
rect 271786 492623 271842 492632
rect 271800 487830 271828 492623
rect 271512 487824 271564 487830
rect 271512 487766 271564 487772
rect 271788 487824 271840 487830
rect 271788 487766 271840 487772
rect 271524 483138 271552 487766
rect 271512 483132 271564 483138
rect 271512 483074 271564 483080
rect 271696 483132 271748 483138
rect 271696 483074 271748 483080
rect 271708 483002 271736 483074
rect 271696 482996 271748 483002
rect 271696 482938 271748 482944
rect 271788 482996 271840 483002
rect 271788 482938 271840 482944
rect 271800 476134 271828 482938
rect 271788 476128 271840 476134
rect 271788 476070 271840 476076
rect 271696 476060 271748 476066
rect 271696 476002 271748 476008
rect 271708 473362 271736 476002
rect 271708 473334 271828 473362
rect 271800 468518 271828 473334
rect 271512 468512 271564 468518
rect 271512 468454 271564 468460
rect 271788 468512 271840 468518
rect 271788 468454 271840 468460
rect 271524 463826 271552 468454
rect 271512 463820 271564 463826
rect 271512 463762 271564 463768
rect 271696 463820 271748 463826
rect 271696 463762 271748 463768
rect 271708 463690 271736 463762
rect 271696 463684 271748 463690
rect 271696 463626 271748 463632
rect 271788 463684 271840 463690
rect 271788 463626 271840 463632
rect 271800 456822 271828 463626
rect 271788 456816 271840 456822
rect 271788 456758 271840 456764
rect 271696 456748 271748 456754
rect 271696 456690 271748 456696
rect 271708 454050 271736 456690
rect 271708 454022 271828 454050
rect 271800 449206 271828 454022
rect 271512 449200 271564 449206
rect 271512 449142 271564 449148
rect 271788 449200 271840 449206
rect 271788 449142 271840 449148
rect 271524 444514 271552 449142
rect 271512 444508 271564 444514
rect 271512 444450 271564 444456
rect 271696 444508 271748 444514
rect 271696 444450 271748 444456
rect 271708 444378 271736 444450
rect 271696 444372 271748 444378
rect 271696 444314 271748 444320
rect 271788 444372 271840 444378
rect 271788 444314 271840 444320
rect 271800 437510 271828 444314
rect 271788 437504 271840 437510
rect 271788 437446 271840 437452
rect 271696 437436 271748 437442
rect 271696 437378 271748 437384
rect 271708 434738 271736 437378
rect 271708 434710 271828 434738
rect 271800 429894 271828 434710
rect 271512 429888 271564 429894
rect 271512 429830 271564 429836
rect 271788 429888 271840 429894
rect 271788 429830 271840 429836
rect 271524 425202 271552 429830
rect 271512 425196 271564 425202
rect 271512 425138 271564 425144
rect 271696 425196 271748 425202
rect 271696 425138 271748 425144
rect 271708 425066 271736 425138
rect 271696 425060 271748 425066
rect 271696 425002 271748 425008
rect 271788 425060 271840 425066
rect 271788 425002 271840 425008
rect 271800 419529 271828 425002
rect 271786 419520 271842 419529
rect 271786 419455 271842 419464
rect 271970 419520 272026 419529
rect 271970 419455 272026 419464
rect 270776 410916 270828 410922
rect 270776 410858 270828 410864
rect 270684 410780 270736 410786
rect 270684 410722 270736 410728
rect 270500 410644 270552 410650
rect 270500 410586 270552 410592
rect 270512 201618 270540 410586
rect 270592 410236 270644 410242
rect 270592 410178 270644 410184
rect 270604 201754 270632 410178
rect 270696 201890 270724 410722
rect 270684 201884 270736 201890
rect 270684 201826 270736 201832
rect 270592 201748 270644 201754
rect 270592 201690 270644 201696
rect 270788 201686 270816 410858
rect 270868 410304 270920 410310
rect 270868 410246 270920 410252
rect 270880 201822 270908 410246
rect 271984 408542 272012 419455
rect 271604 408536 271656 408542
rect 271604 408478 271656 408484
rect 271972 408536 272024 408542
rect 271972 408478 272024 408484
rect 271616 398818 271644 408478
rect 271604 398812 271656 398818
rect 271604 398754 271656 398760
rect 271788 398812 271840 398818
rect 271788 398754 271840 398760
rect 271800 389201 271828 398754
rect 271602 389192 271658 389201
rect 271512 389156 271564 389162
rect 271602 389127 271604 389136
rect 271512 389098 271564 389104
rect 271656 389127 271658 389136
rect 271786 389192 271842 389201
rect 271786 389127 271842 389136
rect 271604 389098 271656 389104
rect 271524 384266 271552 389098
rect 271512 384260 271564 384266
rect 271512 384202 271564 384208
rect 271696 384260 271748 384266
rect 271696 384202 271748 384208
rect 271708 379522 271736 384202
rect 271708 379506 271828 379522
rect 271696 379500 271840 379506
rect 271748 379494 271788 379500
rect 271696 379442 271748 379448
rect 271788 379442 271840 379448
rect 271708 360262 271736 379442
rect 271800 379411 271828 379442
rect 271696 360256 271748 360262
rect 271696 360198 271748 360204
rect 271788 360256 271840 360262
rect 271788 360198 271840 360204
rect 271800 336938 271828 360198
rect 271788 336932 271840 336938
rect 271788 336874 271840 336880
rect 271696 336864 271748 336870
rect 271696 336806 271748 336812
rect 271708 332602 271736 336806
rect 271616 332574 271736 332602
rect 271616 330546 271644 332574
rect 271420 330540 271472 330546
rect 271420 330482 271472 330488
rect 271604 330540 271656 330546
rect 271604 330482 271656 330488
rect 271432 325718 271460 330482
rect 271420 325712 271472 325718
rect 271420 325654 271472 325660
rect 271512 325712 271564 325718
rect 271512 325654 271564 325660
rect 271524 322930 271552 325654
rect 271512 322924 271564 322930
rect 271512 322866 271564 322872
rect 271696 322924 271748 322930
rect 271696 322866 271748 322872
rect 271708 313290 271736 322866
rect 271708 313262 271828 313290
rect 271800 303618 271828 313262
rect 271788 303612 271840 303618
rect 271788 303554 271840 303560
rect 271972 303612 272024 303618
rect 271972 303554 272024 303560
rect 271984 294137 272012 303554
rect 271970 294128 272026 294137
rect 271970 294063 272026 294072
rect 271786 293992 271842 294001
rect 271786 293927 271842 293936
rect 271800 284306 271828 293927
rect 271788 284300 271840 284306
rect 271788 284242 271840 284248
rect 271972 284300 272024 284306
rect 271972 284242 272024 284248
rect 271984 274825 272012 284242
rect 271970 274816 272026 274825
rect 271970 274751 272026 274760
rect 271786 274680 271842 274689
rect 271786 274615 271842 274624
rect 271800 264926 271828 274615
rect 271604 264920 271656 264926
rect 271604 264862 271656 264868
rect 271788 264920 271840 264926
rect 271788 264862 271840 264868
rect 271616 255377 271644 264862
rect 271602 255368 271658 255377
rect 271602 255303 271658 255312
rect 271786 255368 271842 255377
rect 271786 255303 271842 255312
rect 271800 255270 271828 255303
rect 271420 255264 271472 255270
rect 271420 255206 271472 255212
rect 271788 255264 271840 255270
rect 271788 255206 271840 255212
rect 271432 245682 271460 255206
rect 271420 245676 271472 245682
rect 271420 245618 271472 245624
rect 271512 245676 271564 245682
rect 271512 245618 271564 245624
rect 271524 242214 271552 245618
rect 271512 242208 271564 242214
rect 271512 242150 271564 242156
rect 271788 242208 271840 242214
rect 271788 242150 271840 242156
rect 271800 227746 271828 242150
rect 271800 227730 271920 227746
rect 271696 227724 271748 227730
rect 271800 227724 271932 227730
rect 271800 227718 271880 227724
rect 271696 227666 271748 227672
rect 271880 227666 271932 227672
rect 271708 218074 271736 227666
rect 271892 227635 271920 227666
rect 271696 218068 271748 218074
rect 271696 218010 271748 218016
rect 271972 218068 272024 218074
rect 271972 218010 272024 218016
rect 271984 212566 272012 218010
rect 271512 212560 271564 212566
rect 271512 212502 271564 212508
rect 271972 212560 272024 212566
rect 271972 212502 272024 212508
rect 271524 205714 271552 212502
rect 271432 205686 271552 205714
rect 270960 202224 271012 202230
rect 270960 202166 271012 202172
rect 270868 201816 270920 201822
rect 270868 201758 270920 201764
rect 270776 201680 270828 201686
rect 270776 201622 270828 201628
rect 270500 201612 270552 201618
rect 270500 201554 270552 201560
rect 270972 200002 271000 202166
rect 271432 200002 271460 205686
rect 271788 203652 271840 203658
rect 271788 203594 271840 203600
rect 271800 200002 271828 203594
rect 273180 201754 273208 556174
rect 274456 347064 274508 347070
rect 274456 347006 274508 347012
rect 273258 340504 273314 340513
rect 273258 340439 273260 340448
rect 273312 340439 273314 340448
rect 273260 340410 273312 340416
rect 273996 202496 274048 202502
rect 273996 202438 274048 202444
rect 272248 201748 272300 201754
rect 272248 201690 272300 201696
rect 273168 201748 273220 201754
rect 273168 201690 273220 201696
rect 273628 201748 273680 201754
rect 273628 201690 273680 201696
rect 272260 200002 272288 201690
rect 273640 200002 273668 201690
rect 274008 200002 274036 202438
rect 274468 201754 274496 347006
rect 274560 202502 274588 582694
rect 275836 497208 275888 497214
rect 275836 497150 275888 497156
rect 275652 212560 275704 212566
rect 275652 212502 275704 212508
rect 274548 202496 274600 202502
rect 274548 202438 274600 202444
rect 274456 201748 274508 201754
rect 274456 201690 274508 201696
rect 275284 201748 275336 201754
rect 275284 201690 275336 201696
rect 275296 200002 275324 201690
rect 275664 200002 275692 212502
rect 275848 201754 275876 497150
rect 275940 212566 275968 583102
rect 281172 583092 281224 583098
rect 281172 583034 281224 583040
rect 281184 580666 281212 583034
rect 281184 580638 281304 580666
rect 277952 578944 278004 578950
rect 277952 578886 278004 578892
rect 277964 578474 277992 578886
rect 278044 578876 278096 578882
rect 278044 578818 278096 578824
rect 278056 578678 278084 578818
rect 278044 578672 278096 578678
rect 278044 578614 278096 578620
rect 277952 578468 278004 578474
rect 277952 578410 278004 578416
rect 281276 572762 281304 580638
rect 281264 572756 281316 572762
rect 281264 572698 281316 572704
rect 281264 572620 281316 572626
rect 281264 572562 281316 572568
rect 281276 569838 281304 572562
rect 281080 569832 281132 569838
rect 281080 569774 281132 569780
rect 281264 569832 281316 569838
rect 281264 569774 281316 569780
rect 281092 560318 281120 569774
rect 281080 560312 281132 560318
rect 281080 560254 281132 560260
rect 281264 560312 281316 560318
rect 281264 560254 281316 560260
rect 281276 553450 281304 560254
rect 281264 553444 281316 553450
rect 281264 553386 281316 553392
rect 281356 553376 281408 553382
rect 281356 553318 281408 553324
rect 281368 550662 281396 553318
rect 281264 550656 281316 550662
rect 281264 550598 281316 550604
rect 281356 550656 281408 550662
rect 281356 550598 281408 550604
rect 281276 550526 281304 550598
rect 281080 550520 281132 550526
rect 281080 550462 281132 550468
rect 281264 550520 281316 550526
rect 281264 550462 281316 550468
rect 281092 541006 281120 550462
rect 281080 541000 281132 541006
rect 281080 540942 281132 540948
rect 281264 541000 281316 541006
rect 281264 540942 281316 540948
rect 281276 534138 281304 540942
rect 281264 534132 281316 534138
rect 281264 534074 281316 534080
rect 281356 534064 281408 534070
rect 281356 534006 281408 534012
rect 281368 531350 281396 534006
rect 281264 531344 281316 531350
rect 281264 531286 281316 531292
rect 281356 531344 281408 531350
rect 281356 531286 281408 531292
rect 281276 524550 281304 531286
rect 281264 524544 281316 524550
rect 281264 524486 281316 524492
rect 281264 524408 281316 524414
rect 281264 524350 281316 524356
rect 281276 521937 281304 524350
rect 281262 521928 281318 521937
rect 281262 521863 281318 521872
rect 280068 521688 280120 521694
rect 281354 521690 281410 521699
rect 280068 521630 280120 521636
rect 281276 521634 281354 521642
rect 278688 518968 278740 518974
rect 278688 518910 278740 518916
rect 277308 497140 277360 497146
rect 277308 497082 277360 497088
rect 275928 212560 275980 212566
rect 275928 212502 275980 212508
rect 277320 202314 277348 497082
rect 276952 202286 277348 202314
rect 275836 201748 275888 201754
rect 275836 201690 275888 201696
rect 276952 200002 276980 202286
rect 277306 202192 277362 202201
rect 277306 202127 277362 202136
rect 277320 200002 277348 202127
rect 278700 200002 278728 518910
rect 280080 201754 280108 521630
rect 281276 521625 281410 521634
rect 281276 521614 281396 521625
rect 281276 514826 281304 521614
rect 282736 516180 282788 516186
rect 282736 516122 282788 516128
rect 281264 514820 281316 514826
rect 281264 514762 281316 514768
rect 281356 514752 281408 514758
rect 281356 514694 281408 514700
rect 281368 512038 281396 514694
rect 281264 512032 281316 512038
rect 281264 511974 281316 511980
rect 281356 512032 281408 512038
rect 281356 511974 281408 511980
rect 281276 511902 281304 511974
rect 281080 511896 281132 511902
rect 281080 511838 281132 511844
rect 281264 511896 281316 511902
rect 281264 511838 281316 511844
rect 281092 502382 281120 511838
rect 281080 502376 281132 502382
rect 281080 502318 281132 502324
rect 281264 502376 281316 502382
rect 281264 502318 281316 502324
rect 281276 497622 281304 502318
rect 281080 497616 281132 497622
rect 281080 497558 281132 497564
rect 281264 497616 281316 497622
rect 281264 497558 281316 497564
rect 281092 492697 281120 497558
rect 281078 492688 281134 492697
rect 281078 492623 281134 492632
rect 281262 492688 281318 492697
rect 281262 492623 281318 492632
rect 281276 485926 281304 492623
rect 281264 485920 281316 485926
rect 281264 485862 281316 485868
rect 281264 485784 281316 485790
rect 281264 485726 281316 485732
rect 281276 476134 281304 485726
rect 281264 476128 281316 476134
rect 281264 476070 281316 476076
rect 281356 476128 281408 476134
rect 281356 476070 281408 476076
rect 281368 473414 281396 476070
rect 281264 473408 281316 473414
rect 281264 473350 281316 473356
rect 281356 473408 281408 473414
rect 281356 473350 281408 473356
rect 281276 466546 281304 473350
rect 281264 466540 281316 466546
rect 281264 466482 281316 466488
rect 281264 466404 281316 466410
rect 281264 466346 281316 466352
rect 281276 458862 281304 466346
rect 281080 458856 281132 458862
rect 281080 458798 281132 458804
rect 281264 458856 281316 458862
rect 281264 458798 281316 458804
rect 281092 454073 281120 458798
rect 281078 454064 281134 454073
rect 281078 453999 281134 454008
rect 281262 454064 281318 454073
rect 281262 453999 281318 454008
rect 281276 447234 281304 453999
rect 281264 447228 281316 447234
rect 281264 447170 281316 447176
rect 281264 447092 281316 447098
rect 281264 447034 281316 447040
rect 281276 439550 281304 447034
rect 281080 439544 281132 439550
rect 281080 439486 281132 439492
rect 281264 439544 281316 439550
rect 281264 439486 281316 439492
rect 281092 434761 281120 439486
rect 281078 434752 281134 434761
rect 281078 434687 281134 434696
rect 281262 434752 281318 434761
rect 281262 434687 281318 434696
rect 281276 427922 281304 434687
rect 281264 427916 281316 427922
rect 281264 427858 281316 427864
rect 281264 427780 281316 427786
rect 281264 427722 281316 427728
rect 281276 423638 281304 427722
rect 281264 423632 281316 423638
rect 281264 423574 281316 423580
rect 281540 423632 281592 423638
rect 281540 423574 281592 423580
rect 281552 414066 281580 423574
rect 281552 414038 281672 414066
rect 281644 413982 281672 414038
rect 281632 413976 281684 413982
rect 281632 413918 281684 413924
rect 281816 413976 281868 413982
rect 281816 413918 281868 413924
rect 281828 404954 281856 413918
rect 281644 404926 281856 404954
rect 281644 396137 281672 404926
rect 281630 396128 281686 396137
rect 281630 396063 281686 396072
rect 281630 395992 281686 396001
rect 281630 395927 281686 395936
rect 281644 386458 281672 395927
rect 281368 386430 281672 386458
rect 281368 386374 281396 386430
rect 281356 386368 281408 386374
rect 281356 386310 281408 386316
rect 281540 386368 281592 386374
rect 281540 386310 281592 386316
rect 281552 376854 281580 386310
rect 281172 376848 281224 376854
rect 281172 376790 281224 376796
rect 281540 376848 281592 376854
rect 281540 376790 281592 376796
rect 281184 376718 281212 376790
rect 281080 376712 281132 376718
rect 281080 376654 281132 376660
rect 281172 376712 281224 376718
rect 281172 376654 281224 376660
rect 281092 367198 281120 376654
rect 281080 367192 281132 367198
rect 281080 367134 281132 367140
rect 281356 367192 281408 367198
rect 281356 367134 281408 367140
rect 281368 367062 281396 367134
rect 281080 367056 281132 367062
rect 281080 366998 281132 367004
rect 281356 367056 281408 367062
rect 281356 366998 281408 367004
rect 281092 357542 281120 366998
rect 281080 357536 281132 357542
rect 281080 357478 281132 357484
rect 281172 357536 281224 357542
rect 281172 357478 281224 357484
rect 281184 357406 281212 357478
rect 281080 357400 281132 357406
rect 281080 357342 281132 357348
rect 281172 357400 281224 357406
rect 281172 357342 281224 357348
rect 281092 347886 281120 357342
rect 281080 347880 281132 347886
rect 281080 347822 281132 347828
rect 281356 347880 281408 347886
rect 281356 347822 281408 347828
rect 281368 347750 281396 347822
rect 281080 347744 281132 347750
rect 281080 347686 281132 347692
rect 281356 347744 281408 347750
rect 281356 347686 281408 347692
rect 280160 340536 280212 340542
rect 280160 340478 280212 340484
rect 280172 340338 280200 340478
rect 280160 340332 280212 340338
rect 280160 340274 280212 340280
rect 281092 338162 281120 347686
rect 281080 338156 281132 338162
rect 281080 338098 281132 338104
rect 281264 338156 281316 338162
rect 281264 338098 281316 338104
rect 281276 338042 281304 338098
rect 281184 338014 281304 338042
rect 281184 328506 281212 338014
rect 281172 328500 281224 328506
rect 281172 328442 281224 328448
rect 281264 328500 281316 328506
rect 281264 328442 281316 328448
rect 281276 321570 281304 328442
rect 281264 321564 281316 321570
rect 281264 321506 281316 321512
rect 281356 321564 281408 321570
rect 281356 321506 281408 321512
rect 281368 318782 281396 321506
rect 281080 318776 281132 318782
rect 281080 318718 281132 318724
rect 281356 318776 281408 318782
rect 281356 318718 281408 318724
rect 281092 309194 281120 318718
rect 281080 309188 281132 309194
rect 281080 309130 281132 309136
rect 281264 309188 281316 309194
rect 281264 309130 281316 309136
rect 281276 302258 281304 309130
rect 281264 302252 281316 302258
rect 281264 302194 281316 302200
rect 281356 302184 281408 302190
rect 281356 302126 281408 302132
rect 281368 299470 281396 302126
rect 281080 299464 281132 299470
rect 281080 299406 281132 299412
rect 281356 299464 281408 299470
rect 281356 299406 281408 299412
rect 281092 289882 281120 299406
rect 281080 289876 281132 289882
rect 281080 289818 281132 289824
rect 281264 289876 281316 289882
rect 281264 289818 281316 289824
rect 281276 282946 281304 289818
rect 281264 282940 281316 282946
rect 281264 282882 281316 282888
rect 281356 282872 281408 282878
rect 281356 282814 281408 282820
rect 281368 280158 281396 282814
rect 281356 280152 281408 280158
rect 281356 280094 281408 280100
rect 281632 280152 281684 280158
rect 281632 280094 281684 280100
rect 281644 270638 281672 280094
rect 281356 270632 281408 270638
rect 281356 270574 281408 270580
rect 281632 270632 281684 270638
rect 281632 270574 281684 270580
rect 281368 270502 281396 270574
rect 281080 270496 281132 270502
rect 281080 270438 281132 270444
rect 281356 270496 281408 270502
rect 281356 270438 281408 270444
rect 281092 260914 281120 270438
rect 281080 260908 281132 260914
rect 281080 260850 281132 260856
rect 281264 260908 281316 260914
rect 281264 260850 281316 260856
rect 281170 260808 281226 260817
rect 281276 260794 281304 260850
rect 281226 260766 281304 260794
rect 281170 260743 281226 260752
rect 281078 251152 281134 251161
rect 281078 251087 281134 251096
rect 281092 241534 281120 251087
rect 281080 241528 281132 241534
rect 281080 241470 281132 241476
rect 281264 241528 281316 241534
rect 281264 241470 281316 241476
rect 281276 241398 281304 241470
rect 281080 241392 281132 241398
rect 281080 241334 281132 241340
rect 281264 241392 281316 241398
rect 281264 241334 281316 241340
rect 281092 231878 281120 241334
rect 281080 231872 281132 231878
rect 281080 231814 281132 231820
rect 281264 231872 281316 231878
rect 281264 231814 281316 231820
rect 281276 227066 281304 231814
rect 281092 227038 281304 227066
rect 281092 222222 281120 227038
rect 281080 222216 281132 222222
rect 281080 222158 281132 222164
rect 281172 222216 281224 222222
rect 281172 222158 281224 222164
rect 281184 215354 281212 222158
rect 281172 215348 281224 215354
rect 281172 215290 281224 215296
rect 281264 215212 281316 215218
rect 281264 215154 281316 215160
rect 280528 203584 280580 203590
rect 280528 203526 280580 203532
rect 279240 201748 279292 201754
rect 279240 201690 279292 201696
rect 280068 201748 280120 201754
rect 280068 201690 280120 201696
rect 279252 200002 279280 201690
rect 280540 200002 280568 203526
rect 281276 202502 281304 215154
rect 282748 202502 282776 516122
rect 280988 202496 281040 202502
rect 280988 202438 281040 202444
rect 281264 202496 281316 202502
rect 281264 202438 281316 202444
rect 282276 202496 282328 202502
rect 282276 202438 282328 202444
rect 282736 202496 282788 202502
rect 282736 202438 282788 202444
rect 281000 200002 281028 202438
rect 282288 200002 282316 202438
rect 282840 200138 282868 583510
rect 289728 583228 289780 583234
rect 289728 583170 289780 583176
rect 282920 579012 282972 579018
rect 282920 578954 282972 578960
rect 282932 578814 282960 578954
rect 287704 578876 287756 578882
rect 287704 578818 287756 578824
rect 282920 578808 282972 578814
rect 282920 578750 282972 578756
rect 287716 578610 287744 578818
rect 287704 578604 287756 578610
rect 287704 578546 287756 578552
rect 286968 538280 287020 538286
rect 286968 538222 287020 538228
rect 284208 497752 284260 497758
rect 284208 497694 284260 497700
rect 284116 497616 284168 497622
rect 284116 497558 284168 497564
rect 283932 202632 283984 202638
rect 283932 202574 283984 202580
rect 283564 202156 283616 202162
rect 283564 202098 283616 202104
rect 282748 200110 282868 200138
rect 282748 200002 282776 200110
rect 283576 200002 283604 202098
rect 283944 200002 283972 202574
rect 269776 199974 269836 200002
rect 270296 199974 270448 200002
rect 270664 199974 271000 200002
rect 271124 199974 271460 200002
rect 271584 199974 271828 200002
rect 272044 199974 272288 200002
rect 273332 199974 273668 200002
rect 273792 199974 274036 200002
rect 275080 199974 275324 200002
rect 275448 199974 275692 200002
rect 276828 199974 276980 200002
rect 277196 199974 277348 200002
rect 278576 199974 278728 200002
rect 278944 199974 279280 200002
rect 280232 199974 280568 200002
rect 280692 199974 281028 200002
rect 281980 199974 282316 200002
rect 282440 199974 282776 200002
rect 283360 199974 283604 200002
rect 283728 199974 283972 200002
rect 284128 200002 284156 497558
rect 284220 202638 284248 497694
rect 285588 497344 285640 497350
rect 285588 497286 285640 497292
rect 284208 202632 284260 202638
rect 284208 202574 284260 202580
rect 285600 200002 285628 497286
rect 286232 204944 286284 204950
rect 286232 204886 286284 204892
rect 286244 200002 286272 204886
rect 286980 200002 287008 538222
rect 289636 497412 289688 497418
rect 289636 497354 289688 497360
rect 288256 497072 288308 497078
rect 288256 497014 288308 497020
rect 288268 215234 288296 497014
rect 288084 215206 288296 215234
rect 288084 205714 288112 215206
rect 287992 205686 288112 205714
rect 287520 203720 287572 203726
rect 287520 203662 287572 203668
rect 287532 200002 287560 203662
rect 287992 200002 288020 205686
rect 289268 202836 289320 202842
rect 289268 202778 289320 202784
rect 288808 202496 288860 202502
rect 288808 202438 288860 202444
rect 288820 200002 288848 202438
rect 289280 200002 289308 202778
rect 289648 200002 289676 497354
rect 289740 202842 289768 583170
rect 293868 583024 293920 583030
rect 293868 582966 293920 582972
rect 291108 582820 291160 582826
rect 291108 582762 291160 582768
rect 289818 578912 289874 578921
rect 289818 578847 289820 578856
rect 289872 578847 289874 578856
rect 289820 578818 289872 578824
rect 291016 497684 291068 497690
rect 291016 497626 291068 497632
rect 290924 210452 290976 210458
rect 290924 210394 290976 210400
rect 289728 202836 289780 202842
rect 289728 202778 289780 202784
rect 290556 202836 290608 202842
rect 290556 202778 290608 202784
rect 290568 200002 290596 202778
rect 290936 200138 290964 210394
rect 291028 202842 291056 497626
rect 291120 210458 291148 582762
rect 293776 509312 293828 509318
rect 293776 509254 293828 509260
rect 292396 497276 292448 497282
rect 292396 497218 292448 497224
rect 291108 210452 291160 210458
rect 291108 210394 291160 210400
rect 292408 202842 292436 497218
rect 292488 340400 292540 340406
rect 292540 340348 292712 340354
rect 292488 340342 292712 340348
rect 292500 340338 292712 340342
rect 292500 340332 292724 340338
rect 292500 340326 292672 340332
rect 292672 340274 292724 340280
rect 292488 203788 292540 203794
rect 292488 203730 292540 203736
rect 291016 202836 291068 202842
rect 291016 202778 291068 202784
rect 291384 202836 291436 202842
rect 291384 202778 291436 202784
rect 292396 202836 292448 202842
rect 292396 202778 292448 202784
rect 290936 200110 291056 200138
rect 291028 200002 291056 200110
rect 291396 200002 291424 202778
rect 292304 202292 292356 202298
rect 292304 202234 292356 202240
rect 292316 200002 292344 202234
rect 292500 200002 292528 203730
rect 293132 202836 293184 202842
rect 293132 202778 293184 202784
rect 293144 200002 293172 202778
rect 293788 200002 293816 509254
rect 293880 202842 293908 582966
rect 300400 582956 300452 582962
rect 300400 582898 300452 582904
rect 298928 582684 298980 582690
rect 298928 582626 298980 582632
rect 298744 582480 298796 582486
rect 298744 582422 298796 582428
rect 297180 579012 297232 579018
rect 297180 578954 297232 578960
rect 294604 578944 294656 578950
rect 294604 578886 294656 578892
rect 294512 578604 294564 578610
rect 294512 578546 294564 578552
rect 294524 578474 294552 578546
rect 294616 578474 294644 578886
rect 297088 578740 297140 578746
rect 297088 578682 297140 578688
rect 297100 578474 297128 578682
rect 297192 578678 297220 578954
rect 298008 578876 298060 578882
rect 298008 578818 298060 578824
rect 297180 578672 297232 578678
rect 297180 578614 297232 578620
rect 294512 578468 294564 578474
rect 294512 578410 294564 578416
rect 294604 578468 294656 578474
rect 294604 578410 294656 578416
rect 297088 578468 297140 578474
rect 297088 578410 297140 578416
rect 296718 575784 296774 575793
rect 296718 575719 296774 575728
rect 296732 575550 296760 575719
rect 296720 575544 296772 575550
rect 296720 575486 296772 575492
rect 297362 572928 297418 572937
rect 297362 572863 297418 572872
rect 296718 570072 296774 570081
rect 296718 570007 296774 570016
rect 296732 569974 296760 570007
rect 296720 569968 296772 569974
rect 296720 569910 296772 569916
rect 296442 566128 296498 566137
rect 296442 566063 296498 566072
rect 294604 532772 294656 532778
rect 294604 532714 294656 532720
rect 294616 521626 294644 532714
rect 293960 521620 294012 521626
rect 293960 521562 294012 521568
rect 294604 521620 294656 521626
rect 294604 521562 294656 521568
rect 293972 521286 294000 521562
rect 293960 521280 294012 521286
rect 293960 521222 294012 521228
rect 293972 406570 294000 521222
rect 293960 406564 294012 406570
rect 293960 406506 294012 406512
rect 293972 406434 294000 406506
rect 293960 406428 294012 406434
rect 293960 406370 294012 406376
rect 294604 406428 294656 406434
rect 294604 406370 294656 406376
rect 294616 385694 294644 406370
rect 294604 385688 294656 385694
rect 294604 385630 294656 385636
rect 294880 205012 294932 205018
rect 294880 204954 294932 204960
rect 294420 203448 294472 203454
rect 294420 203390 294472 203396
rect 293868 202836 293920 202842
rect 293868 202778 293920 202784
rect 294432 200002 294460 203390
rect 294892 200002 294920 204954
rect 296168 203516 296220 203522
rect 296168 203458 296220 203464
rect 295800 202836 295852 202842
rect 295800 202778 295852 202784
rect 295812 200002 295840 202778
rect 296180 200002 296208 203458
rect 296456 202842 296484 566063
rect 296718 563272 296774 563281
rect 296718 563207 296774 563216
rect 296732 563106 296760 563207
rect 296720 563100 296772 563106
rect 296720 563042 296772 563048
rect 297270 541104 297326 541113
rect 297270 541039 297326 541048
rect 296534 531584 296590 531593
rect 296534 531519 296590 531528
rect 296444 202836 296496 202842
rect 296444 202778 296496 202784
rect 296548 200002 296576 531519
rect 296718 509552 296774 509561
rect 296718 509487 296774 509496
rect 296732 509318 296760 509487
rect 296720 509312 296772 509318
rect 296720 509254 296772 509260
rect 296718 506560 296774 506569
rect 296718 506495 296720 506504
rect 296772 506495 296774 506504
rect 296720 506466 296772 506472
rect 297180 505096 297232 505102
rect 297180 505038 297232 505044
rect 297192 495514 297220 505038
rect 297180 495508 297232 495514
rect 297180 495450 297232 495456
rect 297180 389156 297232 389162
rect 297180 389098 297232 389104
rect 297192 379574 297220 389098
rect 297180 379568 297232 379574
rect 297180 379510 297232 379516
rect 297284 337618 297312 541039
rect 297376 532778 297404 572863
rect 297914 560416 297970 560425
rect 297914 560351 297970 560360
rect 297822 556880 297878 556889
rect 297822 556815 297878 556824
rect 297836 556238 297864 556815
rect 297824 556232 297876 556238
rect 297824 556174 297876 556180
rect 297822 553616 297878 553625
rect 297822 553551 297878 553560
rect 297730 550760 297786 550769
rect 297730 550695 297786 550704
rect 297638 538384 297694 538393
rect 297638 538319 297694 538328
rect 297652 538286 297680 538319
rect 297640 538280 297692 538286
rect 297640 538222 297692 538228
rect 297638 534848 297694 534857
rect 297638 534783 297694 534792
rect 297364 532772 297416 532778
rect 297364 532714 297416 532720
rect 297362 528592 297418 528601
rect 297362 528527 297418 528536
rect 297376 518226 297404 528527
rect 297454 525872 297510 525881
rect 297454 525807 297510 525816
rect 297468 521506 297496 525807
rect 297546 522064 297602 522073
rect 297546 521999 297602 522008
rect 297560 521694 297588 521999
rect 297548 521688 297600 521694
rect 297548 521630 297600 521636
rect 297468 521478 297588 521506
rect 297454 519072 297510 519081
rect 297454 519007 297510 519016
rect 297468 518974 297496 519007
rect 297456 518968 297508 518974
rect 297456 518910 297508 518916
rect 297364 518220 297416 518226
rect 297364 518162 297416 518168
rect 297454 516216 297510 516225
rect 297454 516151 297456 516160
rect 297508 516151 297510 516160
rect 297456 516122 297508 516128
rect 297454 513496 297510 513505
rect 297454 513431 297510 513440
rect 297362 503840 297418 503849
rect 297362 503775 297418 503784
rect 297272 337612 297324 337618
rect 297272 337554 297324 337560
rect 297272 215280 297324 215286
rect 297272 215222 297324 215228
rect 297284 205698 297312 215222
rect 297272 205692 297324 205698
rect 297272 205634 297324 205640
rect 297272 201884 297324 201890
rect 297272 201826 297324 201832
rect 297284 200002 297312 201826
rect 297376 201686 297404 503775
rect 297468 202094 297496 513431
rect 297560 202366 297588 521478
rect 297548 202360 297600 202366
rect 297548 202302 297600 202308
rect 297456 202088 297508 202094
rect 297456 202030 297508 202036
rect 297364 201680 297416 201686
rect 297364 201622 297416 201628
rect 297652 201550 297680 534783
rect 297744 210458 297772 550695
rect 297836 211138 297864 553551
rect 297824 211132 297876 211138
rect 297824 211074 297876 211080
rect 297732 210452 297784 210458
rect 297732 210394 297784 210400
rect 297824 205692 297876 205698
rect 297824 205634 297876 205640
rect 297640 201544 297692 201550
rect 297640 201486 297692 201492
rect 297836 200138 297864 205634
rect 297928 203318 297956 560351
rect 298020 505102 298048 578818
rect 298008 505096 298060 505102
rect 298008 505038 298060 505044
rect 298008 495508 298060 495514
rect 298008 495450 298060 495456
rect 298020 389162 298048 495450
rect 298008 389156 298060 389162
rect 298008 389098 298060 389104
rect 298008 379568 298060 379574
rect 298008 379510 298060 379516
rect 298020 215286 298048 379510
rect 298008 215280 298060 215286
rect 298008 215222 298060 215228
rect 297916 203312 297968 203318
rect 297916 203254 297968 203260
rect 298376 201748 298428 201754
rect 298376 201690 298428 201696
rect 297836 200110 297956 200138
rect 297928 200002 297956 200110
rect 298388 200002 298416 201690
rect 298756 201618 298784 582422
rect 298836 582412 298888 582418
rect 298836 582354 298888 582360
rect 298848 499458 298876 582354
rect 298836 499452 298888 499458
rect 298836 499394 298888 499400
rect 298940 499050 298968 582626
rect 300308 582616 300360 582622
rect 300308 582558 300360 582564
rect 299296 582548 299348 582554
rect 299296 582490 299348 582496
rect 299204 579692 299256 579698
rect 299204 579634 299256 579640
rect 299110 547904 299166 547913
rect 299110 547839 299166 547848
rect 299018 544096 299074 544105
rect 299018 544031 299074 544040
rect 298928 499044 298980 499050
rect 298928 498986 298980 498992
rect 299032 202638 299060 544031
rect 299124 202706 299152 547839
rect 299112 202700 299164 202706
rect 299112 202642 299164 202648
rect 299020 202632 299072 202638
rect 299020 202574 299072 202580
rect 299216 202434 299244 579634
rect 299308 202570 299336 582490
rect 300216 579488 300268 579494
rect 300216 579430 300268 579436
rect 299480 579352 299532 579358
rect 299480 579294 299532 579300
rect 299386 578912 299442 578921
rect 299386 578847 299442 578856
rect 299400 578814 299428 578847
rect 299388 578808 299440 578814
rect 299388 578750 299440 578756
rect 299388 203856 299440 203862
rect 299388 203798 299440 203804
rect 299296 202564 299348 202570
rect 299296 202506 299348 202512
rect 299204 202428 299256 202434
rect 299204 202370 299256 202376
rect 299204 201952 299256 201958
rect 299204 201894 299256 201900
rect 298744 201612 298796 201618
rect 298744 201554 298796 201560
rect 299216 200002 299244 201894
rect 299400 200002 299428 203798
rect 299492 202774 299520 579294
rect 299572 579216 299624 579222
rect 299572 579158 299624 579164
rect 299584 579018 299612 579158
rect 300228 579086 300256 579430
rect 300216 579080 300268 579086
rect 300216 579022 300268 579028
rect 299572 579012 299624 579018
rect 299572 578954 299624 578960
rect 300216 578944 300268 578950
rect 300216 578886 300268 578892
rect 300228 578814 300256 578886
rect 300216 578808 300268 578814
rect 300216 578750 300268 578756
rect 300124 578740 300176 578746
rect 300124 578682 300176 578688
rect 300136 578542 300164 578682
rect 300124 578536 300176 578542
rect 300124 578478 300176 578484
rect 300320 498982 300348 582558
rect 300308 498976 300360 498982
rect 300308 498918 300360 498924
rect 299572 490612 299624 490618
rect 299572 490554 299624 490560
rect 299584 337550 299612 490554
rect 299572 337544 299624 337550
rect 299572 337486 299624 337492
rect 300124 202836 300176 202842
rect 300124 202778 300176 202784
rect 299480 202768 299532 202774
rect 299480 202710 299532 202716
rect 300136 200002 300164 202778
rect 300412 201822 300440 582898
rect 300492 582888 300544 582894
rect 300492 582830 300544 582836
rect 300504 202026 300532 582830
rect 302804 579972 302832 583646
rect 307024 583636 307076 583642
rect 307024 583578 307076 583584
rect 307036 579972 307064 583578
rect 313464 583568 313516 583574
rect 313464 583510 313516 583516
rect 309232 582412 309284 582418
rect 309232 582354 309284 582360
rect 309244 579972 309272 582354
rect 313476 579972 313504 583510
rect 317696 583500 317748 583506
rect 317696 583442 317748 583448
rect 317708 579972 317736 583442
rect 347504 583432 347556 583438
rect 347504 583374 347556 583380
rect 324136 583364 324188 583370
rect 324136 583306 324188 583312
rect 319720 583160 319772 583166
rect 319720 583102 319772 583108
rect 319732 579972 319760 583102
rect 321928 582480 321980 582486
rect 321928 582422 321980 582428
rect 321940 579972 321968 582422
rect 324148 579972 324176 583306
rect 328368 583228 328420 583234
rect 328368 583170 328420 583176
rect 326160 583092 326212 583098
rect 326160 583034 326212 583040
rect 326172 579972 326200 583034
rect 328380 579972 328408 583170
rect 338856 583024 338908 583030
rect 338856 582966 338908 582972
rect 332600 582548 332652 582554
rect 332600 582490 332652 582496
rect 332612 579972 332640 582490
rect 338868 579972 338896 582966
rect 341064 582684 341116 582690
rect 341064 582626 341116 582632
rect 341076 579972 341104 582626
rect 347516 579972 347544 583374
rect 349528 583296 349580 583302
rect 349528 583238 349580 583244
rect 349540 579972 349568 583238
rect 353760 582956 353812 582962
rect 353760 582898 353812 582904
rect 351736 582820 351788 582826
rect 351736 582762 351788 582768
rect 351748 579972 351776 582762
rect 353772 579972 353800 582898
rect 355968 582888 356020 582894
rect 355968 582830 356020 582836
rect 355980 579972 356008 582830
rect 368664 582752 368716 582758
rect 368664 582694 368716 582700
rect 357992 582684 358044 582690
rect 357992 582626 358044 582632
rect 358004 579972 358032 582626
rect 362408 582616 362460 582622
rect 362408 582558 362460 582564
rect 366640 582616 366692 582622
rect 366640 582558 366692 582564
rect 362420 579972 362448 582558
rect 366652 579972 366680 582558
rect 368676 579972 368704 582694
rect 379060 582684 379112 582690
rect 379060 582626 379112 582632
rect 377588 582616 377640 582622
rect 377588 582558 377640 582564
rect 370872 582548 370924 582554
rect 370872 582490 370924 582496
rect 377312 582548 377364 582554
rect 377312 582490 377364 582496
rect 370884 579972 370912 582490
rect 372896 582480 372948 582486
rect 372896 582422 372948 582428
rect 372908 579972 372936 582422
rect 304828 579698 305026 579714
rect 304816 579692 305026 579698
rect 304868 579686 305026 579692
rect 334728 579686 334940 579714
rect 304816 579634 304868 579640
rect 305092 579624 305144 579630
rect 305092 579566 305144 579572
rect 315212 579624 315264 579630
rect 330760 579624 330812 579630
rect 315264 579572 315514 579578
rect 315212 579566 315514 579572
rect 330760 579566 330812 579572
rect 305104 579358 305132 579566
rect 315224 579550 315514 579566
rect 330668 579556 330720 579562
rect 330668 579498 330720 579504
rect 310980 579488 311032 579494
rect 330576 579488 330628 579494
rect 311032 579436 311282 579442
rect 310980 579430 311282 579436
rect 330576 579430 330628 579436
rect 310992 579414 311282 579430
rect 330588 579358 330616 579430
rect 330680 579358 330708 579498
rect 330772 579358 330800 579566
rect 334728 579358 334756 579686
rect 334808 579624 334860 579630
rect 334808 579566 334860 579572
rect 334820 579358 334848 579566
rect 334912 579358 334940 579686
rect 335176 579556 335228 579562
rect 335176 579498 335228 579504
rect 335188 579358 335216 579498
rect 338672 579488 338724 579494
rect 336568 579426 336858 579442
rect 338672 579430 338724 579436
rect 336556 579420 336858 579426
rect 336608 579414 336858 579420
rect 336556 579362 336608 579368
rect 338684 579358 338712 579430
rect 343008 579426 343298 579442
rect 342996 579420 343298 579426
rect 343048 579414 343298 579420
rect 342996 579362 343048 579368
rect 300676 579352 300728 579358
rect 300610 579300 300676 579306
rect 300610 579294 300728 579300
rect 305092 579352 305144 579358
rect 305184 579352 305236 579358
rect 305092 579294 305144 579300
rect 305182 579320 305184 579329
rect 309784 579352 309836 579358
rect 305236 579320 305238 579329
rect 300610 579278 300716 579294
rect 309968 579352 310020 579358
rect 309836 579312 309968 579340
rect 309784 579294 309836 579300
rect 315856 579352 315908 579358
rect 309968 579294 310020 579300
rect 315854 579320 315856 579329
rect 330024 579352 330076 579358
rect 315908 579320 315910 579329
rect 305182 579255 305238 579264
rect 330576 579352 330628 579358
rect 330076 579300 330418 579306
rect 330024 579294 330418 579300
rect 330576 579294 330628 579300
rect 330668 579352 330720 579358
rect 330668 579294 330720 579300
rect 330760 579352 330812 579358
rect 330760 579294 330812 579300
rect 334440 579352 334492 579358
rect 334716 579352 334768 579358
rect 334492 579300 334650 579306
rect 334440 579294 334650 579300
rect 334716 579294 334768 579300
rect 334808 579352 334860 579358
rect 334808 579294 334860 579300
rect 334900 579352 334952 579358
rect 334900 579294 334952 579300
rect 335176 579352 335228 579358
rect 335176 579294 335228 579300
rect 338672 579352 338724 579358
rect 338672 579294 338724 579300
rect 345112 579352 345164 579358
rect 360384 579352 360436 579358
rect 345164 579300 345322 579306
rect 345112 579294 345322 579300
rect 330036 579278 330418 579294
rect 334452 579278 334650 579294
rect 345124 579278 345322 579294
rect 360226 579300 360384 579306
rect 360226 579294 360436 579300
rect 364248 579352 364300 579358
rect 375380 579352 375432 579358
rect 364300 579300 364458 579306
rect 364248 579294 364458 579300
rect 360226 579278 360424 579294
rect 364260 579278 364458 579294
rect 375130 579300 375380 579306
rect 375130 579294 375432 579300
rect 375130 579278 375420 579294
rect 377154 579278 377260 579306
rect 315854 579255 315910 579264
rect 300596 490618 300624 500004
rect 302252 499990 302634 500018
rect 302252 499882 302280 499990
rect 302068 499854 302280 499882
rect 302068 498846 302096 499854
rect 302424 499452 302476 499458
rect 302424 499394 302476 499400
rect 302056 498840 302108 498846
rect 302056 498782 302108 498788
rect 302068 492658 302096 498782
rect 302056 492652 302108 492658
rect 302056 492594 302108 492600
rect 302148 492652 302200 492658
rect 302148 492594 302200 492600
rect 302160 491298 302188 492594
rect 301964 491292 302016 491298
rect 301964 491234 302016 491240
rect 302148 491292 302200 491298
rect 302148 491234 302200 491240
rect 300584 490612 300636 490618
rect 300584 490554 300636 490560
rect 301976 481710 302004 491234
rect 301872 481704 301924 481710
rect 301872 481646 301924 481652
rect 301964 481704 302016 481710
rect 301964 481646 302016 481652
rect 301884 473385 301912 481646
rect 301870 473376 301926 473385
rect 301870 473311 301926 473320
rect 302054 473376 302110 473385
rect 302054 473311 302110 473320
rect 302068 469130 302096 473311
rect 302056 469124 302108 469130
rect 302056 469066 302108 469072
rect 302056 468988 302108 468994
rect 302056 468930 302108 468936
rect 302068 462346 302096 468930
rect 302068 462318 302280 462346
rect 302252 448594 302280 462318
rect 302056 448588 302108 448594
rect 302056 448530 302108 448536
rect 302240 448588 302292 448594
rect 302240 448530 302292 448536
rect 302068 438870 302096 448530
rect 301872 438864 301924 438870
rect 301872 438806 301924 438812
rect 302056 438864 302108 438870
rect 302056 438806 302108 438812
rect 301884 429214 301912 438806
rect 302068 429214 302096 429245
rect 301872 429208 301924 429214
rect 301872 429150 301924 429156
rect 302056 429208 302108 429214
rect 302108 429156 302188 429162
rect 302056 429150 302188 429156
rect 302068 429134 302188 429150
rect 302160 427854 302188 429134
rect 302148 427848 302200 427854
rect 302148 427790 302200 427796
rect 302056 427780 302108 427786
rect 302056 427722 302108 427728
rect 302068 418198 302096 427722
rect 302056 418192 302108 418198
rect 302056 418134 302108 418140
rect 302056 418056 302108 418062
rect 302056 417998 302108 418004
rect 302068 401674 302096 417998
rect 301780 401668 301832 401674
rect 301780 401610 301832 401616
rect 302056 401668 302108 401674
rect 302056 401610 302108 401616
rect 301792 401554 301820 401610
rect 301792 401526 301912 401554
rect 301884 392018 301912 401526
rect 301872 392012 301924 392018
rect 301872 391954 301924 391960
rect 302056 392012 302108 392018
rect 302056 391954 302108 391960
rect 302068 389178 302096 391954
rect 301976 389150 302096 389178
rect 301976 381546 302004 389150
rect 301504 381540 301556 381546
rect 301504 381482 301556 381488
rect 301964 381540 302016 381546
rect 301964 381482 302016 381488
rect 301516 338094 301544 381482
rect 301504 338088 301556 338094
rect 301504 338030 301556 338036
rect 300768 291916 300820 291922
rect 300768 291858 300820 291864
rect 300676 291848 300728 291854
rect 300676 291790 300728 291796
rect 300688 202842 300716 291790
rect 300676 202836 300728 202842
rect 300676 202778 300728 202784
rect 300492 202020 300544 202026
rect 300492 201962 300544 201968
rect 300400 201816 300452 201822
rect 300400 201758 300452 201764
rect 300780 200002 300808 291858
rect 301412 203924 301464 203930
rect 301412 203866 301464 203872
rect 301044 202768 301096 202774
rect 301044 202710 301096 202716
rect 301056 201754 301084 202710
rect 301044 201748 301096 201754
rect 301044 201690 301096 201696
rect 301424 200002 301452 203866
rect 302238 202600 302294 202609
rect 302238 202535 302240 202544
rect 302292 202535 302294 202544
rect 302332 202564 302384 202570
rect 302240 202506 302292 202512
rect 302332 202506 302384 202512
rect 302344 202450 302372 202506
rect 302252 202422 302372 202450
rect 302252 202366 302280 202422
rect 302240 202360 302292 202366
rect 302240 202302 302292 202308
rect 301872 201680 301924 201686
rect 301872 201622 301924 201628
rect 301884 200002 301912 201622
rect 302436 200002 302464 499394
rect 304828 496942 304856 500004
rect 306852 497214 306880 500004
rect 308968 499990 309074 500018
rect 310624 499990 311098 500018
rect 306840 497208 306892 497214
rect 306840 497150 306892 497156
rect 307024 497208 307076 497214
rect 307024 497150 307076 497156
rect 304816 496936 304868 496942
rect 304816 496878 304868 496884
rect 307036 483177 307064 497150
rect 307576 497004 307628 497010
rect 307576 496946 307628 496952
rect 307022 483168 307078 483177
rect 307022 483103 307078 483112
rect 307022 483032 307078 483041
rect 307022 482967 307078 482976
rect 307036 463865 307064 482967
rect 307022 463856 307078 463865
rect 307022 463791 307078 463800
rect 307022 463720 307078 463729
rect 306840 463684 306892 463690
rect 307022 463655 307024 463664
rect 306840 463626 306892 463632
rect 307076 463655 307078 463664
rect 307024 463626 307076 463632
rect 306852 454073 306880 463626
rect 306838 454064 306894 454073
rect 306838 453999 306894 454008
rect 307022 454064 307078 454073
rect 307022 453999 307078 454008
rect 307036 444378 307064 453999
rect 306840 444372 306892 444378
rect 306840 444314 306892 444320
rect 307024 444372 307076 444378
rect 307024 444314 307076 444320
rect 306852 434790 306880 444314
rect 306840 434784 306892 434790
rect 306840 434726 306892 434732
rect 307024 434784 307076 434790
rect 307024 434726 307076 434732
rect 307036 386374 307064 434726
rect 306840 386368 306892 386374
rect 306840 386310 306892 386316
rect 307024 386368 307076 386374
rect 307024 386310 307076 386316
rect 306852 376786 306880 386310
rect 306840 376780 306892 376786
rect 306840 376722 306892 376728
rect 307024 376780 307076 376786
rect 307024 376722 307076 376728
rect 307036 367062 307064 376722
rect 306840 367056 306892 367062
rect 306840 366998 306892 367004
rect 307024 367056 307076 367062
rect 307024 366998 307076 367004
rect 306852 357474 306880 366998
rect 306840 357468 306892 357474
rect 306840 357410 306892 357416
rect 307024 357468 307076 357474
rect 307024 357410 307076 357416
rect 307036 347970 307064 357410
rect 306944 347942 307064 347970
rect 306944 347750 306972 347942
rect 306840 347744 306892 347750
rect 306840 347686 306892 347692
rect 306932 347744 306984 347750
rect 306932 347686 306984 347692
rect 306852 338162 306880 347686
rect 306840 338156 306892 338162
rect 306840 338098 306892 338104
rect 307024 338156 307076 338162
rect 307024 338098 307076 338104
rect 307036 328438 307064 338098
rect 307024 328432 307076 328438
rect 307024 328374 307076 328380
rect 307024 328296 307076 328302
rect 307024 328238 307076 328244
rect 307036 309194 307064 328238
rect 307024 309188 307076 309194
rect 307024 309130 307076 309136
rect 307116 309120 307168 309126
rect 307116 309062 307168 309068
rect 307128 307834 307156 309062
rect 307116 307828 307168 307834
rect 307116 307770 307168 307776
rect 307208 307828 307260 307834
rect 307208 307770 307260 307776
rect 307220 299538 307248 307770
rect 307024 299532 307076 299538
rect 307024 299474 307076 299480
rect 307208 299532 307260 299538
rect 307208 299474 307260 299480
rect 307036 270570 307064 299474
rect 307024 270564 307076 270570
rect 307024 270506 307076 270512
rect 306932 270496 306984 270502
rect 306932 270438 306984 270444
rect 306944 269074 306972 270438
rect 306748 269068 306800 269074
rect 306748 269010 306800 269016
rect 306932 269068 306984 269074
rect 306932 269010 306984 269016
rect 306760 259486 306788 269010
rect 306748 259480 306800 259486
rect 306748 259422 306800 259428
rect 307024 259480 307076 259486
rect 307024 259422 307076 259428
rect 307036 251530 307064 259422
rect 307024 251524 307076 251530
rect 307024 251466 307076 251472
rect 307024 251388 307076 251394
rect 307024 251330 307076 251336
rect 307036 251002 307064 251330
rect 307036 250974 307248 251002
rect 307220 241602 307248 250974
rect 307024 241596 307076 241602
rect 307024 241538 307076 241544
rect 307208 241596 307260 241602
rect 307208 241538 307260 241544
rect 307036 240122 307064 241538
rect 306944 240094 307064 240122
rect 306944 231878 306972 240094
rect 306932 231872 306984 231878
rect 306932 231814 306984 231820
rect 307024 231804 307076 231810
rect 307024 231746 307076 231752
rect 307036 230518 307064 231746
rect 306932 230512 306984 230518
rect 306932 230454 306984 230460
rect 307024 230512 307076 230518
rect 307024 230454 307076 230460
rect 306944 224890 306972 230454
rect 306944 224862 307156 224890
rect 307128 222154 307156 224862
rect 307024 222148 307076 222154
rect 307024 222090 307076 222096
rect 307116 222148 307168 222154
rect 307116 222090 307168 222096
rect 307036 212566 307064 222090
rect 307024 212560 307076 212566
rect 307024 212502 307076 212508
rect 307208 212560 307260 212566
rect 307208 212502 307260 212508
rect 303896 211132 303948 211138
rect 303896 211074 303948 211080
rect 302884 203380 302936 203386
rect 302884 203322 302936 203328
rect 302896 200002 302924 203322
rect 302976 202564 303028 202570
rect 302976 202506 303028 202512
rect 284128 199974 284188 200002
rect 285476 199974 285628 200002
rect 285936 199974 286272 200002
rect 286764 199974 287008 200002
rect 287224 199974 287560 200002
rect 287684 199974 288020 200002
rect 288512 199974 288848 200002
rect 288972 199974 289308 200002
rect 289432 199974 289676 200002
rect 290260 199974 290596 200002
rect 290720 199974 291056 200002
rect 291180 199974 291424 200002
rect 292008 199974 292344 200002
rect 292468 199974 292528 200002
rect 292928 199974 293172 200002
rect 293756 199974 293816 200002
rect 294216 199974 294460 200002
rect 294584 199974 294920 200002
rect 295504 199974 295840 200002
rect 295964 199974 296208 200002
rect 296332 199974 296576 200002
rect 297252 199974 297312 200002
rect 297712 199974 297956 200002
rect 298080 199974 298416 200002
rect 299000 199974 299244 200002
rect 299368 199974 299428 200002
rect 299828 199974 300164 200002
rect 300748 199974 300808 200002
rect 301116 199974 301452 200002
rect 301576 199974 301912 200002
rect 302404 199974 302464 200002
rect 302864 199974 302924 200002
rect 302988 200002 303016 202506
rect 303908 202178 303936 211074
rect 306656 203992 306708 203998
rect 306656 203934 306708 203940
rect 305000 202700 305052 202706
rect 305000 202642 305052 202648
rect 303908 202150 304488 202178
rect 303896 202088 303948 202094
rect 303896 202030 303948 202036
rect 304262 202056 304318 202065
rect 303908 200002 303936 202030
rect 304262 201991 304318 202000
rect 304276 201958 304304 201991
rect 304264 201952 304316 201958
rect 304264 201894 304316 201900
rect 304460 200002 304488 202150
rect 305012 200002 305040 202642
rect 305644 202632 305696 202638
rect 305644 202574 305696 202580
rect 305552 202360 305604 202366
rect 305552 202302 305604 202308
rect 305564 201890 305592 202302
rect 305552 201884 305604 201890
rect 305552 201826 305604 201832
rect 305656 200002 305684 202574
rect 306668 200002 306696 203934
rect 307116 202836 307168 202842
rect 307116 202778 307168 202784
rect 306932 202700 306984 202706
rect 306932 202642 306984 202648
rect 306944 202434 306972 202642
rect 306932 202428 306984 202434
rect 306932 202370 306984 202376
rect 307024 202428 307076 202434
rect 307024 202370 307076 202376
rect 306932 202088 306984 202094
rect 306932 202030 306984 202036
rect 306944 201550 306972 202030
rect 306932 201544 306984 201550
rect 306932 201486 306984 201492
rect 307036 200002 307064 202370
rect 307128 201822 307156 202778
rect 307220 202774 307248 212502
rect 307208 202768 307260 202774
rect 307208 202710 307260 202716
rect 307208 202632 307260 202638
rect 307206 202600 307208 202609
rect 307260 202600 307262 202609
rect 307206 202535 307262 202544
rect 307300 202564 307352 202570
rect 307300 202506 307352 202512
rect 307312 202065 307340 202506
rect 307588 202434 307616 496946
rect 308864 492788 308916 492794
rect 308864 492730 308916 492736
rect 308876 486418 308904 492730
rect 308784 486390 308904 486418
rect 308784 481642 308812 486390
rect 308772 481636 308824 481642
rect 308772 481578 308824 481584
rect 308864 481636 308916 481642
rect 308864 481578 308916 481584
rect 308876 473414 308904 481578
rect 308864 473408 308916 473414
rect 308864 473350 308916 473356
rect 308772 473340 308824 473346
rect 308772 473282 308824 473288
rect 308784 472002 308812 473282
rect 308784 471974 308904 472002
rect 308876 452554 308904 471974
rect 308784 452526 308904 452554
rect 308784 443018 308812 452526
rect 308772 443012 308824 443018
rect 308772 442954 308824 442960
rect 308864 443012 308916 443018
rect 308864 442954 308916 442960
rect 308876 433242 308904 442954
rect 308784 433214 308904 433242
rect 308784 423706 308812 433214
rect 308772 423700 308824 423706
rect 308772 423642 308824 423648
rect 308864 423700 308916 423706
rect 308864 423642 308916 423648
rect 308876 413930 308904 423642
rect 308784 413902 308904 413930
rect 308784 404394 308812 413902
rect 308772 404388 308824 404394
rect 308772 404330 308824 404336
rect 308864 404388 308916 404394
rect 308864 404330 308916 404336
rect 308876 394602 308904 404330
rect 308588 394596 308640 394602
rect 308588 394538 308640 394544
rect 308864 394596 308916 394602
rect 308864 394538 308916 394544
rect 308600 376786 308628 394538
rect 308588 376780 308640 376786
rect 308588 376722 308640 376728
rect 308680 376780 308732 376786
rect 308680 376722 308732 376728
rect 308692 365838 308720 376722
rect 308680 365832 308732 365838
rect 308680 365774 308732 365780
rect 308864 365832 308916 365838
rect 308864 365774 308916 365780
rect 308876 365702 308904 365774
rect 308680 365696 308732 365702
rect 308680 365638 308732 365644
rect 308864 365696 308916 365702
rect 308864 365638 308916 365644
rect 308692 357474 308720 365638
rect 308680 357468 308732 357474
rect 308680 357410 308732 357416
rect 308864 357400 308916 357406
rect 308864 357342 308916 357348
rect 308876 351234 308904 357342
rect 308692 351206 308904 351234
rect 308692 346458 308720 351206
rect 308680 346452 308732 346458
rect 308680 346394 308732 346400
rect 308772 346452 308824 346458
rect 308772 346394 308824 346400
rect 308784 338162 308812 346394
rect 308772 338156 308824 338162
rect 308772 338098 308824 338104
rect 308864 338020 308916 338026
rect 308864 337962 308916 337968
rect 308876 336682 308904 337962
rect 308784 336654 308904 336682
rect 308784 327214 308812 336654
rect 308772 327208 308824 327214
rect 308772 327150 308824 327156
rect 308864 327140 308916 327146
rect 308864 327082 308916 327088
rect 308876 317370 308904 327082
rect 308784 317342 308904 317370
rect 308784 299538 308812 317342
rect 308680 299532 308732 299538
rect 308680 299474 308732 299480
rect 308772 299532 308824 299538
rect 308772 299474 308824 299480
rect 308692 292602 308720 299474
rect 308680 292596 308732 292602
rect 308680 292538 308732 292544
rect 308864 292596 308916 292602
rect 308864 292538 308916 292544
rect 308876 283626 308904 292538
rect 308588 283620 308640 283626
rect 308588 283562 308640 283568
rect 308864 283620 308916 283626
rect 308864 283562 308916 283568
rect 308600 278798 308628 283562
rect 308588 278792 308640 278798
rect 308588 278734 308640 278740
rect 308680 278792 308732 278798
rect 308680 278734 308732 278740
rect 308692 269142 308720 278734
rect 308680 269136 308732 269142
rect 308680 269078 308732 269084
rect 308864 269136 308916 269142
rect 308864 269078 308916 269084
rect 308876 251433 308904 269078
rect 308862 251424 308918 251433
rect 308862 251359 308918 251368
rect 308862 251288 308918 251297
rect 308862 251223 308918 251232
rect 308876 245410 308904 251223
rect 308588 245404 308640 245410
rect 308588 245346 308640 245352
rect 308864 245404 308916 245410
rect 308864 245346 308916 245352
rect 308600 235346 308628 245346
rect 308588 235340 308640 235346
rect 308588 235282 308640 235288
rect 308772 235340 308824 235346
rect 308772 235282 308824 235288
rect 308784 230466 308812 235282
rect 308692 230438 308812 230466
rect 308692 222222 308720 230438
rect 308680 222216 308732 222222
rect 308680 222158 308732 222164
rect 308772 222148 308824 222154
rect 308772 222090 308824 222096
rect 308784 220862 308812 222090
rect 308680 220856 308732 220862
rect 308680 220798 308732 220804
rect 308772 220856 308824 220862
rect 308772 220798 308824 220804
rect 308692 216034 308720 220798
rect 308312 216028 308364 216034
rect 308312 215970 308364 215976
rect 308680 216028 308732 216034
rect 308680 215970 308732 215976
rect 308324 212378 308352 215970
rect 308324 212350 308444 212378
rect 308416 205630 308444 212350
rect 308404 205624 308456 205630
rect 308404 205566 308456 205572
rect 308588 205624 308640 205630
rect 308588 205566 308640 205572
rect 308404 204060 308456 204066
rect 308404 204002 308456 204008
rect 307576 202428 307628 202434
rect 307576 202370 307628 202376
rect 307298 202056 307354 202065
rect 307298 201991 307354 202000
rect 307116 201816 307168 201822
rect 307116 201758 307168 201764
rect 307300 201612 307352 201618
rect 307300 201554 307352 201560
rect 302988 199974 303324 200002
rect 303908 199974 304152 200002
rect 304460 199974 304612 200002
rect 305012 199974 305072 200002
rect 305656 199974 305900 200002
rect 306360 199974 306696 200002
rect 306820 199974 307064 200002
rect 307312 200002 307340 201554
rect 308416 200002 308444 204002
rect 308600 202858 308628 205566
rect 308968 203182 308996 499990
rect 310520 499044 310572 499050
rect 310520 498986 310572 498992
rect 309048 498908 309100 498914
rect 309048 498850 309100 498856
rect 309060 492794 309088 498850
rect 309324 496936 309376 496942
rect 309324 496878 309376 496884
rect 309048 492788 309100 492794
rect 309048 492730 309100 492736
rect 308956 203176 309008 203182
rect 308956 203118 309008 203124
rect 308600 202830 308812 202858
rect 308784 200258 308812 202830
rect 308542 200252 308594 200258
rect 308542 200194 308594 200200
rect 308772 200252 308824 200258
rect 308772 200194 308824 200200
rect 307312 199974 307648 200002
rect 308108 199974 308444 200002
rect 308554 199988 308582 200194
rect 309336 200002 309364 496878
rect 310428 202768 310480 202774
rect 310428 202710 310480 202716
rect 309508 202632 309560 202638
rect 309508 202574 309560 202580
rect 309520 200002 309548 202574
rect 310440 200002 310468 202710
rect 310532 202434 310560 498986
rect 310624 347070 310652 499990
rect 311900 498976 311952 498982
rect 311900 498918 311952 498924
rect 310612 347064 310664 347070
rect 310612 347006 310664 347012
rect 311912 202842 311940 498918
rect 313292 497894 313320 500004
rect 315040 499990 315330 500018
rect 313280 497888 313332 497894
rect 313280 497830 313332 497836
rect 315040 497010 315068 499990
rect 317328 498976 317380 498982
rect 317328 498918 317380 498924
rect 315028 497004 315080 497010
rect 315028 496946 315080 496952
rect 315304 497004 315356 497010
rect 315304 496946 315356 496952
rect 311992 210452 312044 210458
rect 311992 210394 312044 210400
rect 311900 202836 311952 202842
rect 311900 202778 311952 202784
rect 311164 202632 311216 202638
rect 311164 202574 311216 202580
rect 310520 202428 310572 202434
rect 310520 202370 310572 202376
rect 311176 200002 311204 202574
rect 311256 202428 311308 202434
rect 311256 202370 311308 202376
rect 311348 202428 311400 202434
rect 311348 202370 311400 202376
rect 309336 199974 309396 200002
rect 309520 199974 309856 200002
rect 310316 199974 310468 200002
rect 311144 199974 311204 200002
rect 311268 200002 311296 202370
rect 311360 201754 311388 202370
rect 311348 201748 311400 201754
rect 311348 201690 311400 201696
rect 312004 200002 312032 210394
rect 313556 204196 313608 204202
rect 313556 204138 313608 204144
rect 312544 202836 312596 202842
rect 312544 202778 312596 202784
rect 312636 202836 312688 202842
rect 312636 202778 312688 202784
rect 311268 199974 311604 200002
rect 311972 199974 312032 200002
rect 312556 200002 312584 202778
rect 312648 201686 312676 202778
rect 312636 201680 312688 201686
rect 312636 201622 312688 201628
rect 313568 200002 313596 204138
rect 314936 204128 314988 204134
rect 314936 204070 314988 204076
rect 313648 201816 313700 201822
rect 313648 201758 313700 201764
rect 312556 199974 312892 200002
rect 313352 199974 313596 200002
rect 313660 200002 313688 201758
rect 314948 200002 314976 204070
rect 315212 203244 315264 203250
rect 315212 203186 315264 203192
rect 315224 200002 315252 203186
rect 315316 202502 315344 496946
rect 317340 204762 317368 498918
rect 317524 497146 317552 500004
rect 318708 497888 318760 497894
rect 318708 497830 318760 497836
rect 317512 497140 317564 497146
rect 317512 497082 317564 497088
rect 317064 204734 317368 204762
rect 315304 202496 315356 202502
rect 315304 202438 315356 202444
rect 315304 202088 315356 202094
rect 315304 202030 315356 202036
rect 313660 199974 313720 200002
rect 314640 199974 314976 200002
rect 315100 199974 315252 200002
rect 315316 200002 315344 202030
rect 315580 201952 315632 201958
rect 315580 201894 315632 201900
rect 315592 200002 315620 201894
rect 317064 200002 317092 204734
rect 317144 202020 317196 202026
rect 317144 201962 317196 201968
rect 315316 199974 315468 200002
rect 315592 199974 315928 200002
rect 316756 199974 317092 200002
rect 317156 200002 317184 201962
rect 318720 200002 318748 497830
rect 319732 497826 319760 500004
rect 321468 499044 321520 499050
rect 321468 498986 321520 498992
rect 319720 497820 319772 497826
rect 319720 497762 319772 497768
rect 320088 497820 320140 497826
rect 320088 497762 320140 497768
rect 318892 340400 318944 340406
rect 318812 340348 318892 340354
rect 318812 340342 318944 340348
rect 318812 340338 318932 340342
rect 318800 340332 318932 340338
rect 318852 340326 318932 340332
rect 318800 340274 318852 340280
rect 319168 204264 319220 204270
rect 319168 204206 319220 204212
rect 319180 202842 319208 204206
rect 320100 202842 320128 497762
rect 319168 202836 319220 202842
rect 319168 202778 319220 202784
rect 319260 202836 319312 202842
rect 319260 202778 319312 202784
rect 320088 202836 320140 202842
rect 320088 202778 320140 202784
rect 319272 200002 319300 202778
rect 320640 202700 320692 202706
rect 320640 202642 320692 202648
rect 320548 202020 320600 202026
rect 320548 201962 320600 201968
rect 320560 200002 320588 201962
rect 317156 199974 317216 200002
rect 318504 199974 318748 200002
rect 318964 199974 319300 200002
rect 320252 199974 320588 200002
rect 320652 200002 320680 202642
rect 321480 202026 321508 498986
rect 321756 497078 321784 500004
rect 321744 497072 321796 497078
rect 321744 497014 321796 497020
rect 323964 497010 323992 500004
rect 325712 499990 326002 500018
rect 324228 499112 324280 499118
rect 324228 499054 324280 499060
rect 323952 497004 324004 497010
rect 323952 496946 324004 496952
rect 322848 291984 322900 291990
rect 322848 291926 322900 291932
rect 321744 203176 321796 203182
rect 321744 203118 321796 203124
rect 321468 202020 321520 202026
rect 321468 201962 321520 201968
rect 321756 200002 321784 203118
rect 322860 200138 322888 291926
rect 324044 202020 324096 202026
rect 324044 201962 324096 201968
rect 322676 200110 322888 200138
rect 322676 200002 322704 200110
rect 324056 200002 324084 201962
rect 324240 200002 324268 499054
rect 324964 496936 325016 496942
rect 324964 496878 325016 496884
rect 324976 202026 325004 496878
rect 325148 203312 325200 203318
rect 325148 203254 325200 203260
rect 324964 202020 325016 202026
rect 324964 201962 325016 201968
rect 320652 199974 320712 200002
rect 321756 199974 322000 200002
rect 322460 199974 322704 200002
rect 323748 199974 324084 200002
rect 324208 199974 324268 200002
rect 325160 200002 325188 203254
rect 325712 202570 325740 499990
rect 328196 496942 328224 500004
rect 329852 499990 330234 500018
rect 331232 499990 332442 500018
rect 328184 496936 328236 496942
rect 328184 496878 328236 496884
rect 329852 337482 329880 499990
rect 331128 340400 331180 340406
rect 331128 340342 331180 340348
rect 331140 340270 331168 340342
rect 331128 340264 331180 340270
rect 331128 340206 331180 340212
rect 329840 337476 329892 337482
rect 329840 337418 329892 337424
rect 331232 203386 331260 499990
rect 334452 497962 334480 500004
rect 334440 497956 334492 497962
rect 334440 497898 334492 497904
rect 336004 497956 336056 497962
rect 336004 497898 336056 497904
rect 334624 497140 334676 497146
rect 334624 497082 334676 497088
rect 331864 496936 331916 496942
rect 331864 496878 331916 496884
rect 331220 203380 331272 203386
rect 331220 203322 331272 203328
rect 331876 202638 331904 496878
rect 333888 362976 333940 362982
rect 333888 362918 333940 362924
rect 333796 347064 333848 347070
rect 333796 347006 333848 347012
rect 333244 340468 333296 340474
rect 333244 340410 333296 340416
rect 333256 340270 333284 340410
rect 333244 340264 333296 340270
rect 333244 340206 333296 340212
rect 331864 202632 331916 202638
rect 331864 202574 331916 202580
rect 325700 202564 325752 202570
rect 325700 202506 325752 202512
rect 333152 202496 333204 202502
rect 333152 202438 333204 202444
rect 325700 202428 325752 202434
rect 325700 202370 325752 202376
rect 332508 202428 332560 202434
rect 332508 202370 332560 202376
rect 325712 200002 325740 202370
rect 332520 200002 332548 202370
rect 333164 200002 333192 202438
rect 333808 200138 333836 347006
rect 333900 202502 333928 362918
rect 333888 202496 333940 202502
rect 333888 202438 333940 202444
rect 334636 202026 334664 497082
rect 336016 203250 336044 497898
rect 336660 496942 336688 500004
rect 338868 498030 338896 500004
rect 338856 498024 338908 498030
rect 338856 497966 338908 497972
rect 336648 496936 336700 496942
rect 336648 496878 336700 496884
rect 340892 203454 340920 500004
rect 343100 497146 343128 500004
rect 345124 497350 345152 500004
rect 347332 498098 347360 500004
rect 347320 498092 347372 498098
rect 347320 498034 347372 498040
rect 349356 497962 349384 500004
rect 349344 497956 349396 497962
rect 349344 497898 349396 497904
rect 345112 497344 345164 497350
rect 345112 497286 345164 497292
rect 351564 497282 351592 500004
rect 353312 499990 353602 500018
rect 351552 497276 351604 497282
rect 351552 497218 351604 497224
rect 343088 497140 343140 497146
rect 343088 497082 343140 497088
rect 344928 385756 344980 385762
rect 344928 385698 344980 385704
rect 343548 385212 343600 385218
rect 343548 385154 343600 385160
rect 342168 347336 342220 347342
rect 342168 347278 342220 347284
rect 340880 203448 340932 203454
rect 340880 203390 340932 203396
rect 336004 203244 336056 203250
rect 336004 203186 336056 203192
rect 342076 202632 342128 202638
rect 342076 202574 342128 202580
rect 341432 202496 341484 202502
rect 341432 202438 341484 202444
rect 334624 202020 334676 202026
rect 334624 201962 334676 201968
rect 333532 200110 333836 200138
rect 333532 200002 333560 200110
rect 341444 200002 341472 202438
rect 342088 200002 342116 202574
rect 342180 202502 342208 347278
rect 343560 202502 343588 385154
rect 344008 202700 344060 202706
rect 344008 202642 344060 202648
rect 342168 202496 342220 202502
rect 342168 202438 342220 202444
rect 343180 202496 343232 202502
rect 343180 202438 343232 202444
rect 343548 202496 343600 202502
rect 343548 202438 343600 202444
rect 343192 200002 343220 202438
rect 344020 200002 344048 202642
rect 344940 200002 344968 385698
rect 349068 385552 349120 385558
rect 349068 385494 349120 385500
rect 347688 385280 347740 385286
rect 347688 385222 347740 385228
rect 347596 369912 347648 369918
rect 347596 369854 347648 369860
rect 347608 202502 347636 369854
rect 346676 202496 346728 202502
rect 346676 202438 346728 202444
rect 347596 202496 347648 202502
rect 347596 202438 347648 202444
rect 345756 202156 345808 202162
rect 345756 202098 345808 202104
rect 345768 200002 345796 202098
rect 346688 200002 346716 202438
rect 347700 200138 347728 385222
rect 348332 202632 348384 202638
rect 348332 202574 348384 202580
rect 347516 200110 347728 200138
rect 347516 200002 347544 200110
rect 348344 200002 348372 202574
rect 349080 200002 349108 385494
rect 353208 385416 353260 385422
rect 353208 385358 353260 385364
rect 351828 376780 351880 376786
rect 351828 376722 351880 376728
rect 350540 347404 350592 347410
rect 350540 347346 350592 347352
rect 350552 338162 350580 347346
rect 350264 338156 350316 338162
rect 350264 338098 350316 338104
rect 350540 338156 350592 338162
rect 350540 338098 350592 338104
rect 350276 331242 350304 338098
rect 350276 331214 350488 331242
rect 350460 202706 350488 331214
rect 351840 202842 351868 376722
rect 353220 202842 353248 385358
rect 353312 203522 353340 499990
rect 355796 497894 355824 500004
rect 355784 497888 355836 497894
rect 355784 497830 355836 497836
rect 358004 497826 358032 500004
rect 357992 497820 358044 497826
rect 357992 497762 358044 497768
rect 360028 497554 360056 500004
rect 360016 497548 360068 497554
rect 360016 497490 360068 497496
rect 362236 497214 362264 500004
rect 362224 497208 362276 497214
rect 362224 497150 362276 497156
rect 364260 496874 364288 500004
rect 366468 497418 366496 500004
rect 368492 497758 368520 500004
rect 369872 499990 370714 500018
rect 368480 497752 368532 497758
rect 368480 497694 368532 497700
rect 366456 497412 366508 497418
rect 366456 497354 366508 497360
rect 364248 496868 364300 496874
rect 364248 496810 364300 496816
rect 365628 385620 365680 385626
rect 365628 385562 365680 385568
rect 355876 385484 355928 385490
rect 355876 385426 355928 385432
rect 354588 353320 354640 353326
rect 354588 353262 354640 353268
rect 354496 347200 354548 347206
rect 354496 347142 354548 347148
rect 353300 203516 353352 203522
rect 353300 203458 353352 203464
rect 351000 202836 351052 202842
rect 351000 202778 351052 202784
rect 351828 202836 351880 202842
rect 351828 202778 351880 202784
rect 352748 202836 352800 202842
rect 352748 202778 352800 202784
rect 353208 202836 353260 202842
rect 353208 202778 353260 202784
rect 353300 202836 353352 202842
rect 353300 202778 353352 202784
rect 349988 202700 350040 202706
rect 349988 202642 350040 202648
rect 350448 202700 350500 202706
rect 350448 202642 350500 202648
rect 350000 200002 350028 202642
rect 351012 200002 351040 202778
rect 351736 202700 351788 202706
rect 351736 202642 351788 202648
rect 351748 200002 351776 202642
rect 352760 200002 352788 202778
rect 353312 202706 353340 202778
rect 353300 202700 353352 202706
rect 353300 202642 353352 202648
rect 353484 202632 353536 202638
rect 353484 202574 353536 202580
rect 353496 202162 353524 202574
rect 353484 202156 353536 202162
rect 353484 202098 353536 202104
rect 353576 202156 353628 202162
rect 353576 202098 353628 202104
rect 353588 200002 353616 202098
rect 354508 200002 354536 347142
rect 354600 202162 354628 353262
rect 354588 202156 354640 202162
rect 354588 202098 354640 202104
rect 355324 201544 355376 201550
rect 355324 201486 355376 201492
rect 355336 200002 355364 201486
rect 325160 199974 325496 200002
rect 325712 199974 325956 200002
rect 332488 199974 332548 200002
rect 332856 199974 333192 200002
rect 333316 199974 333560 200002
rect 341136 199974 341472 200002
rect 342056 199974 342116 200002
rect 342884 199974 343220 200002
rect 343712 199974 344048 200002
rect 344632 199974 344968 200002
rect 345460 199974 345796 200002
rect 346380 199974 346716 200002
rect 347208 199974 347544 200002
rect 348128 199974 348372 200002
rect 348956 199974 349108 200002
rect 349876 199974 350028 200002
rect 350704 199974 351040 200002
rect 351624 199974 351776 200002
rect 352452 199974 352788 200002
rect 353280 199974 353616 200002
rect 354200 199974 354536 200002
rect 355028 199974 355364 200002
rect 355888 200002 355916 385426
rect 357348 385348 357400 385354
rect 357348 385290 357400 385296
rect 355968 385144 356020 385150
rect 355968 385086 356020 385092
rect 355980 201550 356008 385086
rect 355968 201544 356020 201550
rect 355968 201486 356020 201492
rect 357360 200138 357388 385290
rect 364248 374060 364300 374066
rect 364248 374002 364300 374008
rect 360108 347676 360160 347682
rect 360108 347618 360160 347624
rect 358728 347608 358780 347614
rect 358728 347550 358780 347556
rect 357440 340400 357492 340406
rect 357440 340342 357492 340348
rect 357452 340270 357480 340342
rect 357440 340264 357492 340270
rect 357440 340206 357492 340212
rect 357900 202088 357952 202094
rect 357900 202030 357952 202036
rect 357084 200110 357388 200138
rect 357084 200002 357112 200110
rect 357912 200002 357940 202030
rect 358740 200002 358768 347550
rect 360120 201550 360148 347618
rect 362868 347540 362920 347546
rect 362868 347482 362920 347488
rect 362776 347472 362828 347478
rect 362776 347414 362828 347420
rect 361488 347268 361540 347274
rect 361488 347210 361540 347216
rect 361396 347132 361448 347138
rect 361396 347074 361448 347080
rect 361408 201550 361436 347074
rect 359648 201544 359700 201550
rect 359648 201486 359700 201492
rect 360108 201544 360160 201550
rect 360108 201486 360160 201492
rect 360568 201544 360620 201550
rect 360568 201486 360620 201492
rect 361396 201544 361448 201550
rect 361396 201486 361448 201492
rect 359660 200002 359688 201486
rect 360580 200002 360608 201486
rect 361500 200138 361528 347210
rect 362224 340400 362276 340406
rect 362224 340342 362276 340348
rect 362236 340270 362264 340342
rect 362224 340264 362276 340270
rect 362224 340206 362276 340212
rect 362788 201550 362816 347414
rect 362316 201544 362368 201550
rect 362316 201486 362368 201492
rect 362776 201544 362828 201550
rect 362776 201486 362828 201492
rect 361408 200110 361528 200138
rect 361408 200002 361436 200110
rect 362328 200002 362356 201486
rect 362880 200002 362908 347482
rect 364260 200138 364288 374002
rect 365536 347744 365588 347750
rect 365536 347686 365588 347692
rect 365548 202162 365576 347686
rect 364892 202156 364944 202162
rect 364892 202098 364944 202104
rect 365536 202156 365588 202162
rect 365536 202098 365588 202104
rect 364076 200110 364288 200138
rect 364076 200002 364104 200110
rect 364904 200002 364932 202098
rect 365640 202042 365668 385562
rect 367008 385076 367060 385082
rect 367008 385018 367060 385024
rect 367020 202162 367048 385018
rect 369872 203658 369900 499990
rect 372724 497486 372752 500004
rect 374932 497622 374960 500004
rect 375288 498840 375340 498846
rect 375288 498782 375340 498788
rect 374920 497616 374972 497622
rect 374920 497558 374972 497564
rect 372712 497480 372764 497486
rect 372712 497422 372764 497428
rect 369860 203652 369912 203658
rect 369860 203594 369912 203600
rect 375300 202230 375328 498782
rect 377140 497690 377168 500004
rect 377128 497684 377180 497690
rect 377128 497626 377180 497632
rect 377232 204066 377260 579278
rect 377220 204060 377272 204066
rect 377220 204002 377272 204008
rect 375656 202768 375708 202774
rect 375656 202710 375708 202716
rect 375748 202768 375800 202774
rect 375748 202710 375800 202716
rect 375668 202366 375696 202710
rect 375656 202360 375708 202366
rect 375656 202302 375708 202308
rect 374368 202224 374420 202230
rect 374368 202166 374420 202172
rect 374460 202224 374512 202230
rect 374460 202166 374512 202172
rect 375288 202224 375340 202230
rect 375288 202166 375340 202172
rect 366180 202156 366232 202162
rect 366180 202098 366232 202104
rect 367008 202156 367060 202162
rect 367008 202098 367060 202104
rect 365364 202014 365668 202042
rect 365364 200002 365392 202014
rect 366192 200002 366220 202098
rect 366916 202020 366968 202026
rect 366916 201962 366968 201968
rect 366928 200002 366956 201962
rect 374380 201958 374408 202166
rect 374368 201952 374420 201958
rect 374368 201894 374420 201900
rect 374472 200002 374500 202166
rect 375760 200002 375788 202710
rect 377324 202366 377352 582490
rect 377496 582480 377548 582486
rect 377496 582422 377548 582428
rect 377402 572112 377458 572121
rect 377402 572047 377458 572056
rect 377416 500478 377444 572047
rect 377404 500472 377456 500478
rect 377404 500414 377456 500420
rect 377508 498914 377536 582422
rect 377600 498982 377628 582558
rect 378968 579352 379020 579358
rect 378968 579294 379020 579300
rect 378138 569732 378194 569741
rect 378138 569667 378194 569676
rect 377678 519208 377734 519217
rect 377678 519143 377734 519152
rect 377692 500886 377720 519143
rect 377680 500880 377732 500886
rect 377680 500822 377732 500828
rect 377588 498976 377640 498982
rect 377588 498918 377640 498924
rect 377496 498908 377548 498914
rect 377496 498850 377548 498856
rect 378152 204202 378180 569667
rect 378230 566468 378286 566477
rect 378230 566403 378286 566412
rect 378244 204950 378272 566403
rect 378322 563476 378378 563485
rect 378322 563411 378378 563420
rect 378336 205018 378364 563411
rect 378414 559600 378470 559609
rect 378414 559535 378470 559544
rect 378324 205012 378376 205018
rect 378324 204954 378376 204960
rect 378232 204944 378284 204950
rect 378232 204886 378284 204892
rect 378140 204196 378192 204202
rect 378140 204138 378192 204144
rect 377312 202360 377364 202366
rect 377312 202302 377364 202308
rect 378428 202201 378456 559535
rect 378598 556608 378654 556617
rect 378598 556543 378654 556552
rect 378506 521792 378562 521801
rect 378506 521727 378562 521736
rect 378520 202298 378548 521727
rect 378612 291922 378640 556543
rect 378784 556232 378836 556238
rect 378784 556174 378836 556180
rect 378690 550760 378746 550769
rect 378690 550695 378746 550704
rect 378704 291990 378732 550695
rect 378692 291984 378744 291990
rect 378692 291926 378744 291932
rect 378600 291916 378652 291922
rect 378600 291858 378652 291864
rect 378796 202774 378824 556174
rect 378874 547088 378930 547097
rect 378874 547023 378930 547032
rect 378888 291854 378916 547023
rect 378980 499050 379008 579294
rect 379072 499118 379100 582626
rect 380530 575512 380586 575521
rect 380530 575447 380586 575456
rect 379518 553480 379574 553489
rect 379518 553415 379574 553424
rect 379060 499112 379112 499118
rect 379060 499054 379112 499060
rect 378968 499044 379020 499050
rect 378968 498986 379020 498992
rect 378876 291848 378928 291854
rect 378876 291790 378928 291796
rect 379532 203930 379560 553415
rect 379610 543824 379666 543833
rect 379610 543759 379666 543768
rect 379520 203924 379572 203930
rect 379520 203866 379572 203872
rect 379624 203726 379652 543759
rect 380346 541104 380402 541113
rect 380346 541039 380402 541048
rect 379702 537568 379758 537577
rect 379702 537503 379758 537512
rect 379612 203720 379664 203726
rect 379612 203662 379664 203668
rect 378784 202768 378836 202774
rect 378784 202710 378836 202716
rect 378508 202292 378560 202298
rect 378508 202234 378560 202240
rect 379716 202230 379744 537503
rect 379794 534576 379850 534585
rect 379794 534511 379850 534520
rect 379808 203794 379836 534511
rect 379886 531448 379942 531457
rect 379886 531383 379942 531392
rect 379796 203788 379848 203794
rect 379796 203730 379848 203736
rect 379900 203590 379928 531383
rect 379978 525056 380034 525065
rect 379978 524991 380034 525000
rect 379888 203584 379940 203590
rect 379888 203526 379940 203532
rect 379704 202224 379756 202230
rect 378414 202192 378470 202201
rect 376484 202156 376536 202162
rect 379704 202166 379756 202172
rect 378414 202127 378470 202136
rect 376484 202098 376536 202104
rect 376496 200002 376524 202098
rect 379992 201958 380020 524991
rect 380070 515536 380126 515545
rect 380070 515471 380126 515480
rect 380084 204270 380112 515471
rect 380162 512544 380218 512553
rect 380162 512479 380218 512488
rect 380072 204264 380124 204270
rect 380072 204206 380124 204212
rect 380176 204134 380204 512479
rect 380254 509552 380310 509561
rect 380254 509487 380310 509496
rect 380164 204128 380216 204134
rect 380164 204070 380216 204076
rect 380268 203862 380296 509487
rect 380360 506666 380388 541039
rect 380438 528728 380494 528737
rect 380438 528663 380494 528672
rect 380348 506660 380400 506666
rect 380348 506602 380400 506608
rect 380346 506560 380402 506569
rect 380346 506495 380402 506504
rect 380360 500954 380388 506495
rect 380348 500948 380400 500954
rect 380348 500890 380400 500896
rect 380452 337414 380480 528663
rect 380544 407862 380572 575447
rect 418804 556300 418856 556306
rect 418804 556242 418856 556248
rect 380624 506660 380676 506666
rect 380624 506602 380676 506608
rect 380636 500410 380664 506602
rect 380714 503024 380770 503033
rect 380714 502959 380770 502968
rect 380624 500404 380676 500410
rect 380624 500346 380676 500352
rect 380532 407856 380584 407862
rect 380532 407798 380584 407804
rect 380440 337408 380492 337414
rect 380440 337350 380492 337356
rect 380728 203998 380756 502959
rect 416780 407788 416832 407794
rect 416780 407730 416832 407736
rect 411260 407176 411312 407182
rect 411260 407118 411312 407124
rect 402980 406496 403032 406502
rect 402980 406438 403032 406444
rect 402992 393310 403020 406438
rect 402980 393304 403032 393310
rect 402980 393246 403032 393252
rect 403900 393304 403952 393310
rect 403900 393246 403952 393252
rect 388260 385688 388312 385694
rect 388260 385630 388312 385636
rect 385868 385552 385920 385558
rect 385868 385494 385920 385500
rect 385880 383316 385908 385494
rect 388272 383316 388300 385630
rect 392860 385620 392912 385626
rect 392860 385562 392912 385568
rect 390468 385076 390520 385082
rect 390468 385018 390520 385024
rect 390480 383316 390508 385018
rect 392872 383316 392900 385562
rect 399668 385484 399720 385490
rect 399668 385426 399720 385432
rect 397460 385280 397512 385286
rect 397460 385222 397512 385228
rect 395068 385212 395120 385218
rect 395068 385154 395120 385160
rect 395080 383316 395108 385154
rect 397472 383316 397500 385222
rect 399680 383316 399708 385426
rect 402060 385416 402112 385422
rect 402060 385358 402112 385364
rect 402072 383316 402100 385358
rect 403912 383330 403940 393246
rect 408868 385756 408920 385762
rect 408868 385698 408920 385704
rect 406660 385348 406712 385354
rect 406660 385290 406712 385296
rect 403912 383302 404294 383330
rect 406672 383316 406700 385290
rect 408880 383316 408908 385698
rect 411272 383316 411300 407118
rect 416688 389360 416740 389366
rect 416688 389302 416740 389308
rect 416596 389224 416648 389230
rect 416596 389166 416648 389172
rect 413468 385144 413520 385150
rect 413468 385086 413520 385092
rect 413480 383316 413508 385086
rect 380900 381540 380952 381546
rect 380900 381482 380952 381488
rect 380912 381449 380940 381482
rect 380898 381440 380954 381449
rect 380898 381375 380954 381384
rect 380898 377224 380954 377233
rect 380898 377159 380954 377168
rect 380912 376786 380940 377159
rect 380900 376780 380952 376786
rect 380900 376722 380952 376728
rect 380898 374096 380954 374105
rect 380898 374031 380900 374040
rect 380952 374031 380954 374040
rect 414664 374060 414716 374066
rect 380900 374002 380952 374008
rect 414664 374002 414716 374008
rect 380898 370424 380954 370433
rect 380898 370359 380954 370368
rect 380912 369918 380940 370359
rect 380900 369912 380952 369918
rect 380900 369854 380952 369860
rect 381542 367432 381598 367441
rect 381542 367367 381598 367376
rect 380898 363624 380954 363633
rect 380898 363559 380954 363568
rect 380912 362982 380940 363559
rect 380900 362976 380952 362982
rect 380900 362918 380952 362924
rect 380898 353560 380954 353569
rect 380898 353495 380954 353504
rect 380912 353326 380940 353495
rect 380900 353320 380952 353326
rect 380900 353262 380952 353268
rect 381556 340678 381584 367367
rect 381634 360360 381690 360369
rect 381634 360295 381690 360304
rect 381648 340746 381676 360295
rect 381726 356824 381782 356833
rect 381726 356759 381782 356768
rect 381636 340740 381688 340746
rect 381636 340682 381688 340688
rect 381544 340672 381596 340678
rect 381544 340614 381596 340620
rect 381740 340406 381768 356759
rect 383672 350118 384606 350146
rect 383672 340610 383700 350118
rect 386800 347750 386828 350132
rect 386788 347744 386840 347750
rect 386788 347686 386840 347692
rect 389008 347342 389036 350132
rect 391400 347682 391428 350132
rect 391388 347676 391440 347682
rect 391388 347618 391440 347624
rect 393608 347614 393636 350132
rect 393596 347608 393648 347614
rect 393596 347550 393648 347556
rect 396000 347410 396028 350132
rect 398208 347546 398236 350132
rect 398196 347540 398248 347546
rect 398196 347482 398248 347488
rect 395988 347404 396040 347410
rect 395988 347346 396040 347352
rect 388996 347336 389048 347342
rect 388996 347278 389048 347284
rect 400600 347206 400628 350132
rect 402808 347478 402836 350132
rect 404372 350118 405214 350146
rect 402796 347472 402848 347478
rect 402796 347414 402848 347420
rect 400588 347200 400640 347206
rect 400588 347142 400640 347148
rect 404372 340814 404400 350118
rect 407408 347274 407436 350132
rect 408512 350118 409814 350146
rect 407396 347268 407448 347274
rect 407396 347210 407448 347216
rect 408512 340882 408540 350118
rect 412008 347070 412036 350132
rect 414400 347138 414428 350132
rect 414388 347132 414440 347138
rect 414388 347074 414440 347080
rect 411996 347064 412048 347070
rect 411996 347006 412048 347012
rect 408500 340876 408552 340882
rect 408500 340818 408552 340824
rect 404360 340808 404412 340814
rect 404360 340750 404412 340756
rect 383660 340604 383712 340610
rect 383660 340546 383712 340552
rect 381728 340400 381780 340406
rect 381728 340342 381780 340348
rect 401508 337612 401560 337618
rect 401508 337554 401560 337560
rect 380716 203992 380768 203998
rect 380716 203934 380768 203940
rect 380256 203856 380308 203862
rect 380256 203798 380308 203804
rect 401520 202774 401548 337554
rect 411168 337544 411220 337550
rect 411168 337486 411220 337492
rect 408408 337476 408460 337482
rect 408408 337418 408460 337424
rect 400588 202768 400640 202774
rect 400588 202710 400640 202716
rect 401508 202768 401560 202774
rect 401508 202710 401560 202716
rect 401600 202768 401652 202774
rect 401600 202710 401652 202716
rect 379980 201952 380032 201958
rect 379980 201894 380032 201900
rect 400600 200002 400628 202710
rect 401612 202586 401640 202710
rect 401520 202558 401640 202586
rect 401520 201550 401548 202558
rect 400956 201544 401008 201550
rect 400956 201486 401008 201492
rect 401508 201544 401560 201550
rect 401508 201486 401560 201492
rect 400968 200002 400996 201486
rect 408420 200002 408448 337418
rect 411180 202366 411208 337486
rect 413928 337408 413980 337414
rect 413928 337350 413980 337356
rect 413008 202836 413060 202842
rect 413008 202778 413060 202784
rect 413100 202836 413152 202842
rect 413100 202778 413152 202784
rect 413020 202706 413048 202778
rect 412916 202700 412968 202706
rect 412916 202642 412968 202648
rect 413008 202700 413060 202706
rect 413008 202642 413060 202648
rect 412928 202502 412956 202642
rect 412824 202496 412876 202502
rect 412824 202438 412876 202444
rect 412916 202496 412968 202502
rect 412916 202438 412968 202444
rect 410156 202360 410208 202366
rect 410156 202302 410208 202308
rect 411168 202360 411220 202366
rect 411168 202302 411220 202308
rect 409236 202224 409288 202230
rect 409236 202166 409288 202172
rect 409248 200002 409276 202166
rect 410168 200002 410196 202302
rect 411076 202292 411128 202298
rect 411076 202234 411128 202240
rect 355888 199974 355948 200002
rect 356776 199974 357112 200002
rect 357696 199974 357940 200002
rect 358524 199974 358768 200002
rect 359444 199974 359688 200002
rect 360272 199974 360608 200002
rect 361192 199974 361436 200002
rect 362020 199974 362356 200002
rect 362848 199974 362908 200002
rect 363768 199974 364104 200002
rect 364596 199974 364932 200002
rect 365056 199974 365392 200002
rect 365976 199974 366220 200002
rect 366804 199974 366956 200002
rect 374164 199974 374500 200002
rect 375452 199974 375788 200002
rect 376372 199974 376524 200002
rect 400292 199974 400628 200002
rect 400752 199974 400996 200002
rect 408112 199974 408448 200002
rect 408940 199974 409276 200002
rect 409860 199974 410196 200002
rect 411088 200002 411116 202234
rect 412272 201952 412324 201958
rect 412272 201894 412324 201900
rect 412284 200002 412312 201894
rect 412836 201890 412864 202438
rect 412824 201884 412876 201890
rect 412824 201826 412876 201832
rect 413112 200002 413140 202778
rect 413940 200002 413968 337350
rect 414676 202842 414704 374002
rect 414664 202836 414716 202842
rect 414664 202778 414716 202784
rect 415032 202836 415084 202842
rect 415032 202778 415084 202784
rect 415044 202434 415072 202778
rect 415032 202428 415084 202434
rect 415032 202370 415084 202376
rect 415768 202428 415820 202434
rect 415768 202370 415820 202376
rect 414940 202088 414992 202094
rect 414940 202030 414992 202036
rect 414664 202020 414716 202026
rect 414664 201962 414716 201968
rect 414676 201822 414704 201962
rect 414664 201816 414716 201822
rect 414664 201758 414716 201764
rect 414952 200002 414980 202030
rect 415780 200002 415808 202370
rect 416608 200002 416636 389166
rect 416700 202434 416728 389302
rect 416792 374649 416820 407730
rect 416872 407244 416924 407250
rect 416872 407186 416924 407192
rect 416884 380905 416912 407186
rect 418068 389292 418120 389298
rect 418068 389234 418120 389240
rect 416870 380896 416926 380905
rect 416870 380831 416926 380840
rect 417422 376952 417478 376961
rect 417422 376887 417478 376896
rect 416778 374640 416834 374649
rect 416778 374575 416834 374584
rect 416870 370152 416926 370161
rect 416870 370087 416926 370096
rect 416884 202570 416912 370087
rect 416962 367160 417018 367169
rect 416962 367095 417018 367104
rect 416872 202564 416924 202570
rect 416872 202506 416924 202512
rect 416688 202428 416740 202434
rect 416688 202370 416740 202376
rect 416976 202026 417004 367095
rect 417054 363352 417110 363361
rect 417054 363287 417110 363296
rect 416964 202020 417016 202026
rect 416964 201962 417016 201968
rect 417068 201890 417096 363287
rect 417146 360224 417202 360233
rect 417146 360159 417202 360168
rect 417160 202638 417188 360159
rect 417238 356552 417294 356561
rect 417238 356487 417294 356496
rect 417148 202632 417200 202638
rect 417148 202574 417200 202580
rect 417252 202502 417280 356487
rect 417330 353424 417386 353433
rect 417330 353359 417386 353368
rect 417344 202706 417372 353359
rect 417436 202842 417464 376887
rect 418080 202842 418108 389234
rect 417424 202836 417476 202842
rect 417424 202778 417476 202784
rect 417516 202836 417568 202842
rect 417516 202778 417568 202784
rect 418068 202836 418120 202842
rect 418068 202778 418120 202784
rect 417332 202700 417384 202706
rect 417332 202642 417384 202648
rect 417240 202496 417292 202502
rect 417240 202438 417292 202444
rect 417148 202360 417200 202366
rect 417148 202302 417200 202308
rect 417160 202094 417188 202302
rect 417148 202088 417200 202094
rect 417148 202030 417200 202036
rect 417056 201884 417108 201890
rect 417056 201826 417108 201832
rect 417528 200002 417556 202778
rect 418816 201822 418844 556242
rect 418804 201816 418856 201822
rect 418804 201758 418856 201764
rect 411088 199974 411148 200002
rect 411976 199974 412312 200002
rect 412896 199974 413140 200002
rect 413724 199974 413968 200002
rect 414644 199974 414980 200002
rect 415472 199974 415808 200002
rect 416392 199974 416636 200002
rect 417220 199974 417556 200002
rect 238760 199912 238812 199918
rect 238760 199854 238812 199860
rect 239496 199912 239548 199918
rect 239548 199860 239844 199866
rect 239496 199854 239844 199860
rect 239508 199838 239844 199854
rect 433904 157321 433932 699654
rect 433996 159361 434024 700878
rect 434088 163577 434116 700946
rect 434168 700800 434220 700806
rect 434168 700742 434220 700748
rect 434180 165617 434208 700742
rect 434352 700664 434404 700670
rect 434352 700606 434404 700612
rect 438124 700664 438176 700670
rect 438124 700606 438176 700612
rect 434260 623824 434312 623830
rect 434260 623766 434312 623772
rect 434272 173913 434300 623766
rect 434258 173904 434314 173913
rect 434258 173839 434314 173848
rect 434364 167793 434392 700606
rect 434444 700460 434496 700466
rect 434444 700402 434496 700408
rect 434456 169697 434484 700402
rect 436100 700188 436152 700194
rect 436100 700130 436152 700136
rect 434536 681760 434588 681766
rect 434536 681702 434588 681708
rect 434548 172009 434576 681702
rect 434720 336796 434772 336802
rect 434720 336738 434772 336744
rect 434732 184657 434760 336738
rect 434812 294024 434864 294030
rect 434812 293966 434864 293972
rect 434824 186289 434852 293966
rect 434904 251252 434956 251258
rect 434904 251194 434956 251200
rect 434916 188873 434944 251194
rect 434996 207052 435048 207058
rect 434996 206994 435048 207000
rect 435008 190233 435036 206994
rect 434994 190224 435050 190233
rect 434994 190159 435050 190168
rect 434902 188864 434958 188873
rect 434902 188799 434958 188808
rect 434810 186280 434866 186289
rect 434810 186215 434866 186224
rect 434718 184648 434774 184657
rect 434718 184583 434774 184592
rect 434534 172000 434590 172009
rect 434534 171935 434590 171944
rect 434442 169688 434498 169697
rect 434442 169623 434498 169632
rect 434350 167784 434406 167793
rect 434350 167719 434406 167728
rect 434166 165608 434222 165617
rect 434166 165543 434222 165552
rect 434074 163568 434130 163577
rect 434074 163503 434130 163512
rect 436112 161265 436140 700130
rect 436192 392624 436244 392630
rect 436192 392566 436244 392572
rect 436204 180305 436232 392566
rect 436652 201204 436704 201210
rect 436652 201146 436704 201152
rect 436560 201136 436612 201142
rect 436560 201078 436612 201084
rect 436284 199844 436336 199850
rect 436284 199786 436336 199792
rect 436296 193089 436324 199786
rect 436374 196208 436430 196217
rect 436374 196143 436430 196152
rect 436282 193080 436338 193089
rect 436282 193015 436338 193024
rect 436284 192976 436336 192982
rect 436284 192918 436336 192924
rect 436190 180296 436246 180305
rect 436190 180231 436246 180240
rect 436098 161256 436154 161265
rect 436098 161191 436154 161200
rect 433982 159352 434038 159361
rect 433982 159287 434038 159296
rect 433890 157312 433946 157321
rect 433890 157247 433946 157256
rect 436100 155644 436152 155650
rect 436100 155586 436152 155592
rect 436112 155145 436140 155586
rect 436098 155136 436154 155145
rect 436098 155071 436154 155080
rect 436192 148912 436244 148918
rect 436190 148880 436192 148889
rect 436244 148880 436246 148889
rect 436190 148815 436246 148824
rect 436098 146296 436154 146305
rect 436098 146231 436100 146240
rect 436152 146231 436154 146240
rect 436100 146202 436152 146208
rect 436100 142112 436152 142118
rect 436098 142080 436100 142089
rect 436152 142080 436154 142089
rect 436098 142015 436154 142024
rect 134062 130384 134118 130393
rect 134062 130319 134118 130328
rect 436100 128308 436152 128314
rect 436100 128250 436152 128256
rect 436112 127809 436140 128250
rect 436098 127800 436154 127809
rect 436098 127735 436154 127744
rect 133970 123040 134026 123049
rect 133970 122975 134026 122984
rect 133984 120766 134012 122975
rect 134062 121952 134118 121961
rect 134062 121887 134118 121896
rect 134076 120834 134104 121887
rect 134064 120828 134116 120834
rect 134064 120770 134116 120776
rect 133972 120760 134024 120766
rect 133972 120702 134024 120708
rect 151096 120278 151432 120306
rect 156616 120278 156952 120306
rect 133984 120006 134320 120034
rect 134536 120006 134872 120034
rect 135364 120006 135516 120034
rect 135732 120006 136068 120034
rect 136712 120006 136864 120034
rect 133788 117292 133840 117298
rect 133788 117234 133840 117240
rect 133880 117224 133932 117230
rect 133880 117166 133932 117172
rect 133892 117094 133920 117166
rect 133880 117088 133932 117094
rect 133880 117030 133932 117036
rect 133880 113892 133932 113898
rect 133880 113834 133932 113840
rect 133512 88324 133564 88330
rect 133512 88266 133564 88272
rect 133144 67652 133196 67658
rect 133144 67594 133196 67600
rect 133236 67652 133288 67658
rect 133236 67594 133288 67600
rect 133156 60738 133184 67594
rect 133156 60710 133276 60738
rect 133248 57934 133276 60710
rect 132960 57928 133012 57934
rect 132960 57870 133012 57876
rect 133236 57928 133288 57934
rect 133236 57870 133288 57876
rect 132972 50946 133000 57870
rect 132972 50918 133184 50946
rect 133156 41426 133184 50918
rect 133156 41398 133276 41426
rect 133248 38622 133276 41398
rect 132960 38616 133012 38622
rect 132960 38558 133012 38564
rect 133236 38616 133288 38622
rect 133236 38558 133288 38564
rect 132972 31634 133000 38558
rect 132972 31606 133184 31634
rect 132132 30320 132184 30326
rect 132132 30262 132184 30268
rect 133156 22114 133184 31606
rect 133156 22086 133276 22114
rect 133248 12458 133276 22086
rect 133064 12430 133276 12458
rect 133064 9110 133092 12430
rect 133052 9104 133104 9110
rect 133052 9046 133104 9052
rect 131396 8764 131448 8770
rect 131396 8706 131448 8712
rect 130476 4548 130528 4554
rect 130476 4490 130528 4496
rect 131408 480 131436 8706
rect 132592 8696 132644 8702
rect 132592 8638 132644 8644
rect 132604 480 132632 8638
rect 133892 7750 133920 113834
rect 133880 7744 133932 7750
rect 133880 7686 133932 7692
rect 133984 7614 134012 120006
rect 134536 113898 134564 120006
rect 134524 113892 134576 113898
rect 134524 113834 134576 113840
rect 135260 113892 135312 113898
rect 135260 113834 135312 113840
rect 134892 9104 134944 9110
rect 134892 9046 134944 9052
rect 133972 7608 134024 7614
rect 133972 7550 134024 7556
rect 133788 7268 133840 7274
rect 133788 7210 133840 7216
rect 133800 480 133828 7210
rect 134904 480 134932 9046
rect 135272 6186 135300 113834
rect 135364 7682 135392 120006
rect 135444 118312 135496 118318
rect 135444 118254 135496 118260
rect 135352 7676 135404 7682
rect 135352 7618 135404 7624
rect 135456 6322 135484 118254
rect 135732 113898 135760 120006
rect 135720 113892 135772 113898
rect 135720 113834 135772 113840
rect 136732 113892 136784 113898
rect 136732 113834 136784 113840
rect 136640 113824 136692 113830
rect 136640 113766 136692 113772
rect 136088 8628 136140 8634
rect 136088 8570 136140 8576
rect 135444 6316 135496 6322
rect 135444 6258 135496 6264
rect 135260 6180 135312 6186
rect 135260 6122 135312 6128
rect 135352 6180 135404 6186
rect 135352 6122 135404 6128
rect 135364 5574 135392 6122
rect 135352 5568 135404 5574
rect 135352 5510 135404 5516
rect 136100 480 136128 8570
rect 136652 7818 136680 113766
rect 136744 9042 136772 113834
rect 136732 9036 136784 9042
rect 136732 8978 136784 8984
rect 136836 8974 136864 120006
rect 137020 120006 137356 120034
rect 137572 120006 137908 120034
rect 138216 120006 138552 120034
rect 138676 120006 139196 120034
rect 139596 120006 139748 120034
rect 140056 120006 140392 120034
rect 140792 120006 141036 120034
rect 141252 120006 141588 120034
rect 142232 120006 142384 120034
rect 137020 113898 137048 120006
rect 137192 118992 137244 118998
rect 137192 118934 137244 118940
rect 137204 118318 137232 118934
rect 137192 118312 137244 118318
rect 137192 118254 137244 118260
rect 137284 118312 137336 118318
rect 137284 118254 137336 118260
rect 137296 117706 137324 118254
rect 137284 117700 137336 117706
rect 137284 117642 137336 117648
rect 137008 113892 137060 113898
rect 137008 113834 137060 113840
rect 137572 113830 137600 120006
rect 138216 118658 138244 120006
rect 138296 118992 138348 118998
rect 138296 118934 138348 118940
rect 138308 118658 138336 118934
rect 138204 118652 138256 118658
rect 138204 118594 138256 118600
rect 138296 118652 138348 118658
rect 138296 118594 138348 118600
rect 137652 117700 137704 117706
rect 138676 117688 138704 120006
rect 139400 119400 139452 119406
rect 139400 119342 139452 119348
rect 137652 117642 137704 117648
rect 138124 117660 138704 117688
rect 137664 117570 137692 117642
rect 137652 117564 137704 117570
rect 137652 117506 137704 117512
rect 137560 113824 137612 113830
rect 137560 113766 137612 113772
rect 138124 99482 138152 117660
rect 139412 117570 139440 119342
rect 138664 117564 138716 117570
rect 138664 117506 138716 117512
rect 139400 117564 139452 117570
rect 139400 117506 139452 117512
rect 138112 99476 138164 99482
rect 138112 99418 138164 99424
rect 138112 99340 138164 99346
rect 138112 99282 138164 99288
rect 138124 71126 138152 99282
rect 138112 71120 138164 71126
rect 138112 71062 138164 71068
rect 138296 71120 138348 71126
rect 138296 71062 138348 71068
rect 138308 66298 138336 71062
rect 138112 66292 138164 66298
rect 138112 66234 138164 66240
rect 138296 66292 138348 66298
rect 138296 66234 138348 66240
rect 138124 31890 138152 66234
rect 138112 31884 138164 31890
rect 138112 31826 138164 31832
rect 138296 31884 138348 31890
rect 138296 31826 138348 31832
rect 138308 26314 138336 31826
rect 138112 26308 138164 26314
rect 138112 26250 138164 26256
rect 138296 26308 138348 26314
rect 138296 26250 138348 26256
rect 138124 14906 138152 26250
rect 138124 14878 138244 14906
rect 136824 8968 136876 8974
rect 136824 8910 136876 8916
rect 136640 7812 136692 7818
rect 136640 7754 136692 7760
rect 137284 7608 137336 7614
rect 137284 7550 137336 7556
rect 137296 480 137324 7550
rect 138216 6934 138244 14878
rect 138676 9586 138704 117506
rect 139492 113892 139544 113898
rect 139492 113834 139544 113840
rect 138664 9580 138716 9586
rect 138664 9522 138716 9528
rect 138480 8968 138532 8974
rect 138480 8910 138532 8916
rect 138020 6928 138072 6934
rect 138020 6870 138072 6876
rect 138204 6928 138256 6934
rect 138204 6870 138256 6876
rect 138032 3534 138060 6870
rect 138020 3528 138072 3534
rect 138020 3470 138072 3476
rect 138492 480 138520 8910
rect 139504 4826 139532 113834
rect 139492 4820 139544 4826
rect 139492 4762 139544 4768
rect 139596 3466 139624 120006
rect 140056 113898 140084 120006
rect 140792 118561 140820 120006
rect 141252 119354 141280 120006
rect 140884 119326 141280 119354
rect 140778 118552 140834 118561
rect 140778 118487 140834 118496
rect 140044 113892 140096 113898
rect 140044 113834 140096 113840
rect 140884 106457 140912 119326
rect 142252 119128 142304 119134
rect 142252 119070 142304 119076
rect 140870 106448 140926 106457
rect 140870 106383 140926 106392
rect 140778 106312 140834 106321
rect 140778 106247 140780 106256
rect 140832 106247 140834 106256
rect 140964 106276 141016 106282
rect 140780 106218 140832 106224
rect 140964 106218 141016 106224
rect 140976 104854 141004 106218
rect 140964 104848 141016 104854
rect 140964 104790 141016 104796
rect 141148 104848 141200 104854
rect 141148 104790 141200 104796
rect 141160 96370 141188 104790
rect 140976 96342 141188 96370
rect 140976 87038 141004 96342
rect 140872 87032 140924 87038
rect 140872 86974 140924 86980
rect 140964 87032 141016 87038
rect 140964 86974 141016 86980
rect 140884 66314 140912 86974
rect 140792 66286 140912 66314
rect 140792 60897 140820 66286
rect 140778 60888 140834 60897
rect 140778 60823 140834 60832
rect 140778 55312 140834 55321
rect 140778 55247 140834 55256
rect 140792 44146 140820 55247
rect 140792 44118 140912 44146
rect 140884 41449 140912 44118
rect 140870 41440 140926 41449
rect 140870 41375 140926 41384
rect 140778 41304 140834 41313
rect 140778 41239 140834 41248
rect 140792 31770 140820 41239
rect 140792 31742 140912 31770
rect 140884 19310 140912 31742
rect 140872 19304 140924 19310
rect 140872 19246 140924 19252
rect 140964 19236 141016 19242
rect 140964 19178 141016 19184
rect 139676 9036 139728 9042
rect 139676 8978 139728 8984
rect 139584 3460 139636 3466
rect 139584 3402 139636 3408
rect 139688 480 139716 8978
rect 140872 7744 140924 7750
rect 140872 7686 140924 7692
rect 140884 480 140912 7686
rect 140976 3670 141004 19178
rect 142264 4894 142292 119070
rect 142252 4888 142304 4894
rect 142252 4830 142304 4836
rect 142068 4820 142120 4826
rect 142068 4762 142120 4768
rect 140964 3664 141016 3670
rect 140964 3606 141016 3612
rect 142080 480 142108 4762
rect 142356 3602 142384 120006
rect 142540 120006 142876 120034
rect 143092 120006 143428 120034
rect 143552 120006 144072 120034
rect 144380 120006 144716 120034
rect 145024 120006 145268 120034
rect 145576 120006 145912 120034
rect 146312 120006 146556 120034
rect 146680 120006 147108 120034
rect 142540 119134 142568 120006
rect 142528 119128 142580 119134
rect 142528 119070 142580 119076
rect 143092 118658 143120 120006
rect 143080 118652 143132 118658
rect 143080 118594 143132 118600
rect 143448 117224 143500 117230
rect 143448 117166 143500 117172
rect 143460 117094 143488 117166
rect 143448 117088 143500 117094
rect 143448 117030 143500 117036
rect 143264 9580 143316 9586
rect 143264 9522 143316 9528
rect 142344 3596 142396 3602
rect 142344 3538 142396 3544
rect 143276 480 143304 9522
rect 143552 3738 143580 120006
rect 144380 119406 144408 120006
rect 143632 119400 143684 119406
rect 143632 119342 143684 119348
rect 144368 119400 144420 119406
rect 144368 119342 144420 119348
rect 143644 115938 143672 119342
rect 145024 118930 145052 120006
rect 145012 118924 145064 118930
rect 145012 118866 145064 118872
rect 145024 115954 145052 118866
rect 145576 118386 145604 120006
rect 145564 118380 145616 118386
rect 145564 118322 145616 118328
rect 144932 115938 145052 115954
rect 143632 115932 143684 115938
rect 143632 115874 143684 115880
rect 143724 115932 143776 115938
rect 143724 115874 143776 115880
rect 144920 115932 145052 115938
rect 144972 115926 145052 115932
rect 145288 115932 145340 115938
rect 144920 115874 144972 115880
rect 145288 115874 145340 115880
rect 143736 106350 143764 115874
rect 144932 115843 144960 115874
rect 143632 106344 143684 106350
rect 143632 106286 143684 106292
rect 143724 106344 143776 106350
rect 145300 106321 145328 115874
rect 143724 106286 143776 106292
rect 145102 106312 145158 106321
rect 143644 104854 143672 106286
rect 145102 106247 145158 106256
rect 145286 106312 145342 106321
rect 145286 106247 145342 106256
rect 143632 104848 143684 104854
rect 143632 104790 143684 104796
rect 143908 104848 143960 104854
rect 143908 104790 143960 104796
rect 143920 87038 143948 104790
rect 143632 87032 143684 87038
rect 143632 86974 143684 86980
rect 143908 87032 143960 87038
rect 143908 86974 143960 86980
rect 143644 85542 143672 86974
rect 145116 85542 145144 106247
rect 143632 85536 143684 85542
rect 143632 85478 143684 85484
rect 143816 85536 143868 85542
rect 143816 85478 143868 85484
rect 144828 85536 144880 85542
rect 144828 85478 144880 85484
rect 145104 85536 145156 85542
rect 145104 85478 145156 85484
rect 143828 75954 143856 85478
rect 144840 75954 144868 85478
rect 143632 75948 143684 75954
rect 143632 75890 143684 75896
rect 143816 75948 143868 75954
rect 143816 75890 143868 75896
rect 144828 75948 144880 75954
rect 144828 75890 144880 75896
rect 145012 75948 145064 75954
rect 145012 75890 145064 75896
rect 143644 66230 143672 75890
rect 145024 75857 145052 75890
rect 144826 75848 144882 75857
rect 144826 75783 144882 75792
rect 145010 75848 145066 75857
rect 145010 75783 145066 75792
rect 144840 66298 144868 75783
rect 144828 66292 144880 66298
rect 144828 66234 144880 66240
rect 145104 66292 145156 66298
rect 145104 66234 145156 66240
rect 143632 66224 143684 66230
rect 143632 66166 143684 66172
rect 143816 66224 143868 66230
rect 145116 66201 145144 66234
rect 143816 66166 143868 66172
rect 145102 66192 145158 66201
rect 143828 56642 143856 66166
rect 145102 66127 145158 66136
rect 145194 66056 145250 66065
rect 145194 65991 145250 66000
rect 145208 56642 145236 65991
rect 143632 56636 143684 56642
rect 143632 56578 143684 56584
rect 143816 56636 143868 56642
rect 143816 56578 143868 56584
rect 145104 56636 145156 56642
rect 145104 56578 145156 56584
rect 145196 56636 145248 56642
rect 145196 56578 145248 56584
rect 143644 56522 143672 56578
rect 143644 56494 143764 56522
rect 143736 44169 143764 56494
rect 145116 53802 145144 56578
rect 145116 53774 145236 53802
rect 145208 51134 145236 53774
rect 145196 51128 145248 51134
rect 145196 51070 145248 51076
rect 145104 51060 145156 51066
rect 145104 51002 145156 51008
rect 143722 44160 143778 44169
rect 143722 44095 143778 44104
rect 143998 44160 144054 44169
rect 143998 44095 144054 44104
rect 144012 34542 144040 44095
rect 145116 41562 145144 51002
rect 144932 41534 145144 41562
rect 144932 35986 144960 41534
rect 144932 35958 145144 35986
rect 145116 35850 145144 35958
rect 144840 35822 145144 35850
rect 143816 34536 143868 34542
rect 143816 34478 143868 34484
rect 144000 34536 144052 34542
rect 144000 34478 144052 34484
rect 143828 19378 143856 34478
rect 144840 31090 144868 35822
rect 144840 31062 144960 31090
rect 144932 19394 144960 31062
rect 143724 19372 143776 19378
rect 143724 19314 143776 19320
rect 143816 19372 143868 19378
rect 144932 19366 145052 19394
rect 143816 19314 143868 19320
rect 143736 3806 143764 19314
rect 145024 19310 145052 19366
rect 145012 19304 145064 19310
rect 145012 19246 145064 19252
rect 145196 19304 145248 19310
rect 145196 19246 145248 19252
rect 145208 12186 145236 19246
rect 145024 12158 145236 12186
rect 144460 7676 144512 7682
rect 144460 7618 144512 7624
rect 143724 3800 143776 3806
rect 143724 3742 143776 3748
rect 143540 3732 143592 3738
rect 143540 3674 143592 3680
rect 144472 480 144500 7618
rect 145024 4962 145052 12158
rect 145012 4956 145064 4962
rect 145012 4898 145064 4904
rect 145656 4888 145708 4894
rect 145656 4830 145708 4836
rect 145668 480 145696 4830
rect 146312 3874 146340 120006
rect 146680 118130 146708 120006
rect 147738 119762 147766 120020
rect 148060 120006 148396 120034
rect 148612 120006 148948 120034
rect 149072 120006 149592 120034
rect 149900 120006 150236 120034
rect 150452 120006 150788 120034
rect 147738 119734 147812 119762
rect 147784 118862 147812 119734
rect 147772 118856 147824 118862
rect 147772 118798 147824 118804
rect 146760 118652 146812 118658
rect 146760 118594 146812 118600
rect 146404 118102 146708 118130
rect 146404 4418 146432 118102
rect 146482 118008 146538 118017
rect 146482 117943 146538 117952
rect 146496 10402 146524 117943
rect 146772 117570 146800 118594
rect 146852 118380 146904 118386
rect 146852 118322 146904 118328
rect 146864 118017 146892 118322
rect 146850 118008 146906 118017
rect 146850 117943 146906 117952
rect 146760 117564 146812 117570
rect 146760 117506 146812 117512
rect 146484 10396 146536 10402
rect 146484 10338 146536 10344
rect 147784 5030 147812 118798
rect 148060 117434 148088 120006
rect 148048 117428 148100 117434
rect 148048 117370 148100 117376
rect 148612 114578 148640 120006
rect 149072 118794 149100 120006
rect 149060 118788 149112 118794
rect 149060 118730 149112 118736
rect 147956 114572 148008 114578
rect 147956 114514 148008 114520
rect 148600 114572 148652 114578
rect 148600 114514 148652 114520
rect 147968 114442 147996 114514
rect 147956 114436 148008 114442
rect 147956 114378 148008 114384
rect 148232 114436 148284 114442
rect 148232 114378 148284 114384
rect 148244 104961 148272 114378
rect 148046 104952 148102 104961
rect 148046 104887 148102 104896
rect 148230 104952 148286 104961
rect 148230 104887 148286 104896
rect 148060 104854 148088 104887
rect 148048 104848 148100 104854
rect 148048 104790 148100 104796
rect 148232 104848 148284 104854
rect 148232 104790 148284 104796
rect 148244 95266 148272 104790
rect 148048 95260 148100 95266
rect 148048 95202 148100 95208
rect 148232 95260 148284 95266
rect 148232 95202 148284 95208
rect 148060 87038 148088 95202
rect 147864 87032 147916 87038
rect 147864 86974 147916 86980
rect 148048 87032 148100 87038
rect 148048 86974 148100 86980
rect 147876 28914 147904 86974
rect 147876 28886 147996 28914
rect 147772 5024 147824 5030
rect 147772 4966 147824 4972
rect 146392 4412 146444 4418
rect 146392 4354 146444 4360
rect 147968 3942 147996 28886
rect 149072 5098 149100 118730
rect 149900 117910 149928 120006
rect 149888 117904 149940 117910
rect 149888 117846 149940 117852
rect 150452 6338 150480 120006
rect 151096 115954 151124 120278
rect 151832 120006 151984 120034
rect 152476 120006 152628 120034
rect 153272 120006 153424 120034
rect 151832 118697 151860 120006
rect 151818 118688 151874 118697
rect 151818 118623 151874 118632
rect 152476 115977 152504 120006
rect 151004 115926 151124 115954
rect 152186 115968 152242 115977
rect 151004 95266 151032 115926
rect 152186 115903 152242 115912
rect 152462 115968 152518 115977
rect 152462 115903 152518 115912
rect 152200 104854 152228 115903
rect 153292 109812 153344 109818
rect 153292 109754 153344 109760
rect 152096 104848 152148 104854
rect 152096 104790 152148 104796
rect 152188 104848 152240 104854
rect 152188 104790 152240 104796
rect 152108 95266 152136 104790
rect 150716 95260 150768 95266
rect 150716 95202 150768 95208
rect 150992 95260 151044 95266
rect 150992 95202 151044 95208
rect 151820 95260 151872 95266
rect 151820 95202 151872 95208
rect 152096 95260 152148 95266
rect 152096 95202 152148 95208
rect 150728 91798 150756 95202
rect 150532 91792 150584 91798
rect 150532 91734 150584 91740
rect 150716 91792 150768 91798
rect 150716 91734 150768 91740
rect 150544 28966 150572 91734
rect 151832 86986 151860 95202
rect 151832 86970 151952 86986
rect 151820 86964 151964 86970
rect 151872 86958 151912 86964
rect 151820 86906 151872 86912
rect 151912 86906 151964 86912
rect 151832 28966 151860 86906
rect 150532 28960 150584 28966
rect 150532 28902 150584 28908
rect 150624 28960 150676 28966
rect 150624 28902 150676 28908
rect 151820 28960 151872 28966
rect 151820 28902 151872 28908
rect 151912 28960 151964 28966
rect 151912 28902 151964 28908
rect 150636 9178 150664 28902
rect 150624 9172 150676 9178
rect 150624 9114 150676 9120
rect 150360 6310 150480 6338
rect 150360 6186 150388 6310
rect 150348 6180 150400 6186
rect 150348 6122 150400 6128
rect 150440 6180 150492 6186
rect 150440 6122 150492 6128
rect 149060 5092 149112 5098
rect 149060 5034 149112 5040
rect 147956 3936 148008 3942
rect 147956 3878 148008 3884
rect 146300 3868 146352 3874
rect 146300 3810 146352 3816
rect 146852 3528 146904 3534
rect 146852 3470 146904 3476
rect 146864 480 146892 3470
rect 149244 3460 149296 3466
rect 149244 3402 149296 3408
rect 148048 3052 148100 3058
rect 148048 2994 148100 3000
rect 148060 480 148088 2994
rect 149256 480 149284 3402
rect 150452 480 150480 6122
rect 151924 4010 151952 28902
rect 153304 6390 153332 109754
rect 153292 6384 153344 6390
rect 153292 6326 153344 6332
rect 153396 5166 153424 120006
rect 153488 120006 153824 120034
rect 154132 120006 154468 120034
rect 154592 120006 155112 120034
rect 155328 120006 155664 120034
rect 155972 120006 156308 120034
rect 153488 118386 153516 120006
rect 153476 118380 153528 118386
rect 153476 118322 153528 118328
rect 154132 109818 154160 120006
rect 154488 117224 154540 117230
rect 154488 117166 154540 117172
rect 154500 116958 154528 117166
rect 154488 116952 154540 116958
rect 154488 116894 154540 116900
rect 154120 109812 154172 109818
rect 154120 109754 154172 109760
rect 154592 9246 154620 120006
rect 155328 118726 155356 120006
rect 154672 118720 154724 118726
rect 154672 118662 154724 118668
rect 155316 118720 155368 118726
rect 155316 118662 155368 118668
rect 154684 10334 154712 118662
rect 154856 17944 154908 17950
rect 154856 17886 154908 17892
rect 154672 10328 154724 10334
rect 154672 10270 154724 10276
rect 154868 9382 154896 17886
rect 154856 9376 154908 9382
rect 154856 9318 154908 9324
rect 154580 9240 154632 9246
rect 154580 9182 154632 9188
rect 153936 6248 153988 6254
rect 153936 6190 153988 6196
rect 153384 5160 153436 5166
rect 153384 5102 153436 5108
rect 151912 4004 151964 4010
rect 151912 3946 151964 3952
rect 152740 3936 152792 3942
rect 152740 3878 152792 3884
rect 151544 3868 151596 3874
rect 151544 3810 151596 3816
rect 151556 480 151584 3810
rect 152752 480 152780 3878
rect 153948 480 153976 6190
rect 155972 4078 156000 120006
rect 156616 117314 156644 120278
rect 159468 120142 159988 120170
rect 161952 120142 162472 120170
rect 163148 120142 163668 120170
rect 164988 120142 165508 120170
rect 181548 120142 182068 120170
rect 218256 120142 218776 120170
rect 275204 120142 275724 120170
rect 316756 120142 317092 120170
rect 157352 120006 157504 120034
rect 157812 120006 158148 120034
rect 157352 118658 157380 120006
rect 157340 118652 157392 118658
rect 157340 118594 157392 118600
rect 156524 117286 156644 117314
rect 156524 106282 156552 117286
rect 157812 114578 157840 120006
rect 158778 119762 158806 120020
rect 159008 120006 159344 120034
rect 158778 119734 158852 119762
rect 157432 114572 157484 114578
rect 157432 114514 157484 114520
rect 157800 114572 157852 114578
rect 157800 114514 157852 114520
rect 156144 106276 156196 106282
rect 156144 106218 156196 106224
rect 156512 106276 156564 106282
rect 156512 106218 156564 106224
rect 156156 80730 156184 106218
rect 156064 80702 156184 80730
rect 156064 28966 156092 80702
rect 157444 53122 157472 114514
rect 157352 53094 157472 53122
rect 157352 38690 157380 53094
rect 157340 38684 157392 38690
rect 157340 38626 157392 38632
rect 157432 38684 157484 38690
rect 157432 38626 157484 38632
rect 157444 28966 157472 38626
rect 158720 37256 158772 37262
rect 158720 37198 158772 37204
rect 156052 28960 156104 28966
rect 156052 28902 156104 28908
rect 156144 28960 156196 28966
rect 156144 28902 156196 28908
rect 157340 28960 157392 28966
rect 157340 28902 157392 28908
rect 157432 28960 157484 28966
rect 157432 28902 157484 28908
rect 156156 6458 156184 28902
rect 157352 19378 157380 28902
rect 158732 27674 158760 37198
rect 158720 27668 158772 27674
rect 158720 27610 158772 27616
rect 157340 19372 157392 19378
rect 157340 19314 157392 19320
rect 157432 19372 157484 19378
rect 157432 19314 157484 19320
rect 157444 12594 157472 19314
rect 158720 17876 158772 17882
rect 158720 17818 158772 17824
rect 157444 12566 157564 12594
rect 157536 12322 157564 12566
rect 157352 12294 157564 12322
rect 157352 6526 157380 12294
rect 158732 6594 158760 17818
rect 158824 7886 158852 119734
rect 159008 117638 159036 120006
rect 159468 119354 159496 120142
rect 159100 119326 159496 119354
rect 160204 120006 160632 120034
rect 160848 120006 161184 120034
rect 161492 120006 161828 120034
rect 158996 117632 159048 117638
rect 158996 117574 159048 117580
rect 159100 109070 159128 119326
rect 159088 109064 159140 109070
rect 159088 109006 159140 109012
rect 158996 108996 159048 109002
rect 158996 108938 159048 108944
rect 159008 86986 159036 108938
rect 159008 86958 159128 86986
rect 159100 80186 159128 86958
rect 159100 80158 159220 80186
rect 159192 80050 159220 80158
rect 159008 80022 159220 80050
rect 159008 72434 159036 80022
rect 159008 72406 159128 72434
rect 159100 56710 159128 72406
rect 159088 56704 159140 56710
rect 159088 56646 159140 56652
rect 159180 56636 159232 56642
rect 159180 56578 159232 56584
rect 159192 56522 159220 56578
rect 159100 56494 159220 56522
rect 159100 48346 159128 56494
rect 159088 48340 159140 48346
rect 159088 48282 159140 48288
rect 159180 48272 159232 48278
rect 159180 48214 159232 48220
rect 159192 46986 159220 48214
rect 158996 46980 159048 46986
rect 158996 46922 159048 46928
rect 159180 46980 159232 46986
rect 159180 46922 159232 46928
rect 159008 37262 159036 46922
rect 158996 37256 159048 37262
rect 158996 37198 159048 37204
rect 158996 27668 159048 27674
rect 158996 27610 159048 27616
rect 159008 17882 159036 27610
rect 158996 17876 159048 17882
rect 158996 17818 159048 17824
rect 160204 9314 160232 120006
rect 160848 117842 160876 120006
rect 160836 117836 160888 117842
rect 160836 117778 160888 117784
rect 161388 117088 161440 117094
rect 161388 117030 161440 117036
rect 161400 116958 161428 117030
rect 161388 116952 161440 116958
rect 161388 116894 161440 116900
rect 160192 9308 160244 9314
rect 160192 9250 160244 9256
rect 158812 7880 158864 7886
rect 158812 7822 158864 7828
rect 161492 6662 161520 120006
rect 161952 119354 161980 120142
rect 161676 119326 161980 119354
rect 162872 120006 163024 120034
rect 161676 114510 161704 119326
rect 162872 117774 162900 120006
rect 163148 119354 163176 120142
rect 164298 119762 164326 120020
rect 164528 120006 164864 120034
rect 164298 119734 164372 119762
rect 162964 119326 163176 119354
rect 162860 117768 162912 117774
rect 162860 117710 162912 117716
rect 161664 114504 161716 114510
rect 161664 114446 161716 114452
rect 161848 114504 161900 114510
rect 161848 114446 161900 114452
rect 161860 104922 161888 114446
rect 161664 104916 161716 104922
rect 161664 104858 161716 104864
rect 161848 104916 161900 104922
rect 161848 104858 161900 104864
rect 161676 80186 161704 104858
rect 162964 99482 162992 119326
rect 162952 99476 163004 99482
rect 162952 99418 163004 99424
rect 162952 99340 163004 99346
rect 162952 99282 163004 99288
rect 161676 80158 161796 80186
rect 161768 79914 161796 80158
rect 161676 79886 161796 79914
rect 161676 67658 161704 79886
rect 162964 71126 162992 99282
rect 162952 71120 163004 71126
rect 162952 71062 163004 71068
rect 163136 71120 163188 71126
rect 163136 71062 163188 71068
rect 161572 67652 161624 67658
rect 161572 67594 161624 67600
rect 161664 67652 161716 67658
rect 161664 67594 161716 67600
rect 161584 61418 161612 67594
rect 163148 66298 163176 71062
rect 162952 66292 163004 66298
rect 162952 66234 163004 66240
rect 163136 66292 163188 66298
rect 163136 66234 163188 66240
rect 161584 61390 161796 61418
rect 161768 60602 161796 61390
rect 161676 60574 161796 60602
rect 161676 53258 161704 60574
rect 162964 56574 162992 66234
rect 162952 56568 163004 56574
rect 162952 56510 163004 56516
rect 163136 56568 163188 56574
rect 163136 56510 163188 56516
rect 161676 53230 161796 53258
rect 161768 48346 161796 53230
rect 161572 48340 161624 48346
rect 161572 48282 161624 48288
rect 161756 48340 161808 48346
rect 161756 48282 161808 48288
rect 161584 38690 161612 48282
rect 163148 46986 163176 56510
rect 162952 46980 163004 46986
rect 162952 46922 163004 46928
rect 163136 46980 163188 46986
rect 163136 46922 163188 46928
rect 161572 38684 161624 38690
rect 161572 38626 161624 38632
rect 161664 38684 161716 38690
rect 161664 38626 161716 38632
rect 161676 29102 161704 38626
rect 161664 29096 161716 29102
rect 161664 29038 161716 29044
rect 161572 29028 161624 29034
rect 161572 28970 161624 28976
rect 161584 19378 161612 28970
rect 162964 19378 162992 46922
rect 161572 19372 161624 19378
rect 161572 19314 161624 19320
rect 161664 19372 161716 19378
rect 161664 19314 161716 19320
rect 162952 19372 163004 19378
rect 162952 19314 163004 19320
rect 161676 17950 161704 19314
rect 163044 19304 163096 19310
rect 163044 19246 163096 19252
rect 163056 18018 163084 19246
rect 163044 18012 163096 18018
rect 163044 17954 163096 17960
rect 163136 18012 163188 18018
rect 163136 17954 163188 17960
rect 161664 17944 161716 17950
rect 161664 17886 161716 17892
rect 163148 9722 163176 17954
rect 162860 9716 162912 9722
rect 162860 9658 162912 9664
rect 163136 9716 163188 9722
rect 163136 9658 163188 9664
rect 162872 6730 162900 9658
rect 164344 9450 164372 119734
rect 164528 118522 164556 120006
rect 164988 119354 165016 120142
rect 164620 119326 165016 119354
rect 165724 120006 166152 120034
rect 166276 120006 166704 120034
rect 167104 120006 167348 120034
rect 167656 120006 167992 120034
rect 168392 120006 168544 120034
rect 168852 120006 169188 120034
rect 169740 120006 169984 120034
rect 164516 118516 164568 118522
rect 164516 118458 164568 118464
rect 164620 113880 164648 119326
rect 164528 113852 164648 113880
rect 164528 82142 164556 113852
rect 164516 82136 164568 82142
rect 164516 82078 164568 82084
rect 164608 82068 164660 82074
rect 164608 82010 164660 82016
rect 164620 77330 164648 82010
rect 164528 77302 164648 77330
rect 164528 77194 164556 77302
rect 164528 77166 164648 77194
rect 164620 66314 164648 77166
rect 164528 66286 164648 66314
rect 164528 64870 164556 66286
rect 164516 64864 164568 64870
rect 164516 64806 164568 64812
rect 164792 64864 164844 64870
rect 164792 64806 164844 64812
rect 164804 46986 164832 64806
rect 164608 46980 164660 46986
rect 164608 46922 164660 46928
rect 164792 46980 164844 46986
rect 164792 46922 164844 46928
rect 164620 29209 164648 46922
rect 164606 29200 164662 29209
rect 164606 29135 164662 29144
rect 164514 29064 164570 29073
rect 164514 28999 164570 29008
rect 164528 28948 164556 28999
rect 164528 28920 164648 28948
rect 164620 24154 164648 28920
rect 164528 24126 164648 24154
rect 164332 9444 164384 9450
rect 164332 9386 164384 9392
rect 164528 6798 164556 24126
rect 165724 9518 165752 120006
rect 166276 117706 166304 120006
rect 166264 117700 166316 117706
rect 166264 117642 166316 117648
rect 167000 113892 167052 113898
rect 167000 113834 167052 113840
rect 165712 9512 165764 9518
rect 165712 9454 165764 9460
rect 164516 6792 164568 6798
rect 164516 6734 164568 6740
rect 162860 6724 162912 6730
rect 162860 6666 162912 6672
rect 161480 6656 161532 6662
rect 161480 6598 161532 6604
rect 158720 6588 158772 6594
rect 158720 6530 158772 6536
rect 157340 6520 157392 6526
rect 157340 6462 157392 6468
rect 156144 6452 156196 6458
rect 156144 6394 156196 6400
rect 157524 6384 157576 6390
rect 157524 6326 157576 6332
rect 155960 4072 156012 4078
rect 155960 4014 156012 4020
rect 156328 4004 156380 4010
rect 156328 3946 156380 3952
rect 155132 3732 155184 3738
rect 155132 3674 155184 3680
rect 155144 480 155172 3674
rect 156340 480 156368 3946
rect 157536 480 157564 6326
rect 161112 6316 161164 6322
rect 161112 6258 161164 6264
rect 160008 5160 160060 5166
rect 160008 5102 160060 5108
rect 158720 4956 158772 4962
rect 158720 4898 158772 4904
rect 158732 480 158760 4898
rect 160020 3466 160048 5102
rect 160008 3460 160060 3466
rect 160008 3402 160060 3408
rect 159916 2984 159968 2990
rect 159916 2926 159968 2932
rect 159928 480 159956 2926
rect 161124 480 161152 6258
rect 167012 5234 167040 113834
rect 167104 10470 167132 120006
rect 167656 113898 167684 120006
rect 167736 117836 167788 117842
rect 167736 117778 167788 117784
rect 167644 113892 167696 113898
rect 167644 113834 167696 113840
rect 167748 113370 167776 117778
rect 168392 117502 168420 120006
rect 168852 119354 168880 120006
rect 168484 119326 168880 119354
rect 168380 117496 168432 117502
rect 168380 117438 168432 117444
rect 168484 115938 168512 119326
rect 169024 117700 169076 117706
rect 169024 117642 169076 117648
rect 168472 115932 168524 115938
rect 168472 115874 168524 115880
rect 168564 115932 168616 115938
rect 168564 115874 168616 115880
rect 167656 113342 167776 113370
rect 167092 10464 167144 10470
rect 167092 10406 167144 10412
rect 167000 5228 167052 5234
rect 167000 5170 167052 5176
rect 167092 5092 167144 5098
rect 167092 5034 167144 5040
rect 163504 5024 163556 5030
rect 163504 4966 163556 4972
rect 162124 4548 162176 4554
rect 162124 4490 162176 4496
rect 162136 3534 162164 4490
rect 162124 3528 162176 3534
rect 162124 3470 162176 3476
rect 162308 3460 162360 3466
rect 162308 3402 162360 3408
rect 162320 480 162348 3402
rect 163516 480 163544 4966
rect 164700 4072 164752 4078
rect 164700 4014 164752 4020
rect 164712 480 164740 4014
rect 165896 3528 165948 3534
rect 165896 3470 165948 3476
rect 165908 480 165936 3470
rect 167104 480 167132 5034
rect 167656 3194 167684 113342
rect 168576 109070 168604 115874
rect 168564 109064 168616 109070
rect 168564 109006 168616 109012
rect 168472 108996 168524 109002
rect 168472 108938 168524 108944
rect 168484 106298 168512 108938
rect 168484 106270 168604 106298
rect 168392 99414 168420 99445
rect 168576 99414 168604 106270
rect 168380 99408 168432 99414
rect 168564 99408 168616 99414
rect 168432 99356 168564 99362
rect 168380 99350 168616 99356
rect 168392 99334 168604 99350
rect 168576 96626 168604 99334
rect 168380 96620 168432 96626
rect 168380 96562 168432 96568
rect 168564 96620 168616 96626
rect 168564 96562 168616 96568
rect 168392 89434 168420 96562
rect 168392 89406 168604 89434
rect 168576 70258 168604 89406
rect 168484 70230 168604 70258
rect 168484 60738 168512 70230
rect 168484 60710 168604 60738
rect 168576 46986 168604 60710
rect 168472 46980 168524 46986
rect 168472 46922 168524 46928
rect 168564 46980 168616 46986
rect 168564 46922 168616 46928
rect 168484 41426 168512 46922
rect 168484 41398 168604 41426
rect 168576 38622 168604 41398
rect 168380 38616 168432 38622
rect 168380 38558 168432 38564
rect 168564 38616 168616 38622
rect 168564 38558 168616 38564
rect 168392 29050 168420 38558
rect 168392 29022 168512 29050
rect 168484 28966 168512 29022
rect 168472 28960 168524 28966
rect 168472 28902 168524 28908
rect 168656 28960 168708 28966
rect 168656 28902 168708 28908
rect 168668 19394 168696 28902
rect 168392 19366 168696 19394
rect 168392 19310 168420 19366
rect 168196 19304 168248 19310
rect 168196 19246 168248 19252
rect 168380 19304 168432 19310
rect 168380 19246 168432 19252
rect 168208 9722 168236 19246
rect 168196 9716 168248 9722
rect 168196 9658 168248 9664
rect 168472 9716 168524 9722
rect 168472 9658 168524 9664
rect 168484 7954 168512 9658
rect 168472 7948 168524 7954
rect 168472 7890 168524 7896
rect 167644 3188 167696 3194
rect 167644 3130 167696 3136
rect 169036 3126 169064 117642
rect 169852 113892 169904 113898
rect 169852 113834 169904 113840
rect 169864 10538 169892 113834
rect 169852 10532 169904 10538
rect 169852 10474 169904 10480
rect 169956 5302 169984 120006
rect 170048 120006 170384 120034
rect 170692 120006 171028 120034
rect 171244 120006 171580 120034
rect 171888 120006 172224 120034
rect 172624 120006 172868 120034
rect 173084 120006 173420 120034
rect 173912 120006 174064 120034
rect 174372 120006 174708 120034
rect 175260 120006 175504 120034
rect 170048 118454 170076 120006
rect 170404 118652 170456 118658
rect 170404 118594 170456 118600
rect 170036 118448 170088 118454
rect 170036 118390 170088 118396
rect 169944 5296 169996 5302
rect 169944 5238 169996 5244
rect 170416 4146 170444 118594
rect 170692 113898 170720 120006
rect 171140 117224 171192 117230
rect 171138 117192 171140 117201
rect 171192 117192 171194 117201
rect 171138 117127 171194 117136
rect 170680 113892 170732 113898
rect 170680 113834 170732 113840
rect 171244 5370 171272 120006
rect 171888 117638 171916 120006
rect 171876 117632 171928 117638
rect 171876 117574 171928 117580
rect 172520 109132 172572 109138
rect 172520 109074 172572 109080
rect 171784 7812 171836 7818
rect 171784 7754 171836 7760
rect 171232 5364 171284 5370
rect 171232 5306 171284 5312
rect 170588 5228 170640 5234
rect 170588 5170 170640 5176
rect 170404 4140 170456 4146
rect 170404 4082 170456 4088
rect 169392 3596 169444 3602
rect 169392 3538 169444 3544
rect 169024 3120 169076 3126
rect 169024 3062 169076 3068
rect 168196 2916 168248 2922
rect 168196 2858 168248 2864
rect 168208 480 168236 2858
rect 169404 480 169432 3538
rect 170600 480 170628 5170
rect 171796 480 171824 7754
rect 172532 5438 172560 109074
rect 172624 8022 172652 120006
rect 173084 109138 173112 120006
rect 173912 118114 173940 120006
rect 174372 119354 174400 120006
rect 174004 119326 174400 119354
rect 173900 118108 173952 118114
rect 173900 118050 173952 118056
rect 173072 109132 173124 109138
rect 173072 109074 173124 109080
rect 174004 98734 174032 119326
rect 175372 111784 175424 111790
rect 175372 111726 175424 111732
rect 173808 98728 173860 98734
rect 173808 98670 173860 98676
rect 173992 98728 174044 98734
rect 173992 98670 174044 98676
rect 173820 93906 173848 98670
rect 173808 93900 173860 93906
rect 173808 93842 173860 93848
rect 173992 93900 174044 93906
rect 173992 93842 174044 93848
rect 174004 84182 174032 93842
rect 173808 84176 173860 84182
rect 173808 84118 173860 84124
rect 173992 84176 174044 84182
rect 173992 84118 174044 84124
rect 173820 74594 173848 84118
rect 173808 74588 173860 74594
rect 173808 74530 173860 74536
rect 173900 74588 173952 74594
rect 173900 74530 173952 74536
rect 173912 66314 173940 74530
rect 173912 66286 174032 66314
rect 174004 64870 174032 66286
rect 173808 64864 173860 64870
rect 173808 64806 173860 64812
rect 173992 64864 174044 64870
rect 173992 64806 174044 64812
rect 173820 55282 173848 64806
rect 173808 55276 173860 55282
rect 173808 55218 173860 55224
rect 174084 55276 174136 55282
rect 174084 55218 174136 55224
rect 174096 46986 174124 55218
rect 173900 46980 173952 46986
rect 173900 46922 173952 46928
rect 174084 46980 174136 46986
rect 174084 46922 174136 46928
rect 173912 45558 173940 46922
rect 173716 45552 173768 45558
rect 173716 45494 173768 45500
rect 173900 45552 173952 45558
rect 173900 45494 173952 45500
rect 173728 35970 173756 45494
rect 173716 35964 173768 35970
rect 173716 35906 173768 35912
rect 173992 35964 174044 35970
rect 173992 35906 174044 35912
rect 174004 28966 174032 35906
rect 173992 28960 174044 28966
rect 173992 28902 174044 28908
rect 173992 28824 174044 28830
rect 173992 28766 174044 28772
rect 174004 19310 174032 28766
rect 173992 19304 174044 19310
rect 173992 19246 174044 19252
rect 174176 19304 174228 19310
rect 174176 19246 174228 19252
rect 174188 10606 174216 19246
rect 174176 10600 174228 10606
rect 174176 10542 174228 10548
rect 174266 9616 174322 9625
rect 174266 9551 174322 9560
rect 172612 8016 172664 8022
rect 172612 7958 172664 7964
rect 172520 5432 172572 5438
rect 172520 5374 172572 5380
rect 173900 5364 173952 5370
rect 173900 5306 173952 5312
rect 172980 3800 173032 3806
rect 172980 3742 173032 3748
rect 172992 480 173020 3742
rect 173912 3738 173940 5306
rect 174176 5296 174228 5302
rect 174176 5238 174228 5244
rect 173900 3732 173952 3738
rect 173900 3674 173952 3680
rect 174188 480 174216 5238
rect 174280 3398 174308 9551
rect 175384 8090 175412 111726
rect 175372 8084 175424 8090
rect 175372 8026 175424 8032
rect 175476 5506 175504 120006
rect 175568 120006 175904 120034
rect 176212 120006 176548 120034
rect 176764 120006 177100 120034
rect 177408 120006 177744 120034
rect 178144 120006 178388 120034
rect 178604 120006 178940 120034
rect 179432 120006 179584 120034
rect 179984 120006 180228 120034
rect 180780 120006 180932 120034
rect 175568 118250 175596 120006
rect 175556 118244 175608 118250
rect 175556 118186 175608 118192
rect 176212 111790 176240 120006
rect 176568 118108 176620 118114
rect 176568 118050 176620 118056
rect 176200 111784 176252 111790
rect 176200 111726 176252 111732
rect 175464 5500 175516 5506
rect 175464 5442 175516 5448
rect 176580 4146 176608 118050
rect 176764 4758 176792 120006
rect 177408 118182 177436 120006
rect 177396 118176 177448 118182
rect 177396 118118 177448 118124
rect 177948 117972 178000 117978
rect 177948 117914 178000 117920
rect 176752 4752 176804 4758
rect 176752 4694 176804 4700
rect 175372 4140 175424 4146
rect 175372 4082 175424 4088
rect 176568 4140 176620 4146
rect 176568 4082 176620 4088
rect 174268 3392 174320 3398
rect 174268 3334 174320 3340
rect 175384 480 175412 4082
rect 176752 3732 176804 3738
rect 176752 3674 176804 3680
rect 176764 3482 176792 3674
rect 176580 3454 176792 3482
rect 176580 480 176608 3454
rect 177960 626 177988 117914
rect 178040 113892 178092 113898
rect 178040 113834 178092 113840
rect 178052 4622 178080 113834
rect 178144 10674 178172 120006
rect 178604 113898 178632 120006
rect 179328 118176 179380 118182
rect 179328 118118 179380 118124
rect 178592 113892 178644 113898
rect 178592 113834 178644 113840
rect 178132 10668 178184 10674
rect 178132 10610 178184 10616
rect 178040 4616 178092 4622
rect 178040 4558 178092 4564
rect 177776 598 177988 626
rect 179340 610 179368 118118
rect 179432 118046 179460 120006
rect 179420 118040 179472 118046
rect 179420 117982 179472 117988
rect 179984 114578 180012 120006
rect 180706 117192 180762 117201
rect 180706 117127 180762 117136
rect 180720 117094 180748 117127
rect 180708 117088 180760 117094
rect 180708 117030 180760 117036
rect 179604 114572 179656 114578
rect 179604 114514 179656 114520
rect 179972 114572 180024 114578
rect 179972 114514 180024 114520
rect 179616 109138 179644 114514
rect 179604 109132 179656 109138
rect 179604 109074 179656 109080
rect 179604 108996 179656 109002
rect 179604 108938 179656 108944
rect 179616 104938 179644 108938
rect 179616 104910 179736 104938
rect 179708 103494 179736 104910
rect 179604 103488 179656 103494
rect 179604 103430 179656 103436
rect 179696 103488 179748 103494
rect 179696 103430 179748 103436
rect 179616 99414 179644 103430
rect 179604 99408 179656 99414
rect 179604 99350 179656 99356
rect 179696 99340 179748 99346
rect 179696 99282 179748 99288
rect 179708 77330 179736 99282
rect 179616 77302 179736 77330
rect 179616 67726 179644 77302
rect 179604 67720 179656 67726
rect 179604 67662 179656 67668
rect 179696 67516 179748 67522
rect 179696 67458 179748 67464
rect 179708 60738 179736 67458
rect 179616 60710 179736 60738
rect 179616 56574 179644 60710
rect 179512 56568 179564 56574
rect 179512 56510 179564 56516
rect 179604 56568 179656 56574
rect 179604 56510 179656 56516
rect 179524 46986 179552 56510
rect 179512 46980 179564 46986
rect 179512 46922 179564 46928
rect 179696 46980 179748 46986
rect 179696 46922 179748 46928
rect 179708 45558 179736 46922
rect 179420 45552 179472 45558
rect 179420 45494 179472 45500
rect 179696 45552 179748 45558
rect 179696 45494 179748 45500
rect 179432 35970 179460 45494
rect 179420 35964 179472 35970
rect 179420 35906 179472 35912
rect 179604 35964 179656 35970
rect 179604 35906 179656 35912
rect 179616 28966 179644 35906
rect 179604 28960 179656 28966
rect 179604 28902 179656 28908
rect 179696 28960 179748 28966
rect 179696 28902 179748 28908
rect 179708 22012 179736 28902
rect 180708 27600 180760 27606
rect 180708 27542 180760 27548
rect 179616 21984 179736 22012
rect 179616 8158 179644 21984
rect 180720 18018 180748 27542
rect 180708 18012 180760 18018
rect 180708 17954 180760 17960
rect 179604 8152 179656 8158
rect 179604 8094 179656 8100
rect 180904 4690 180932 120006
rect 181088 120006 181424 120034
rect 181088 118590 181116 120006
rect 181548 119354 181576 120142
rect 181180 119326 181576 119354
rect 182284 120006 182620 120034
rect 182928 120006 183264 120034
rect 183572 120006 183908 120034
rect 184032 120006 184460 120034
rect 184952 120006 185104 120034
rect 185412 120006 185748 120034
rect 186300 120006 186452 120034
rect 181076 118584 181128 118590
rect 181076 118526 181128 118532
rect 181180 113880 181208 119326
rect 182180 118380 182232 118386
rect 182180 118322 182232 118328
rect 182192 118153 182220 118322
rect 182178 118144 182234 118153
rect 182178 118079 182234 118088
rect 182088 118040 182140 118046
rect 182088 117982 182140 117988
rect 181088 113852 181208 113880
rect 181088 109018 181116 113852
rect 181088 108990 181208 109018
rect 181180 96626 181208 108990
rect 180984 96620 181036 96626
rect 180984 96562 181036 96568
rect 181168 96620 181220 96626
rect 181168 96562 181220 96568
rect 180996 89690 181024 96562
rect 180984 89684 181036 89690
rect 180984 89626 181036 89632
rect 181168 89684 181220 89690
rect 181168 89626 181220 89632
rect 181180 81954 181208 89626
rect 181088 81926 181208 81954
rect 181088 67726 181116 81926
rect 181076 67720 181128 67726
rect 181076 67662 181128 67668
rect 181168 67516 181220 67522
rect 181168 67458 181220 67464
rect 181180 57934 181208 67458
rect 181076 57928 181128 57934
rect 181076 57870 181128 57876
rect 181168 57928 181220 57934
rect 181168 57870 181220 57876
rect 181088 56574 181116 57870
rect 180984 56568 181036 56574
rect 180984 56510 181036 56516
rect 181076 56568 181128 56574
rect 181076 56510 181128 56516
rect 180996 46986 181024 56510
rect 180984 46980 181036 46986
rect 180984 46922 181036 46928
rect 181168 46980 181220 46986
rect 181168 46922 181220 46928
rect 181180 41562 181208 46922
rect 181180 41534 181300 41562
rect 181272 35986 181300 41534
rect 181180 35958 181300 35986
rect 181180 27606 181208 35958
rect 181168 27600 181220 27606
rect 181168 27542 181220 27548
rect 181076 18012 181128 18018
rect 181076 17954 181128 17960
rect 181088 9625 181116 17954
rect 181074 9616 181130 9625
rect 181074 9551 181130 9560
rect 180892 4684 180944 4690
rect 180892 4626 180944 4632
rect 182100 4146 182128 117982
rect 182180 117428 182232 117434
rect 182180 117370 182232 117376
rect 182192 117230 182220 117370
rect 182180 117224 182232 117230
rect 182180 117166 182232 117172
rect 182284 9654 182312 120006
rect 182928 118318 182956 120006
rect 182916 118312 182968 118318
rect 182916 118254 182968 118260
rect 183468 118312 183520 118318
rect 183468 118254 183520 118260
rect 183374 37224 183430 37233
rect 183374 37159 183430 37168
rect 183388 27674 183416 37159
rect 183376 27668 183428 27674
rect 183376 27610 183428 27616
rect 182272 9648 182324 9654
rect 182272 9590 182324 9596
rect 183480 4146 183508 118254
rect 183572 8226 183600 120006
rect 184032 119354 184060 120006
rect 183756 119326 184060 119354
rect 183756 109154 183784 119326
rect 184848 118244 184900 118250
rect 184848 118186 184900 118192
rect 183756 109126 183876 109154
rect 183848 109018 183876 109126
rect 183756 108990 183876 109018
rect 183756 91746 183784 108990
rect 183664 91718 183784 91746
rect 183664 77314 183692 91718
rect 184756 86964 184808 86970
rect 184756 86906 184808 86912
rect 184768 77314 184796 86906
rect 183652 77308 183704 77314
rect 183652 77250 183704 77256
rect 183744 77308 183796 77314
rect 183744 77250 183796 77256
rect 184756 77308 184808 77314
rect 184756 77250 184808 77256
rect 183756 56642 183784 77250
rect 184756 71120 184808 71126
rect 184756 71062 184808 71068
rect 184768 56642 184796 71062
rect 183744 56636 183796 56642
rect 183744 56578 183796 56584
rect 183836 56636 183888 56642
rect 183836 56578 183888 56584
rect 184756 56636 184808 56642
rect 184756 56578 184808 56584
rect 183848 48362 183876 56578
rect 183848 48334 183968 48362
rect 183940 48226 183968 48334
rect 183756 48198 183968 48226
rect 183650 37224 183706 37233
rect 183756 37210 183784 48198
rect 183706 37182 183784 37210
rect 183650 37159 183706 37168
rect 183836 27668 183888 27674
rect 183836 27610 183888 27616
rect 183848 19394 183876 27610
rect 183756 19366 183876 19394
rect 183756 19310 183784 19366
rect 183744 19304 183796 19310
rect 183744 19246 183796 19252
rect 183928 19304 183980 19310
rect 183928 19246 183980 19252
rect 183940 9897 183968 19246
rect 183926 9888 183982 9897
rect 183926 9823 183982 9832
rect 183650 9752 183706 9761
rect 183650 9687 183706 9696
rect 183664 9654 183692 9687
rect 183652 9648 183704 9654
rect 183652 9590 183704 9596
rect 183836 9648 183888 9654
rect 183836 9590 183888 9596
rect 184296 9648 184348 9654
rect 184296 9590 184348 9596
rect 183848 8906 183876 9590
rect 183836 8900 183888 8906
rect 183836 8842 183888 8848
rect 183560 8220 183612 8226
rect 183560 8162 183612 8168
rect 181352 4140 181404 4146
rect 181352 4082 181404 4088
rect 182088 4140 182140 4146
rect 182088 4082 182140 4088
rect 182548 4140 182600 4146
rect 182548 4082 182600 4088
rect 183468 4140 183520 4146
rect 183468 4082 183520 4088
rect 180064 3800 180116 3806
rect 180064 3742 180116 3748
rect 180156 3800 180208 3806
rect 180156 3742 180208 3748
rect 180076 3194 180104 3742
rect 180064 3188 180116 3194
rect 180064 3130 180116 3136
rect 178960 604 179012 610
rect 177776 480 177804 598
rect 178960 546 179012 552
rect 179328 604 179380 610
rect 179328 546 179380 552
rect 178972 480 179000 546
rect 180168 480 180196 3742
rect 181364 480 181392 4082
rect 182560 480 182588 4082
rect 183744 3392 183796 3398
rect 183744 3334 183796 3340
rect 183756 480 183784 3334
rect 184308 3330 184336 9590
rect 184296 3324 184348 3330
rect 184296 3266 184348 3272
rect 184860 480 184888 118186
rect 184952 117881 184980 120006
rect 185412 119354 185440 120006
rect 185044 119326 185440 119354
rect 184938 117872 184994 117881
rect 184938 117807 184994 117816
rect 185044 114510 185072 119326
rect 186228 118448 186280 118454
rect 186228 118390 186280 118396
rect 185032 114504 185084 114510
rect 185032 114446 185084 114452
rect 185124 114504 185176 114510
rect 185124 114446 185176 114452
rect 185136 99090 185164 114446
rect 185044 99062 185164 99090
rect 185044 89826 185072 99062
rect 186240 96626 186268 118390
rect 186320 113892 186372 113898
rect 186320 113834 186372 113840
rect 186044 96620 186096 96626
rect 186044 96562 186096 96568
rect 186228 96620 186280 96626
rect 186228 96562 186280 96568
rect 186056 95198 186084 96562
rect 185952 95192 186004 95198
rect 185952 95134 186004 95140
rect 186044 95192 186096 95198
rect 186044 95134 186096 95140
rect 185032 89820 185084 89826
rect 185032 89762 185084 89768
rect 184940 89684 184992 89690
rect 184940 89626 184992 89632
rect 184952 86970 184980 89626
rect 184940 86964 184992 86970
rect 184940 86906 184992 86912
rect 185964 85610 185992 95134
rect 185952 85604 186004 85610
rect 185952 85546 186004 85552
rect 186228 85604 186280 85610
rect 186228 85546 186280 85552
rect 185032 77308 185084 77314
rect 185032 77250 185084 77256
rect 185044 71126 185072 77250
rect 186240 76022 186268 85546
rect 186332 76022 186360 113834
rect 186424 76022 186452 120006
rect 186516 120006 186944 120034
rect 187160 120006 187496 120034
rect 187712 120006 188140 120034
rect 186516 117434 186544 120006
rect 186504 117428 186556 117434
rect 186504 117370 186556 117376
rect 186516 76022 186544 117370
rect 187160 113898 187188 120006
rect 187148 113892 187200 113898
rect 187148 113834 187200 113840
rect 186228 76016 186280 76022
rect 186228 75958 186280 75964
rect 186320 76016 186372 76022
rect 186320 75958 186372 75964
rect 186412 76016 186464 76022
rect 186412 75958 186464 75964
rect 186504 76016 186556 76022
rect 186504 75958 186556 75964
rect 186228 75880 186280 75886
rect 186228 75822 186280 75828
rect 186320 75880 186372 75886
rect 186320 75822 186372 75828
rect 186412 75880 186464 75886
rect 186412 75822 186464 75828
rect 186504 75880 186556 75886
rect 186504 75822 186556 75828
rect 186240 74594 186268 75822
rect 186228 74588 186280 74594
rect 186228 74530 186280 74536
rect 185032 71120 185084 71126
rect 185032 71062 185084 71068
rect 186228 66360 186280 66366
rect 186228 66302 186280 66308
rect 186240 66230 186268 66302
rect 186136 66224 186188 66230
rect 186136 66166 186188 66172
rect 186228 66224 186280 66230
rect 186228 66166 186280 66172
rect 186148 56642 186176 66166
rect 184940 56636 184992 56642
rect 184940 56578 184992 56584
rect 186136 56636 186188 56642
rect 186136 56578 186188 56584
rect 186228 56636 186280 56642
rect 186228 56578 186280 56584
rect 184952 43466 184980 56578
rect 184952 43438 185072 43466
rect 185044 38622 185072 43438
rect 184940 38616 184992 38622
rect 184940 38558 184992 38564
rect 185032 38616 185084 38622
rect 185032 38558 185084 38564
rect 184952 28914 184980 38558
rect 184952 28886 185072 28914
rect 185044 9654 185072 28886
rect 186240 27554 186268 56578
rect 185872 27526 186268 27554
rect 185872 9722 185900 27526
rect 185860 9716 185912 9722
rect 185860 9658 185912 9664
rect 186044 9716 186096 9722
rect 186044 9658 186096 9664
rect 185032 9648 185084 9654
rect 185032 9590 185084 9596
rect 186056 480 186084 9658
rect 186228 3664 186280 3670
rect 186148 3612 186228 3618
rect 186148 3606 186280 3612
rect 186148 3590 186268 3606
rect 186148 3194 186176 3590
rect 186332 3262 186360 75822
rect 186424 6866 186452 75822
rect 186412 6860 186464 6866
rect 186412 6802 186464 6808
rect 186516 6118 186544 75822
rect 186596 74588 186648 74594
rect 186596 74530 186648 74536
rect 186608 66366 186636 74530
rect 186596 66360 186648 66366
rect 186596 66302 186648 66308
rect 186504 6112 186556 6118
rect 186504 6054 186556 6060
rect 187712 6050 187740 120006
rect 188770 119814 188798 120020
rect 189092 120006 189336 120034
rect 189644 120006 189980 120034
rect 190472 120006 190624 120034
rect 190748 120006 191176 120034
rect 191820 120006 191972 120034
rect 187792 119808 187844 119814
rect 187792 119750 187844 119756
rect 188758 119808 188810 119814
rect 188758 119750 188810 119756
rect 187804 118386 187832 119750
rect 188988 118516 189040 118522
rect 188988 118458 189040 118464
rect 187792 118380 187844 118386
rect 187792 118322 187844 118328
rect 187700 6044 187752 6050
rect 187700 5986 187752 5992
rect 187804 5982 187832 118322
rect 188620 6520 188672 6526
rect 188620 6462 188672 6468
rect 188068 6452 188120 6458
rect 188068 6394 188120 6400
rect 187792 5976 187844 5982
rect 187792 5918 187844 5924
rect 186320 3256 186372 3262
rect 186320 3198 186372 3204
rect 186136 3188 186188 3194
rect 186136 3130 186188 3136
rect 188080 2922 188108 6394
rect 188436 4140 188488 4146
rect 188436 4082 188488 4088
rect 188068 2916 188120 2922
rect 188068 2858 188120 2864
rect 187240 2848 187292 2854
rect 187240 2790 187292 2796
rect 187252 480 187280 2790
rect 188448 480 188476 4082
rect 188632 4078 188660 6462
rect 189000 4146 189028 118458
rect 189092 117842 189120 120006
rect 189644 119354 189672 120006
rect 189276 119326 189672 119354
rect 189080 117836 189132 117842
rect 189080 117778 189132 117784
rect 189276 114510 189304 119326
rect 190472 117366 190500 120006
rect 190460 117360 190512 117366
rect 190460 117302 190512 117308
rect 190552 117360 190604 117366
rect 190552 117302 190604 117308
rect 189080 114504 189132 114510
rect 189080 114446 189132 114452
rect 189264 114504 189316 114510
rect 189264 114446 189316 114452
rect 189092 104990 189120 114446
rect 189080 104984 189132 104990
rect 189080 104926 189132 104932
rect 189172 104984 189224 104990
rect 189172 104926 189224 104932
rect 189184 103494 189212 104926
rect 189172 103488 189224 103494
rect 189172 103430 189224 103436
rect 189540 103488 189592 103494
rect 189540 103430 189592 103436
rect 189552 95130 189580 103430
rect 189356 95124 189408 95130
rect 189356 95066 189408 95072
rect 189540 95124 189592 95130
rect 189540 95066 189592 95072
rect 189368 85610 189396 95066
rect 189264 85604 189316 85610
rect 189264 85546 189316 85552
rect 189356 85604 189408 85610
rect 189356 85546 189408 85552
rect 189276 77314 189304 85546
rect 189080 77308 189132 77314
rect 189080 77250 189132 77256
rect 189264 77308 189316 77314
rect 189264 77250 189316 77256
rect 189092 75886 189120 77250
rect 189080 75880 189132 75886
rect 189080 75822 189132 75828
rect 189172 75880 189224 75886
rect 189172 75822 189224 75828
rect 189184 70446 189212 75822
rect 189172 70440 189224 70446
rect 189172 70382 189224 70388
rect 189172 70304 189224 70310
rect 189172 70246 189224 70252
rect 189184 60722 189212 70246
rect 189172 60716 189224 60722
rect 189172 60658 189224 60664
rect 189356 60716 189408 60722
rect 189356 60658 189408 60664
rect 189368 51134 189396 60658
rect 189356 51128 189408 51134
rect 189356 51070 189408 51076
rect 189356 50992 189408 50998
rect 189356 50934 189408 50940
rect 189368 38690 189396 50934
rect 189080 38684 189132 38690
rect 189080 38626 189132 38632
rect 189356 38684 189408 38690
rect 189356 38626 189408 38632
rect 189092 29073 189120 38626
rect 189078 29064 189134 29073
rect 189078 28999 189134 29008
rect 189354 28928 189410 28937
rect 189354 28863 189410 28872
rect 189368 5914 189396 28863
rect 190564 10742 190592 117302
rect 190748 109138 190776 120006
rect 191104 117768 191156 117774
rect 191104 117710 191156 117716
rect 190736 109132 190788 109138
rect 190736 109074 190788 109080
rect 190644 108996 190696 109002
rect 190644 108938 190696 108944
rect 190656 96558 190684 108938
rect 190644 96552 190696 96558
rect 190644 96494 190696 96500
rect 190736 96552 190788 96558
rect 190736 96494 190788 96500
rect 190748 80186 190776 96494
rect 190656 80158 190776 80186
rect 190656 31754 190684 80158
rect 190644 31748 190696 31754
rect 190644 31690 190696 31696
rect 190828 31748 190880 31754
rect 190828 31690 190880 31696
rect 190840 21978 190868 31690
rect 190748 21950 190868 21978
rect 190748 12458 190776 21950
rect 190656 12430 190776 12458
rect 190552 10736 190604 10742
rect 190552 10678 190604 10684
rect 190656 7546 190684 12430
rect 190644 7540 190696 7546
rect 190644 7482 190696 7488
rect 189356 5908 189408 5914
rect 189356 5850 189408 5856
rect 188988 4140 189040 4146
rect 188988 4082 189040 4088
rect 188620 4072 188672 4078
rect 188620 4014 188672 4020
rect 189632 4072 189684 4078
rect 189632 4014 189684 4020
rect 189644 480 189672 4014
rect 190828 3120 190880 3126
rect 190828 3062 190880 3068
rect 190840 480 190868 3062
rect 191116 3058 191144 117710
rect 191944 5846 191972 120006
rect 192128 120006 192464 120034
rect 192680 120006 193016 120034
rect 193232 120006 193660 120034
rect 193968 120006 194304 120034
rect 194704 120006 194856 120034
rect 195164 120006 195500 120034
rect 195992 120006 196144 120034
rect 196268 120006 196696 120034
rect 197340 120006 197584 120034
rect 192128 117366 192156 120006
rect 192680 117706 192708 120006
rect 192668 117700 192720 117706
rect 192668 117642 192720 117648
rect 192116 117360 192168 117366
rect 192116 117302 192168 117308
rect 191932 5840 191984 5846
rect 191932 5782 191984 5788
rect 193232 5778 193260 120006
rect 193968 117745 193996 120006
rect 194508 118380 194560 118386
rect 194508 118322 194560 118328
rect 193954 117736 194010 117745
rect 193954 117671 194010 117680
rect 193312 6588 193364 6594
rect 193312 6530 193364 6536
rect 193220 5772 193272 5778
rect 193220 5714 193272 5720
rect 193220 3324 193272 3330
rect 193220 3266 193272 3272
rect 192024 3188 192076 3194
rect 192024 3130 192076 3136
rect 191104 3052 191156 3058
rect 191104 2994 191156 3000
rect 192036 480 192064 3130
rect 193232 480 193260 3266
rect 193324 2990 193352 6530
rect 194520 3330 194548 118322
rect 194600 113892 194652 113898
rect 194600 113834 194652 113840
rect 194612 6746 194640 113834
rect 194704 8294 194732 120006
rect 195164 113898 195192 120006
rect 195888 118584 195940 118590
rect 195888 118526 195940 118532
rect 195152 113892 195204 113898
rect 195152 113834 195204 113840
rect 194692 8288 194744 8294
rect 194692 8230 194744 8236
rect 194612 6718 194732 6746
rect 194600 6656 194652 6662
rect 194600 6598 194652 6604
rect 194612 4010 194640 6598
rect 194704 5710 194732 6718
rect 194692 5704 194744 5710
rect 194692 5646 194744 5652
rect 194600 4004 194652 4010
rect 194600 3946 194652 3952
rect 194508 3324 194560 3330
rect 194508 3266 194560 3272
rect 194600 3324 194652 3330
rect 194600 3266 194652 3272
rect 194416 3052 194468 3058
rect 194416 2994 194468 3000
rect 193312 2984 193364 2990
rect 193312 2926 193364 2932
rect 194428 480 194456 2994
rect 194612 2854 194640 3266
rect 194600 2848 194652 2854
rect 194600 2790 194652 2796
rect 195900 626 195928 118526
rect 195992 118289 196020 120006
rect 196268 119354 196296 120006
rect 196084 119326 196296 119354
rect 195978 118280 196034 118289
rect 195978 118215 196034 118224
rect 196084 109138 196112 119326
rect 197268 117904 197320 117910
rect 197268 117846 197320 117852
rect 196624 117632 196676 117638
rect 196624 117574 196676 117580
rect 196072 109132 196124 109138
rect 196072 109074 196124 109080
rect 196072 108996 196124 109002
rect 196072 108938 196124 108944
rect 196084 106298 196112 108938
rect 196084 106270 196204 106298
rect 196176 80238 196204 106270
rect 196164 80232 196216 80238
rect 196164 80174 196216 80180
rect 196164 80096 196216 80102
rect 196164 80038 196216 80044
rect 196176 79914 196204 80038
rect 196084 79886 196204 79914
rect 196084 70394 196112 79886
rect 196084 70366 196204 70394
rect 196176 60874 196204 70366
rect 196084 60846 196204 60874
rect 196084 60738 196112 60846
rect 195992 60710 196112 60738
rect 195992 60602 196020 60710
rect 195992 60574 196112 60602
rect 196084 51066 196112 60574
rect 196072 51060 196124 51066
rect 196072 51002 196124 51008
rect 196164 50992 196216 50998
rect 196164 50934 196216 50940
rect 196176 12594 196204 50934
rect 196084 12566 196204 12594
rect 196084 12458 196112 12566
rect 195992 12430 196112 12458
rect 195992 7478 196020 12430
rect 195980 7472 196032 7478
rect 195980 7414 196032 7420
rect 196636 3874 196664 117574
rect 197176 6724 197228 6730
rect 197176 6666 197228 6672
rect 196808 4140 196860 4146
rect 196808 4082 196860 4088
rect 196624 3868 196676 3874
rect 196624 3810 196676 3816
rect 195624 598 195928 626
rect 195624 480 195652 598
rect 196820 480 196848 4082
rect 197188 3942 197216 6666
rect 197280 4146 197308 117846
rect 197556 5642 197584 120006
rect 197648 120006 197984 120034
rect 198200 120006 198536 120034
rect 198844 120006 199180 120034
rect 199488 120006 199824 120034
rect 200224 120006 200376 120034
rect 200684 120006 201020 120034
rect 197648 118425 197676 120006
rect 198200 118658 198228 120006
rect 198188 118652 198240 118658
rect 198188 118594 198240 118600
rect 197634 118416 197690 118425
rect 197634 118351 197690 118360
rect 198740 110628 198792 110634
rect 198740 110570 198792 110576
rect 198752 7342 198780 110570
rect 198844 7410 198872 120006
rect 199488 110634 199516 120006
rect 200028 118652 200080 118658
rect 200028 118594 200080 118600
rect 199476 110628 199528 110634
rect 199476 110570 199528 110576
rect 198832 7404 198884 7410
rect 198832 7346 198884 7352
rect 198740 7336 198792 7342
rect 198740 7278 198792 7284
rect 197544 5636 197596 5642
rect 197544 5578 197596 5584
rect 200040 4146 200068 118594
rect 200120 111512 200172 111518
rect 200120 111454 200172 111460
rect 200132 7206 200160 111454
rect 200224 8838 200252 120006
rect 200684 111518 200712 120006
rect 201650 119762 201678 120020
rect 201604 119734 201678 119762
rect 201880 120006 202216 120034
rect 201500 113892 201552 113898
rect 201500 113834 201552 113840
rect 200672 111512 200724 111518
rect 200672 111454 200724 111460
rect 200212 8832 200264 8838
rect 200212 8774 200264 8780
rect 201512 8702 201540 113834
rect 201604 8770 201632 119734
rect 201880 113898 201908 120006
rect 202846 119762 202874 120020
rect 202984 120006 203504 120034
rect 203720 120006 204056 120034
rect 204272 120006 204700 120034
rect 204916 120006 205252 120034
rect 205744 120006 205896 120034
rect 206204 120006 206540 120034
rect 202846 119734 202920 119762
rect 201868 113892 201920 113898
rect 201868 113834 201920 113840
rect 201592 8764 201644 8770
rect 201592 8706 201644 8712
rect 201500 8696 201552 8702
rect 201500 8638 201552 8644
rect 202892 7274 202920 119734
rect 202984 9110 203012 120006
rect 203720 115977 203748 120006
rect 203062 115968 203118 115977
rect 203062 115903 203118 115912
rect 203706 115968 203762 115977
rect 203706 115903 203762 115912
rect 203076 96626 203104 115903
rect 203064 96620 203116 96626
rect 203064 96562 203116 96568
rect 203248 96620 203300 96626
rect 203248 96562 203300 96568
rect 203260 86970 203288 96562
rect 203248 86964 203300 86970
rect 203248 86906 203300 86912
rect 203432 86964 203484 86970
rect 203432 86906 203484 86912
rect 203444 77314 203472 86906
rect 203064 77308 203116 77314
rect 203064 77250 203116 77256
rect 203432 77308 203484 77314
rect 203432 77250 203484 77256
rect 203076 70378 203104 77250
rect 203064 70372 203116 70378
rect 203064 70314 203116 70320
rect 203156 70304 203208 70310
rect 203156 70246 203208 70252
rect 203168 67590 203196 70246
rect 203064 67584 203116 67590
rect 203064 67526 203116 67532
rect 203156 67584 203208 67590
rect 203156 67526 203208 67532
rect 203076 58002 203104 67526
rect 203064 57996 203116 58002
rect 203064 57938 203116 57944
rect 203248 57996 203300 58002
rect 203248 57938 203300 57944
rect 203260 41426 203288 57938
rect 203168 41398 203288 41426
rect 203168 41290 203196 41398
rect 203168 41262 203288 41290
rect 203260 22080 203288 41262
rect 203168 22052 203288 22080
rect 202972 9104 203024 9110
rect 202972 9046 203024 9052
rect 203168 8634 203196 22052
rect 203156 8628 203208 8634
rect 203156 8570 203208 8576
rect 204272 7614 204300 120006
rect 204916 115977 204944 120006
rect 205180 119808 205232 119814
rect 205180 119750 205232 119756
rect 205192 117774 205220 119750
rect 205180 117768 205232 117774
rect 205180 117710 205232 117716
rect 205640 116612 205692 116618
rect 205640 116554 205692 116560
rect 204534 115968 204590 115977
rect 204534 115903 204590 115912
rect 204902 115968 204958 115977
rect 204902 115903 204958 115912
rect 204548 99498 204576 115903
rect 204456 99470 204576 99498
rect 204456 99362 204484 99470
rect 204456 99334 204668 99362
rect 204640 96626 204668 99334
rect 204628 96620 204680 96626
rect 204628 96562 204680 96568
rect 204812 96620 204864 96626
rect 204812 96562 204864 96568
rect 204824 87009 204852 96562
rect 204626 87000 204682 87009
rect 204626 86935 204682 86944
rect 204810 87000 204866 87009
rect 204810 86935 204866 86944
rect 204640 77314 204668 86935
rect 204352 77308 204404 77314
rect 204352 77250 204404 77256
rect 204628 77308 204680 77314
rect 204628 77250 204680 77256
rect 204364 70394 204392 77250
rect 204364 70366 204576 70394
rect 204548 63458 204576 70366
rect 204456 63430 204576 63458
rect 204456 60602 204484 63430
rect 204456 60574 204576 60602
rect 204548 41426 204576 60574
rect 204456 41398 204576 41426
rect 204456 41290 204484 41398
rect 204456 41262 204576 41290
rect 204548 28966 204576 41262
rect 204352 28960 204404 28966
rect 204352 28902 204404 28908
rect 204536 28960 204588 28966
rect 204536 28902 204588 28908
rect 204364 19378 204392 28902
rect 204352 19372 204404 19378
rect 204352 19314 204404 19320
rect 204444 19372 204496 19378
rect 204444 19314 204496 19320
rect 204456 12510 204484 19314
rect 204444 12504 204496 12510
rect 204444 12446 204496 12452
rect 204352 12436 204404 12442
rect 204352 12378 204404 12384
rect 204364 8974 204392 12378
rect 204352 8968 204404 8974
rect 204352 8910 204404 8916
rect 205652 7750 205680 116554
rect 205744 9042 205772 120006
rect 206204 116618 206232 120006
rect 207078 119762 207106 120020
rect 207032 119734 207106 119762
rect 207308 120006 207736 120034
rect 208380 120006 208624 120034
rect 206192 116612 206244 116618
rect 206192 116554 206244 116560
rect 205732 9036 205784 9042
rect 205732 8978 205784 8984
rect 205640 7744 205692 7750
rect 205640 7686 205692 7692
rect 204260 7608 204312 7614
rect 204260 7550 204312 7556
rect 202880 7268 202932 7274
rect 202880 7210 202932 7216
rect 200120 7200 200172 7206
rect 200120 7142 200172 7148
rect 207032 4826 207060 119734
rect 207308 116634 207336 120006
rect 207124 116606 207336 116634
rect 208492 116680 208544 116686
rect 208492 116622 208544 116628
rect 208400 116612 208452 116618
rect 207124 9586 207152 116606
rect 208400 116554 208452 116560
rect 207112 9580 207164 9586
rect 207112 9522 207164 9528
rect 208308 5432 208360 5438
rect 208308 5374 208360 5380
rect 207020 4820 207072 4826
rect 207020 4762 207072 4768
rect 206928 4752 206980 4758
rect 206928 4694 206980 4700
rect 204352 4684 204404 4690
rect 204352 4626 204404 4632
rect 204260 4616 204312 4622
rect 204260 4558 204312 4564
rect 202972 4480 203024 4486
rect 202972 4422 203024 4428
rect 202880 4412 202932 4418
rect 202880 4354 202932 4360
rect 197268 4140 197320 4146
rect 197268 4082 197320 4088
rect 199200 4140 199252 4146
rect 199200 4082 199252 4088
rect 200028 4140 200080 4146
rect 200028 4082 200080 4088
rect 197176 3936 197228 3942
rect 197176 3878 197228 3884
rect 198004 3868 198056 3874
rect 198004 3810 198056 3816
rect 198016 480 198044 3810
rect 199212 480 199240 4082
rect 202696 3936 202748 3942
rect 202696 3878 202748 3884
rect 200396 3256 200448 3262
rect 200396 3198 200448 3204
rect 200408 480 200436 3198
rect 201500 2916 201552 2922
rect 201500 2858 201552 2864
rect 201512 480 201540 2858
rect 202708 480 202736 3878
rect 202892 3398 202920 4354
rect 202880 3392 202932 3398
rect 202880 3334 202932 3340
rect 202984 3330 203012 4422
rect 203892 4140 203944 4146
rect 203892 4082 203944 4088
rect 202972 3324 203024 3330
rect 202972 3266 203024 3272
rect 203904 480 203932 4082
rect 204272 3126 204300 4558
rect 204260 3120 204312 3126
rect 204260 3062 204312 3068
rect 204364 3058 204392 4626
rect 206940 3874 206968 4694
rect 206928 3868 206980 3874
rect 206928 3810 206980 3816
rect 206284 3392 206336 3398
rect 206284 3334 206336 3340
rect 204352 3052 204404 3058
rect 204352 2994 204404 3000
rect 205088 2848 205140 2854
rect 205088 2790 205140 2796
rect 205100 480 205128 2790
rect 206296 480 206324 3334
rect 207480 3324 207532 3330
rect 207480 3266 207532 3272
rect 207492 480 207520 3266
rect 208320 2922 208348 5374
rect 208412 4894 208440 116554
rect 208400 4888 208452 4894
rect 208400 4830 208452 4836
rect 208504 4554 208532 116622
rect 208596 7682 208624 120006
rect 208688 120006 208932 120034
rect 209240 120006 209576 120034
rect 208688 116618 208716 120006
rect 209240 116686 209268 120006
rect 210206 119814 210234 120020
rect 210436 120006 210772 120034
rect 211264 120006 211416 120034
rect 211724 120006 212060 120034
rect 210194 119808 210246 119814
rect 210194 119750 210246 119756
rect 209228 116680 209280 116686
rect 210436 116634 210464 120006
rect 209228 116622 209280 116628
rect 208676 116612 208728 116618
rect 208676 116554 208728 116560
rect 209884 116606 210464 116634
rect 209884 99498 209912 116606
rect 209792 99470 209912 99498
rect 209792 99362 209820 99470
rect 209792 99334 210004 99362
rect 209976 96626 210004 99334
rect 209964 96620 210016 96626
rect 209964 96562 210016 96568
rect 210148 96620 210200 96626
rect 210148 96562 210200 96568
rect 210160 87009 210188 96562
rect 209962 87000 210018 87009
rect 209962 86935 210018 86944
rect 210146 87000 210202 87009
rect 210146 86935 210202 86944
rect 209976 67658 210004 86935
rect 209872 67652 209924 67658
rect 209872 67594 209924 67600
rect 209964 67652 210016 67658
rect 209964 67594 210016 67600
rect 209884 60738 209912 67594
rect 209884 60710 210004 60738
rect 209976 57934 210004 60710
rect 209688 57928 209740 57934
rect 209688 57870 209740 57876
rect 209964 57928 210016 57934
rect 209964 57870 210016 57876
rect 209700 50946 209728 57870
rect 209700 50918 209912 50946
rect 209884 41426 209912 50918
rect 209884 41398 210004 41426
rect 209976 29034 210004 41398
rect 209596 29028 209648 29034
rect 209596 28970 209648 28976
rect 209964 29028 210016 29034
rect 209964 28970 210016 28976
rect 209608 19378 209636 28970
rect 209596 19372 209648 19378
rect 209596 19314 209648 19320
rect 209780 19372 209832 19378
rect 209780 19314 209832 19320
rect 209792 19258 209820 19314
rect 209792 19230 209912 19258
rect 208584 7676 208636 7682
rect 208584 7618 208636 7624
rect 209228 5500 209280 5506
rect 209228 5442 209280 5448
rect 208676 4888 208728 4894
rect 208676 4830 208728 4836
rect 208492 4548 208544 4554
rect 208492 4490 208544 4496
rect 208308 2916 208360 2922
rect 208308 2858 208360 2864
rect 208688 480 208716 4830
rect 209240 2854 209268 5442
rect 209884 5166 209912 19230
rect 211264 6186 211292 120006
rect 211724 117638 211752 120006
rect 212598 119762 212626 120020
rect 212920 120006 213256 120034
rect 212598 119734 212672 119762
rect 211712 117632 211764 117638
rect 211712 117574 211764 117580
rect 212540 116612 212592 116618
rect 212540 116554 212592 116560
rect 212552 6254 212580 116554
rect 212644 6730 212672 119734
rect 212920 116618 212948 120006
rect 213886 119762 213914 120020
rect 214116 120006 214452 120034
rect 214760 120006 215096 120034
rect 215312 120006 215740 120034
rect 216140 120006 216292 120034
rect 216784 120006 216936 120034
rect 217428 120006 217580 120034
rect 213886 119734 213960 119762
rect 213828 117836 213880 117842
rect 213828 117778 213880 117784
rect 213184 117700 213236 117706
rect 213184 117642 213236 117648
rect 212908 116612 212960 116618
rect 212908 116554 212960 116560
rect 212632 6724 212684 6730
rect 212632 6666 212684 6672
rect 212540 6248 212592 6254
rect 212540 6190 212592 6196
rect 211252 6180 211304 6186
rect 211252 6122 211304 6128
rect 209872 5160 209924 5166
rect 209872 5102 209924 5108
rect 212264 4820 212316 4826
rect 212264 4762 212316 4768
rect 209872 4004 209924 4010
rect 209872 3946 209924 3952
rect 209228 2848 209280 2854
rect 209228 2790 209280 2796
rect 209884 480 209912 3946
rect 211068 3868 211120 3874
rect 211068 3810 211120 3816
rect 211080 480 211108 3810
rect 212276 480 212304 4762
rect 213196 3194 213224 117642
rect 213184 3188 213236 3194
rect 213184 3130 213236 3136
rect 213840 626 213868 117778
rect 213932 5370 213960 119734
rect 214012 116612 214064 116618
rect 214012 116554 214064 116560
rect 214024 6390 214052 116554
rect 214116 6662 214144 120006
rect 214760 116618 214788 120006
rect 214748 116612 214800 116618
rect 214748 116554 214800 116560
rect 214104 6656 214156 6662
rect 214104 6598 214156 6604
rect 214012 6384 214064 6390
rect 214012 6326 214064 6332
rect 213920 5364 213972 5370
rect 213920 5306 213972 5312
rect 215312 4962 215340 120006
rect 216140 115977 216168 120006
rect 215942 115968 215998 115977
rect 215942 115903 215998 115912
rect 216126 115968 216182 115977
rect 216126 115903 216182 115912
rect 215956 95266 215984 115903
rect 215576 95260 215628 95266
rect 215576 95202 215628 95208
rect 215944 95260 215996 95266
rect 215944 95202 215996 95208
rect 215588 86970 215616 95202
rect 215484 86964 215536 86970
rect 215484 86906 215536 86912
rect 215576 86964 215628 86970
rect 215576 86906 215628 86912
rect 215496 6594 215524 86906
rect 215484 6588 215536 6594
rect 215484 6530 215536 6536
rect 216784 6322 216812 120006
rect 217428 115977 217456 120006
rect 218118 119762 218146 120020
rect 218072 119734 218146 119762
rect 217968 117768 218020 117774
rect 217968 117710 218020 117716
rect 217046 115968 217102 115977
rect 217046 115903 217102 115912
rect 217414 115968 217470 115977
rect 217414 115903 217470 115912
rect 217060 106486 217088 115903
rect 217048 106480 217100 106486
rect 217048 106422 217100 106428
rect 216956 106344 217008 106350
rect 216956 106286 217008 106292
rect 216968 99482 216996 106286
rect 216956 99476 217008 99482
rect 216956 99418 217008 99424
rect 216956 99340 217008 99346
rect 216956 99282 217008 99288
rect 216968 95266 216996 99282
rect 216956 95260 217008 95266
rect 216956 95202 217008 95208
rect 217048 95260 217100 95266
rect 217048 95202 217100 95208
rect 217060 86970 217088 95202
rect 216956 86964 217008 86970
rect 216956 86906 217008 86912
rect 217048 86964 217100 86970
rect 217048 86906 217100 86912
rect 216772 6316 216824 6322
rect 216772 6258 216824 6264
rect 215300 4956 215352 4962
rect 215300 4898 215352 4904
rect 215852 4956 215904 4962
rect 215852 4898 215904 4904
rect 214656 3120 214708 3126
rect 214656 3062 214708 3068
rect 213472 598 213868 626
rect 213472 480 213500 598
rect 214668 480 214696 3062
rect 215864 480 215892 4898
rect 216968 3466 216996 86906
rect 216956 3460 217008 3466
rect 216956 3402 217008 3408
rect 217980 3058 218008 117710
rect 218072 5030 218100 119734
rect 218256 115954 218284 120142
rect 219406 119762 219434 120020
rect 219544 120006 219972 120034
rect 220372 120006 220616 120034
rect 220832 120006 221260 120034
rect 221660 120006 221812 120034
rect 222304 120006 222456 120034
rect 222672 120006 223008 120034
rect 219406 119734 219480 119762
rect 218256 115926 218376 115954
rect 218348 104922 218376 115926
rect 218244 104916 218296 104922
rect 218244 104858 218296 104864
rect 218336 104916 218388 104922
rect 218336 104858 218388 104864
rect 218256 104825 218284 104858
rect 218242 104816 218298 104825
rect 218242 104751 218298 104760
rect 218426 104680 218482 104689
rect 218426 104615 218482 104624
rect 218440 95266 218468 104615
rect 218336 95260 218388 95266
rect 218336 95202 218388 95208
rect 218428 95260 218480 95266
rect 218428 95202 218480 95208
rect 218348 86970 218376 95202
rect 218244 86964 218296 86970
rect 218244 86906 218296 86912
rect 218336 86964 218388 86970
rect 218336 86906 218388 86912
rect 218256 85542 218284 86906
rect 218244 85536 218296 85542
rect 218244 85478 218296 85484
rect 218428 85536 218480 85542
rect 218428 85478 218480 85484
rect 218440 75954 218468 85478
rect 218244 75948 218296 75954
rect 218244 75890 218296 75896
rect 218428 75948 218480 75954
rect 218428 75890 218480 75896
rect 218256 56574 218284 75890
rect 218152 56568 218204 56574
rect 218152 56510 218204 56516
rect 218244 56568 218296 56574
rect 218244 56510 218296 56516
rect 218164 46986 218192 56510
rect 218152 46980 218204 46986
rect 218152 46922 218204 46928
rect 218428 46980 218480 46986
rect 218428 46922 218480 46928
rect 218440 29034 218468 46922
rect 218244 29028 218296 29034
rect 218244 28970 218296 28976
rect 218428 29028 218480 29034
rect 218428 28970 218480 28976
rect 218256 6526 218284 28970
rect 218244 6520 218296 6526
rect 218244 6462 218296 6468
rect 218060 5024 218112 5030
rect 218060 4966 218112 4972
rect 219348 5024 219400 5030
rect 219348 4966 219400 4972
rect 218152 3460 218204 3466
rect 218152 3402 218204 3408
rect 217048 3052 217100 3058
rect 217048 2994 217100 3000
rect 217968 3052 218020 3058
rect 217968 2994 218020 3000
rect 217060 480 217088 2994
rect 218164 480 218192 3402
rect 219360 480 219388 4966
rect 219452 3534 219480 119734
rect 219544 5098 219572 120006
rect 220372 115977 220400 120006
rect 220174 115968 220230 115977
rect 220174 115903 220230 115912
rect 220358 115968 220414 115977
rect 220358 115903 220414 115912
rect 220188 99090 220216 115903
rect 219820 99062 220216 99090
rect 219820 86970 219848 99062
rect 219716 86964 219768 86970
rect 219716 86906 219768 86912
rect 219808 86964 219860 86970
rect 219808 86906 219860 86912
rect 219728 66298 219756 86906
rect 219624 66292 219676 66298
rect 219624 66234 219676 66240
rect 219716 66292 219768 66298
rect 219716 66234 219768 66240
rect 219636 56710 219664 66234
rect 219624 56704 219676 56710
rect 219624 56646 219676 56652
rect 219808 56704 219860 56710
rect 219808 56646 219860 56652
rect 219820 53258 219848 56646
rect 219820 53230 220032 53258
rect 220004 47002 220032 53230
rect 219912 46974 220032 47002
rect 219912 45558 219940 46974
rect 219716 45552 219768 45558
rect 219716 45494 219768 45500
rect 219900 45552 219952 45558
rect 219900 45494 219952 45500
rect 219728 35970 219756 45494
rect 219716 35964 219768 35970
rect 219716 35906 219768 35912
rect 219992 35964 220044 35970
rect 219992 35906 220044 35912
rect 220004 29102 220032 35906
rect 219992 29096 220044 29102
rect 219992 29038 220044 29044
rect 219808 28960 219860 28966
rect 219808 28902 219860 28908
rect 219820 18018 219848 28902
rect 219716 18012 219768 18018
rect 219716 17954 219768 17960
rect 219808 18012 219860 18018
rect 219808 17954 219860 17960
rect 219728 6458 219756 17954
rect 219716 6452 219768 6458
rect 219716 6394 219768 6400
rect 219532 5092 219584 5098
rect 219532 5034 219584 5040
rect 220832 3602 220860 120006
rect 221660 115977 221688 120006
rect 221462 115968 221518 115977
rect 221462 115903 221518 115912
rect 221646 115968 221702 115977
rect 221646 115903 221702 115912
rect 221476 104854 221504 115903
rect 222200 113756 222252 113762
rect 222200 113698 222252 113704
rect 221280 104848 221332 104854
rect 221280 104790 221332 104796
rect 221464 104848 221516 104854
rect 221464 104790 221516 104796
rect 221292 99090 221320 104790
rect 221108 99062 221320 99090
rect 221108 80050 221136 99062
rect 221016 80022 221136 80050
rect 221016 75886 221044 80022
rect 221004 75880 221056 75886
rect 221004 75822 221056 75828
rect 221280 75880 221332 75886
rect 221280 75822 221332 75828
rect 221292 66337 221320 75822
rect 221094 66328 221150 66337
rect 221094 66263 221150 66272
rect 221278 66328 221334 66337
rect 221278 66263 221334 66272
rect 221108 66230 221136 66263
rect 221004 66224 221056 66230
rect 221004 66166 221056 66172
rect 221096 66224 221148 66230
rect 221096 66166 221148 66172
rect 221016 64870 221044 66166
rect 221004 64864 221056 64870
rect 221004 64806 221056 64812
rect 221188 64864 221240 64870
rect 221188 64806 221240 64812
rect 221200 55282 221228 64806
rect 221004 55276 221056 55282
rect 221004 55218 221056 55224
rect 221188 55276 221240 55282
rect 221188 55218 221240 55224
rect 221016 45558 221044 55218
rect 221004 45552 221056 45558
rect 221004 45494 221056 45500
rect 221280 45552 221332 45558
rect 221280 45494 221332 45500
rect 221292 27674 221320 45494
rect 221096 27668 221148 27674
rect 221096 27610 221148 27616
rect 221280 27668 221332 27674
rect 221280 27610 221332 27616
rect 221108 18018 221136 27610
rect 221004 18012 221056 18018
rect 221004 17954 221056 17960
rect 221096 18012 221148 18018
rect 221096 17954 221148 17960
rect 221016 5234 221044 17954
rect 221004 5228 221056 5234
rect 221004 5170 221056 5176
rect 222108 3800 222160 3806
rect 222108 3742 222160 3748
rect 220820 3596 220872 3602
rect 220820 3538 220872 3544
rect 222120 3534 222148 3742
rect 222212 3670 222240 113698
rect 222304 7818 222332 120006
rect 222672 113762 222700 120006
rect 223638 119762 223666 120020
rect 223960 120006 224296 120034
rect 224420 120006 224848 120034
rect 225156 120006 225492 120034
rect 225800 120006 226136 120034
rect 226444 120006 226688 120034
rect 226996 120006 227332 120034
rect 227732 120006 227976 120034
rect 228284 120006 228528 120034
rect 223638 119734 223712 119762
rect 222660 113756 222712 113762
rect 222660 113698 222712 113704
rect 222292 7812 222344 7818
rect 222292 7754 222344 7760
rect 223684 5302 223712 119734
rect 223960 118114 223988 120006
rect 223948 118108 224000 118114
rect 223948 118050 224000 118056
rect 224420 117722 224448 120006
rect 225156 117978 225184 120006
rect 225800 118182 225828 120006
rect 225788 118176 225840 118182
rect 225788 118118 225840 118124
rect 225144 117972 225196 117978
rect 225144 117914 225196 117920
rect 226248 117972 226300 117978
rect 226248 117914 226300 117920
rect 223776 117694 224448 117722
rect 223672 5296 223724 5302
rect 223672 5238 223724 5244
rect 222844 3800 222896 3806
rect 222844 3742 222896 3748
rect 222200 3664 222252 3670
rect 222200 3606 222252 3612
rect 222856 3534 222884 3742
rect 223776 3738 223804 117694
rect 224224 117632 224276 117638
rect 224224 117574 224276 117580
rect 223764 3732 223816 3738
rect 223764 3674 223816 3680
rect 219440 3528 219492 3534
rect 219440 3470 219492 3476
rect 222108 3528 222160 3534
rect 222108 3470 222160 3476
rect 222844 3528 222896 3534
rect 222844 3470 222896 3476
rect 222936 3528 222988 3534
rect 222936 3470 222988 3476
rect 220544 3188 220596 3194
rect 220544 3130 220596 3136
rect 220556 480 220584 3130
rect 221740 2984 221792 2990
rect 221740 2926 221792 2932
rect 221752 480 221780 2926
rect 222948 480 222976 3470
rect 224236 3262 224264 117574
rect 225604 117360 225656 117366
rect 225604 117302 225656 117308
rect 225616 4078 225644 117302
rect 225604 4072 225656 4078
rect 225604 4014 225656 4020
rect 226260 3330 226288 117914
rect 226444 3806 226472 120006
rect 226996 118046 227024 120006
rect 227732 118318 227760 120006
rect 227720 118312 227772 118318
rect 227720 118254 227772 118260
rect 226984 118040 227036 118046
rect 226984 117982 227036 117988
rect 228284 115977 228312 120006
rect 229158 119762 229186 120020
rect 229480 120006 229816 120034
rect 229940 120006 230368 120034
rect 230676 120006 231012 120034
rect 231320 120006 231656 120034
rect 231964 120006 232208 120034
rect 232516 120006 232852 120034
rect 233252 120006 233496 120034
rect 233712 120006 234048 120034
rect 229158 119734 229232 119762
rect 229204 118250 229232 119734
rect 229480 118454 229508 120006
rect 229468 118448 229520 118454
rect 229468 118390 229520 118396
rect 229192 118244 229244 118250
rect 229192 118186 229244 118192
rect 229008 118040 229060 118046
rect 229008 117982 229060 117988
rect 227994 115968 228050 115977
rect 227994 115903 228050 115912
rect 228270 115968 228326 115977
rect 228270 115903 228326 115912
rect 228008 109018 228036 115903
rect 227916 108990 228036 109018
rect 227916 99482 227944 108990
rect 227904 99476 227956 99482
rect 227904 99418 227956 99424
rect 227812 99340 227864 99346
rect 227812 99282 227864 99288
rect 227824 89758 227852 99282
rect 227812 89752 227864 89758
rect 227812 89694 227864 89700
rect 227904 89616 227956 89622
rect 227904 89558 227956 89564
rect 227916 85542 227944 89558
rect 227536 85536 227588 85542
rect 227536 85478 227588 85484
rect 227904 85536 227956 85542
rect 227904 85478 227956 85484
rect 227548 75954 227576 85478
rect 227536 75948 227588 75954
rect 227536 75890 227588 75896
rect 227720 75948 227772 75954
rect 227720 75890 227772 75896
rect 227732 70258 227760 75890
rect 227732 70230 227852 70258
rect 227824 60722 227852 70230
rect 227812 60716 227864 60722
rect 227812 60658 227864 60664
rect 227996 60716 228048 60722
rect 227996 60658 228048 60664
rect 228008 57934 228036 60658
rect 227720 57928 227772 57934
rect 227720 57870 227772 57876
rect 227996 57928 228048 57934
rect 227996 57870 228048 57876
rect 227732 48346 227760 57870
rect 227720 48340 227772 48346
rect 227720 48282 227772 48288
rect 227904 48340 227956 48346
rect 227904 48282 227956 48288
rect 227916 41614 227944 48282
rect 227904 41608 227956 41614
rect 227904 41550 227956 41556
rect 227904 41472 227956 41478
rect 227904 41414 227956 41420
rect 227916 31822 227944 41414
rect 227904 31816 227956 31822
rect 227904 31758 227956 31764
rect 227904 31680 227956 31686
rect 227904 31622 227956 31628
rect 227916 29034 227944 31622
rect 227812 29028 227864 29034
rect 227812 28970 227864 28976
rect 227904 29028 227956 29034
rect 227904 28970 227956 28976
rect 227824 28937 227852 28970
rect 227810 28928 227866 28937
rect 227810 28863 227866 28872
rect 227994 28928 228050 28937
rect 227994 28863 228050 28872
rect 228008 4418 228036 28863
rect 227996 4412 228048 4418
rect 227996 4354 228048 4360
rect 226432 3800 226484 3806
rect 226432 3742 226484 3748
rect 228916 3800 228968 3806
rect 228916 3742 228968 3748
rect 226524 3732 226576 3738
rect 226524 3674 226576 3680
rect 225236 3324 225288 3330
rect 225236 3266 225288 3272
rect 225328 3324 225380 3330
rect 225328 3266 225380 3272
rect 226248 3324 226300 3330
rect 226248 3266 226300 3272
rect 224224 3256 224276 3262
rect 224224 3198 224276 3204
rect 224132 3052 224184 3058
rect 224132 2994 224184 3000
rect 224144 480 224172 2994
rect 225248 2990 225276 3266
rect 225236 2984 225288 2990
rect 225236 2926 225288 2932
rect 225340 480 225368 3266
rect 226536 480 226564 3674
rect 227720 3664 227772 3670
rect 227720 3606 227772 3612
rect 227732 480 227760 3606
rect 228928 480 228956 3742
rect 229020 3670 229048 117982
rect 229940 117586 229968 120006
rect 230676 118522 230704 120006
rect 230664 118516 230716 118522
rect 230664 118458 230716 118464
rect 231124 118312 231176 118318
rect 231124 118254 231176 118260
rect 229204 117558 229968 117586
rect 229204 4486 229232 117558
rect 229744 117496 229796 117502
rect 229744 117438 229796 117444
rect 229192 4480 229244 4486
rect 229192 4422 229244 4428
rect 229756 4146 229784 117438
rect 229744 4140 229796 4146
rect 229744 4082 229796 4088
rect 231136 3942 231164 118254
rect 231320 117366 231348 120006
rect 231768 118108 231820 118114
rect 231768 118050 231820 118056
rect 231308 117360 231360 117366
rect 231308 117302 231360 117308
rect 231780 4146 231808 118050
rect 231964 4622 231992 120006
rect 232516 117706 232544 120006
rect 233252 118386 233280 120006
rect 233240 118380 233292 118386
rect 233240 118322 233292 118328
rect 233148 118244 233200 118250
rect 233148 118186 233200 118192
rect 232504 117700 232556 117706
rect 232504 117642 232556 117648
rect 232504 117428 232556 117434
rect 232504 117370 232556 117376
rect 231952 4616 232004 4622
rect 231952 4558 232004 4564
rect 232516 4298 232544 117370
rect 232596 117360 232648 117366
rect 232596 117302 232648 117308
rect 232332 4270 232544 4298
rect 231308 4140 231360 4146
rect 231308 4082 231360 4088
rect 231768 4140 231820 4146
rect 231768 4082 231820 4088
rect 231124 3936 231176 3942
rect 231124 3878 231176 3884
rect 230112 3732 230164 3738
rect 230112 3674 230164 3680
rect 229008 3664 229060 3670
rect 229008 3606 229060 3612
rect 230124 480 230152 3674
rect 231320 480 231348 4082
rect 232332 3398 232360 4270
rect 232504 4140 232556 4146
rect 232504 4082 232556 4088
rect 232320 3392 232372 3398
rect 232320 3334 232372 3340
rect 232516 480 232544 4082
rect 232608 2990 232636 117302
rect 232872 9648 232924 9654
rect 232872 9590 232924 9596
rect 232884 5506 232912 9590
rect 232872 5500 232924 5506
rect 232872 5442 232924 5448
rect 233160 4146 233188 118186
rect 233712 113218 233740 120006
rect 234678 119762 234706 120020
rect 235000 120006 235336 120034
rect 235460 120006 235888 120034
rect 236196 120006 236532 120034
rect 236840 120006 237176 120034
rect 237484 120006 237728 120034
rect 238128 120006 238372 120034
rect 238864 120006 239016 120034
rect 239324 120006 239568 120034
rect 234678 119734 234752 119762
rect 234724 118590 234752 119734
rect 234712 118584 234764 118590
rect 234712 118526 234764 118532
rect 234528 118176 234580 118182
rect 234528 118118 234580 118124
rect 233884 117700 233936 117706
rect 233884 117642 233936 117648
rect 233424 113212 233476 113218
rect 233424 113154 233476 113160
rect 233700 113212 233752 113218
rect 233700 113154 233752 113160
rect 233436 106434 233464 113154
rect 233436 106406 233556 106434
rect 233528 104922 233556 106406
rect 233332 104916 233384 104922
rect 233332 104858 233384 104864
rect 233516 104916 233568 104922
rect 233516 104858 233568 104864
rect 233344 103494 233372 104858
rect 233332 103488 233384 103494
rect 233332 103430 233384 103436
rect 233516 103488 233568 103494
rect 233516 103430 233568 103436
rect 233528 95266 233556 103430
rect 233516 95260 233568 95266
rect 233516 95202 233568 95208
rect 233516 95124 233568 95130
rect 233516 95066 233568 95072
rect 233528 89570 233556 95066
rect 233436 89542 233556 89570
rect 233436 80209 233464 89542
rect 233422 80200 233478 80209
rect 233422 80135 233478 80144
rect 233238 79928 233294 79937
rect 233238 79863 233294 79872
rect 233252 74662 233280 79863
rect 233240 74656 233292 74662
rect 233240 74598 233292 74604
rect 233700 74656 233752 74662
rect 233700 74598 233752 74604
rect 233712 58018 233740 74598
rect 233528 57990 233740 58018
rect 233528 57934 233556 57990
rect 233332 57928 233384 57934
rect 233332 57870 233384 57876
rect 233516 57928 233568 57934
rect 233516 57870 233568 57876
rect 233344 48346 233372 57870
rect 233332 48340 233384 48346
rect 233332 48282 233384 48288
rect 233608 48340 233660 48346
rect 233608 48282 233660 48288
rect 233620 38690 233648 48282
rect 233240 38684 233292 38690
rect 233240 38626 233292 38632
rect 233608 38684 233660 38690
rect 233608 38626 233660 38632
rect 233252 31634 233280 38626
rect 233252 31606 233372 31634
rect 233344 28898 233372 31606
rect 233332 28892 233384 28898
rect 233332 28834 233384 28840
rect 233516 28892 233568 28898
rect 233516 28834 233568 28840
rect 233528 4690 233556 28834
rect 233516 4684 233568 4690
rect 233516 4626 233568 4632
rect 233148 4140 233200 4146
rect 233148 4082 233200 4088
rect 233700 4140 233752 4146
rect 233700 4082 233752 4088
rect 232596 2984 232648 2990
rect 232596 2926 232648 2932
rect 233712 480 233740 4082
rect 233896 3126 233924 117642
rect 234540 4146 234568 118118
rect 235000 117910 235028 120006
rect 234988 117904 235040 117910
rect 234988 117846 235040 117852
rect 235460 117688 235488 120006
rect 236196 118658 236224 120006
rect 236184 118652 236236 118658
rect 236184 118594 236236 118600
rect 235908 118448 235960 118454
rect 235908 118390 235960 118396
rect 234724 117660 235488 117688
rect 234724 4758 234752 117660
rect 235264 117564 235316 117570
rect 235264 117506 235316 117512
rect 234712 4752 234764 4758
rect 234712 4694 234764 4700
rect 234528 4140 234580 4146
rect 234528 4082 234580 4088
rect 234804 4140 234856 4146
rect 234804 4082 234856 4088
rect 233884 3120 233936 3126
rect 233884 3062 233936 3068
rect 234816 480 234844 4082
rect 235276 2854 235304 117506
rect 235920 4146 235948 118390
rect 236840 117638 236868 120006
rect 237288 118516 237340 118522
rect 237288 118458 237340 118464
rect 237196 118312 237248 118318
rect 237196 118254 237248 118260
rect 236828 117632 236880 117638
rect 236828 117574 236880 117580
rect 235908 4140 235960 4146
rect 235908 4082 235960 4088
rect 236000 4140 236052 4146
rect 236000 4082 236052 4088
rect 235264 2848 235316 2854
rect 235264 2790 235316 2796
rect 236012 480 236040 4082
rect 237208 480 237236 118254
rect 237300 117722 237328 118458
rect 237300 117694 237420 117722
rect 237288 117632 237340 117638
rect 237288 117574 237340 117580
rect 237300 117366 237328 117574
rect 237288 117360 237340 117366
rect 237288 117302 237340 117308
rect 237392 117178 237420 117694
rect 237300 117150 237420 117178
rect 237300 4146 237328 117150
rect 237484 5438 237512 120006
rect 238128 118386 238156 120006
rect 238116 118380 238168 118386
rect 238116 118322 238168 118328
rect 238668 118380 238720 118386
rect 238668 118322 238720 118328
rect 238116 117904 238168 117910
rect 238116 117846 238168 117852
rect 238128 96642 238156 117846
rect 238036 96614 238156 96642
rect 238036 70394 238064 96614
rect 237944 70366 238064 70394
rect 237944 70258 237972 70366
rect 237944 70230 238064 70258
rect 238036 51082 238064 70230
rect 237944 51054 238064 51082
rect 237944 50946 237972 51054
rect 237944 50918 238064 50946
rect 238036 31770 238064 50918
rect 237944 31742 238064 31770
rect 237944 31634 237972 31742
rect 237944 31606 238064 31634
rect 238036 22098 238064 31606
rect 238024 22092 238076 22098
rect 238024 22034 238076 22040
rect 238116 22024 238168 22030
rect 238116 21966 238168 21972
rect 237472 5432 237524 5438
rect 237472 5374 237524 5380
rect 237288 4140 237340 4146
rect 237288 4082 237340 4088
rect 238128 4010 238156 21966
rect 238116 4004 238168 4010
rect 238116 3946 238168 3952
rect 238680 610 238708 118322
rect 238864 117502 238892 120006
rect 239324 119354 239352 120006
rect 240198 119762 240226 120020
rect 240428 120006 240764 120034
rect 240888 120006 241408 120034
rect 241716 120006 242052 120034
rect 242268 120006 242604 120034
rect 243004 120006 243248 120034
rect 243648 120006 243892 120034
rect 244292 120006 244444 120034
rect 244568 120006 245088 120034
rect 240198 119734 240272 119762
rect 238956 119326 239352 119354
rect 238852 117496 238904 117502
rect 238852 117438 238904 117444
rect 238956 115938 238984 119326
rect 239404 118652 239456 118658
rect 239404 118594 239456 118600
rect 239416 117978 239444 118594
rect 240048 118584 240100 118590
rect 240048 118526 240100 118532
rect 239404 117972 239456 117978
rect 239404 117914 239456 117920
rect 239404 117360 239456 117366
rect 239404 117302 239456 117308
rect 238944 115932 238996 115938
rect 238944 115874 238996 115880
rect 239128 115932 239180 115938
rect 239128 115874 239180 115880
rect 239140 106321 239168 115874
rect 238942 106312 238998 106321
rect 238942 106247 238998 106256
rect 239126 106312 239182 106321
rect 239126 106247 239182 106256
rect 238956 80186 238984 106247
rect 238864 80158 238984 80186
rect 238864 80050 238892 80158
rect 238864 80022 238984 80050
rect 238956 67590 238984 80022
rect 238944 67584 238996 67590
rect 238944 67526 238996 67532
rect 239128 67584 239180 67590
rect 239128 67526 239180 67532
rect 239140 58002 239168 67526
rect 238944 57996 238996 58002
rect 238944 57938 238996 57944
rect 239128 57996 239180 58002
rect 239128 57938 239180 57944
rect 238956 48278 238984 57938
rect 238760 48272 238812 48278
rect 238760 48214 238812 48220
rect 238944 48272 238996 48278
rect 238944 48214 238996 48220
rect 238772 43330 238800 48214
rect 238772 43302 238984 43330
rect 238956 24206 238984 43302
rect 238944 24200 238996 24206
rect 238944 24142 238996 24148
rect 239128 24200 239180 24206
rect 239128 24142 239180 24148
rect 239140 19378 239168 24142
rect 238944 19372 238996 19378
rect 238944 19314 238996 19320
rect 239128 19372 239180 19378
rect 239128 19314 239180 19320
rect 238956 9654 238984 19314
rect 238944 9648 238996 9654
rect 238944 9590 238996 9596
rect 239416 3874 239444 117302
rect 240060 4146 240088 118526
rect 240244 117502 240272 119734
rect 240428 117638 240456 120006
rect 240888 119354 240916 120006
rect 240520 119326 240916 119354
rect 240416 117632 240468 117638
rect 240416 117574 240468 117580
rect 240232 117496 240284 117502
rect 240232 117438 240284 117444
rect 240520 113914 240548 119326
rect 241716 117978 241744 120006
rect 241704 117972 241756 117978
rect 241704 117914 241756 117920
rect 241428 117904 241480 117910
rect 241428 117846 241480 117852
rect 240244 113886 240548 113914
rect 240244 101402 240272 113886
rect 240244 101374 240456 101402
rect 240428 99226 240456 101374
rect 240336 99198 240456 99226
rect 240336 80170 240364 99198
rect 240324 80164 240376 80170
rect 240324 80106 240376 80112
rect 240232 80096 240284 80102
rect 240232 80038 240284 80044
rect 240244 70394 240272 80038
rect 240152 70366 240272 70394
rect 240152 70258 240180 70366
rect 240152 70230 240272 70258
rect 240244 51082 240272 70230
rect 240152 51054 240272 51082
rect 240152 50946 240180 51054
rect 240152 50918 240272 50946
rect 240244 31770 240272 50918
rect 240152 31742 240272 31770
rect 240152 31634 240180 31742
rect 240152 31606 240272 31634
rect 240244 12458 240272 31606
rect 240152 12430 240272 12458
rect 240152 4894 240180 12430
rect 240140 4888 240192 4894
rect 240140 4830 240192 4836
rect 241440 4146 241468 117846
rect 242164 117428 242216 117434
rect 242164 117370 242216 117376
rect 239588 4140 239640 4146
rect 239588 4082 239640 4088
rect 240048 4140 240100 4146
rect 240048 4082 240100 4088
rect 240784 4140 240836 4146
rect 240784 4082 240836 4088
rect 241428 4140 241480 4146
rect 241428 4082 241480 4088
rect 239404 3868 239456 3874
rect 239404 3810 239456 3816
rect 238392 604 238444 610
rect 238392 546 238444 552
rect 238668 604 238720 610
rect 238668 546 238720 552
rect 238404 480 238432 546
rect 239600 480 239628 4082
rect 240796 480 240824 4082
rect 241980 3188 242032 3194
rect 241980 3130 242032 3136
rect 241992 480 242020 3130
rect 242176 3126 242204 117370
rect 242268 117366 242296 120006
rect 242256 117360 242308 117366
rect 242256 117302 242308 117308
rect 242808 117360 242860 117366
rect 242808 117302 242860 117308
rect 242820 3194 242848 117302
rect 243004 4826 243032 120006
rect 243648 117842 243676 120006
rect 243636 117836 243688 117842
rect 243636 117778 243688 117784
rect 244292 117706 244320 120006
rect 244568 119354 244596 120006
rect 245718 119762 245746 120020
rect 244476 119326 244596 119354
rect 245672 119734 245746 119762
rect 245856 120006 246284 120034
rect 246592 120006 246928 120034
rect 247236 120006 247572 120034
rect 247788 120006 248124 120034
rect 248524 120006 248768 120034
rect 249076 120006 249412 120034
rect 249812 120006 249964 120034
rect 250364 120006 250608 120034
rect 244280 117700 244332 117706
rect 244280 117642 244332 117648
rect 244188 117632 244240 117638
rect 244188 117574 244240 117580
rect 243544 117496 243596 117502
rect 243544 117438 243596 117444
rect 242992 4820 243044 4826
rect 242992 4762 243044 4768
rect 243176 4140 243228 4146
rect 243176 4082 243228 4088
rect 242808 3188 242860 3194
rect 242808 3130 242860 3136
rect 242164 3120 242216 3126
rect 242164 3062 242216 3068
rect 243188 480 243216 4082
rect 243556 3058 243584 117438
rect 244096 37256 244148 37262
rect 244096 37198 244148 37204
rect 244108 27674 244136 37198
rect 244096 27668 244148 27674
rect 244096 27610 244148 27616
rect 244200 4146 244228 117574
rect 244476 111058 244504 119326
rect 245672 117774 245700 119734
rect 245752 117836 245804 117842
rect 245752 117778 245804 117784
rect 245660 117768 245712 117774
rect 245660 117710 245712 117716
rect 245568 117700 245620 117706
rect 245568 117642 245620 117648
rect 245384 114572 245436 114578
rect 245384 114514 245436 114520
rect 244292 111030 244504 111058
rect 244292 99362 244320 111030
rect 245396 106350 245424 114514
rect 245384 106344 245436 106350
rect 245384 106286 245436 106292
rect 245476 106344 245528 106350
rect 245476 106286 245528 106292
rect 244292 99334 244504 99362
rect 244476 75954 244504 99334
rect 244280 75948 244332 75954
rect 244280 75890 244332 75896
rect 244464 75948 244516 75954
rect 244464 75890 244516 75896
rect 244292 75857 244320 75890
rect 244278 75848 244334 75857
rect 244278 75783 244334 75792
rect 244646 75848 244702 75857
rect 244646 75783 244702 75792
rect 244660 66298 244688 75783
rect 244372 66292 244424 66298
rect 244372 66234 244424 66240
rect 244648 66292 244700 66298
rect 244648 66234 244700 66240
rect 244384 66178 244412 66234
rect 244292 66150 244412 66178
rect 244292 56642 244320 66150
rect 244280 56636 244332 56642
rect 244280 56578 244332 56584
rect 244556 56636 244608 56642
rect 244556 56578 244608 56584
rect 244568 38690 244596 56578
rect 244280 38684 244332 38690
rect 244280 38626 244332 38632
rect 244556 38684 244608 38690
rect 244556 38626 244608 38632
rect 244292 37262 244320 38626
rect 244280 37256 244332 37262
rect 244280 37198 244332 37204
rect 244372 27668 244424 27674
rect 244372 27610 244424 27616
rect 244384 22098 244412 27610
rect 244372 22092 244424 22098
rect 244372 22034 244424 22040
rect 244556 22092 244608 22098
rect 244556 22034 244608 22040
rect 244568 12050 244596 22034
rect 245488 12458 245516 106286
rect 245304 12430 245516 12458
rect 244568 12022 244688 12050
rect 244660 11778 244688 12022
rect 244568 11750 244688 11778
rect 244568 4962 244596 11750
rect 245304 9738 245332 12430
rect 245304 9710 245424 9738
rect 245396 9654 245424 9710
rect 245384 9648 245436 9654
rect 245384 9590 245436 9596
rect 245476 9580 245528 9586
rect 245476 9522 245528 9528
rect 244556 4956 244608 4962
rect 244556 4898 244608 4904
rect 244188 4140 244240 4146
rect 244188 4082 244240 4088
rect 244372 4140 244424 4146
rect 244372 4082 244424 4088
rect 243544 3052 243596 3058
rect 243544 2994 243596 3000
rect 244384 480 244412 4082
rect 245488 4026 245516 9522
rect 245580 4146 245608 117642
rect 245764 114578 245792 117778
rect 245752 114572 245804 114578
rect 245752 114514 245804 114520
rect 245752 110016 245804 110022
rect 245752 109958 245804 109964
rect 245764 5030 245792 109958
rect 245752 5024 245804 5030
rect 245752 4966 245804 4972
rect 245568 4140 245620 4146
rect 245568 4082 245620 4088
rect 245488 3998 245608 4026
rect 245580 480 245608 3998
rect 245856 3466 245884 120006
rect 246592 110022 246620 120006
rect 246948 117768 247000 117774
rect 246948 117710 247000 117716
rect 246580 110016 246632 110022
rect 246580 109958 246632 109964
rect 246960 106457 246988 117710
rect 247236 117434 247264 120006
rect 247788 117570 247816 120006
rect 247776 117564 247828 117570
rect 247776 117506 247828 117512
rect 248328 117564 248380 117570
rect 248328 117506 248380 117512
rect 247224 117428 247276 117434
rect 247224 117370 247276 117376
rect 248340 115938 248368 117506
rect 248236 115932 248288 115938
rect 248236 115874 248288 115880
rect 248328 115932 248380 115938
rect 248328 115874 248380 115880
rect 246946 106448 247002 106457
rect 246946 106383 247002 106392
rect 248248 106350 248276 115874
rect 248236 106344 248288 106350
rect 246946 106312 247002 106321
rect 248236 106286 248288 106292
rect 248328 106344 248380 106350
rect 248328 106286 248380 106292
rect 246946 106247 247002 106256
rect 246960 9897 246988 106247
rect 248340 18018 248368 106286
rect 247960 18012 248012 18018
rect 247960 17954 248012 17960
rect 248328 18012 248380 18018
rect 248328 17954 248380 17960
rect 246946 9888 247002 9897
rect 246946 9823 247002 9832
rect 246762 9752 246818 9761
rect 246762 9687 246818 9696
rect 246776 9654 246804 9687
rect 247972 9654 248000 17954
rect 246764 9648 246816 9654
rect 246764 9590 246816 9596
rect 247960 9648 248012 9654
rect 247960 9590 248012 9596
rect 246764 9512 246816 9518
rect 246764 9454 246816 9460
rect 247960 9512 248012 9518
rect 247960 9454 248012 9460
rect 245844 3460 245896 3466
rect 245844 3402 245896 3408
rect 246776 480 246804 9454
rect 247972 480 248000 9454
rect 248524 3534 248552 120006
rect 249076 117502 249104 120006
rect 249812 118658 249840 120006
rect 249800 118652 249852 118658
rect 249800 118594 249852 118600
rect 249892 118652 249944 118658
rect 249892 118594 249944 118600
rect 249064 117496 249116 117502
rect 249064 117438 249116 117444
rect 249708 117496 249760 117502
rect 249708 117438 249760 117444
rect 249720 4146 249748 117438
rect 249904 117366 249932 118594
rect 249892 117360 249944 117366
rect 249892 117302 249944 117308
rect 250364 114578 250392 120006
rect 251238 119762 251266 120020
rect 251468 120006 251804 120034
rect 251928 120006 252448 120034
rect 252756 120006 253092 120034
rect 253308 120006 253644 120034
rect 253952 120006 254288 120034
rect 254596 120006 254932 120034
rect 255332 120006 255484 120034
rect 255792 120006 256128 120034
rect 251238 119734 251312 119762
rect 251284 118046 251312 119734
rect 251272 118040 251324 118046
rect 251272 117982 251324 117988
rect 251088 117972 251140 117978
rect 251088 117914 251140 117920
rect 250444 117360 250496 117366
rect 250444 117302 250496 117308
rect 250076 114572 250128 114578
rect 250076 114514 250128 114520
rect 250352 114572 250404 114578
rect 250352 114514 250404 114520
rect 250088 109018 250116 114514
rect 249996 108990 250116 109018
rect 249996 106264 250024 108990
rect 249904 106236 250024 106264
rect 249904 99414 249932 106236
rect 249892 99408 249944 99414
rect 249892 99350 249944 99356
rect 249984 99340 250036 99346
rect 249984 99282 250036 99288
rect 249996 96642 250024 99282
rect 249904 96614 250024 96642
rect 249904 80170 249932 96614
rect 249892 80164 249944 80170
rect 249892 80106 249944 80112
rect 249800 80096 249852 80102
rect 249800 80038 249852 80044
rect 249812 75886 249840 80038
rect 249800 75880 249852 75886
rect 249800 75822 249852 75828
rect 249892 75880 249944 75886
rect 249892 75822 249944 75828
rect 249904 70446 249932 75822
rect 249892 70440 249944 70446
rect 249892 70382 249944 70388
rect 249984 70372 250036 70378
rect 249984 70314 250036 70320
rect 249996 66314 250024 70314
rect 249904 66286 250024 66314
rect 249904 66230 249932 66286
rect 249892 66224 249944 66230
rect 249892 66166 249944 66172
rect 250168 66156 250220 66162
rect 250168 66098 250220 66104
rect 250180 56642 250208 66098
rect 250076 56636 250128 56642
rect 250076 56578 250128 56584
rect 250168 56636 250220 56642
rect 250168 56578 250220 56584
rect 250088 38690 250116 56578
rect 249800 38684 249852 38690
rect 249800 38626 249852 38632
rect 250076 38684 250128 38690
rect 250076 38626 250128 38632
rect 249812 37262 249840 38626
rect 249800 37256 249852 37262
rect 249800 37198 249852 37204
rect 250168 37256 250220 37262
rect 250168 37198 250220 37204
rect 250180 27674 250208 37198
rect 249892 27668 249944 27674
rect 249892 27610 249944 27616
rect 250168 27668 250220 27674
rect 250168 27610 250220 27616
rect 249904 22098 249932 27610
rect 249892 22092 249944 22098
rect 249892 22034 249944 22040
rect 250076 22092 250128 22098
rect 250076 22034 250128 22040
rect 249156 4140 249208 4146
rect 249156 4082 249208 4088
rect 249708 4140 249760 4146
rect 249708 4082 249760 4088
rect 248512 3528 248564 3534
rect 248512 3470 248564 3476
rect 249168 480 249196 4082
rect 250088 3602 250116 22034
rect 250456 3670 250484 117302
rect 250444 3664 250496 3670
rect 250444 3606 250496 3612
rect 250076 3596 250128 3602
rect 250076 3538 250128 3544
rect 251100 3398 251128 117914
rect 251468 117366 251496 120006
rect 251928 119354 251956 120006
rect 251560 119326 251956 119354
rect 251456 117360 251508 117366
rect 251456 117302 251508 117308
rect 251560 113914 251588 119326
rect 252756 118114 252784 120006
rect 253308 118250 253336 120006
rect 253296 118244 253348 118250
rect 253296 118186 253348 118192
rect 253848 118244 253900 118250
rect 253848 118186 253900 118192
rect 252744 118108 252796 118114
rect 252744 118050 252796 118056
rect 253756 118040 253808 118046
rect 253756 117982 253808 117988
rect 252468 117360 252520 117366
rect 252468 117302 252520 117308
rect 251376 113886 251588 113914
rect 251376 109018 251404 113886
rect 251284 108990 251404 109018
rect 251284 106282 251312 108990
rect 251272 106276 251324 106282
rect 251272 106218 251324 106224
rect 251456 106276 251508 106282
rect 251456 106218 251508 106224
rect 251468 96694 251496 106218
rect 251272 96688 251324 96694
rect 251272 96630 251324 96636
rect 251456 96688 251508 96694
rect 251456 96630 251508 96636
rect 251284 89690 251312 96630
rect 251272 89684 251324 89690
rect 251272 89626 251324 89632
rect 251364 89616 251416 89622
rect 251364 89558 251416 89564
rect 251376 66298 251404 89558
rect 251272 66292 251324 66298
rect 251272 66234 251324 66240
rect 251364 66292 251416 66298
rect 251364 66234 251416 66240
rect 251284 60738 251312 66234
rect 251284 60710 251404 60738
rect 251376 38622 251404 60710
rect 251180 38616 251232 38622
rect 251180 38558 251232 38564
rect 251364 38616 251416 38622
rect 251364 38558 251416 38564
rect 251192 31822 251220 38558
rect 251180 31816 251232 31822
rect 251180 31758 251232 31764
rect 251272 31748 251324 31754
rect 251272 31690 251324 31696
rect 251284 22114 251312 31690
rect 251284 22086 251404 22114
rect 251376 12458 251404 22086
rect 251192 12430 251404 12458
rect 251192 3738 251220 12430
rect 252480 4146 252508 117302
rect 253768 115938 253796 117982
rect 253756 115932 253808 115938
rect 253756 115874 253808 115880
rect 253756 106344 253808 106350
rect 253756 106286 253808 106292
rect 253768 104854 253796 106286
rect 253572 104848 253624 104854
rect 253572 104790 253624 104796
rect 253756 104848 253808 104854
rect 253756 104790 253808 104796
rect 253584 95266 253612 104790
rect 253572 95260 253624 95266
rect 253572 95202 253624 95208
rect 253756 95260 253808 95266
rect 253756 95202 253808 95208
rect 253768 85542 253796 95202
rect 253572 85536 253624 85542
rect 253572 85478 253624 85484
rect 253756 85536 253808 85542
rect 253756 85478 253808 85484
rect 253584 75954 253612 85478
rect 253572 75948 253624 75954
rect 253572 75890 253624 75896
rect 253756 75948 253808 75954
rect 253756 75890 253808 75896
rect 253768 56642 253796 75890
rect 253664 56636 253716 56642
rect 253664 56578 253716 56584
rect 253756 56636 253808 56642
rect 253756 56578 253808 56584
rect 253676 48414 253704 56578
rect 253664 48408 253716 48414
rect 253664 48350 253716 48356
rect 253756 48408 253808 48414
rect 253756 48350 253808 48356
rect 253768 46918 253796 48350
rect 253480 46912 253532 46918
rect 253480 46854 253532 46860
rect 253756 46912 253808 46918
rect 253756 46854 253808 46860
rect 253492 37330 253520 46854
rect 253480 37324 253532 37330
rect 253480 37266 253532 37272
rect 253572 37324 253624 37330
rect 253572 37266 253624 37272
rect 253584 29102 253612 37266
rect 253572 29096 253624 29102
rect 253572 29038 253624 29044
rect 253756 29096 253808 29102
rect 253756 29038 253808 29044
rect 253768 27606 253796 29038
rect 253572 27600 253624 27606
rect 253572 27542 253624 27548
rect 253756 27600 253808 27606
rect 253756 27542 253808 27548
rect 253584 18018 253612 27542
rect 253480 18012 253532 18018
rect 253480 17954 253532 17960
rect 253572 18012 253624 18018
rect 253572 17954 253624 17960
rect 253492 9722 253520 17954
rect 253480 9716 253532 9722
rect 253480 9658 253532 9664
rect 253664 9716 253716 9722
rect 253664 9658 253716 9664
rect 251456 4140 251508 4146
rect 251456 4082 251508 4088
rect 252468 4140 252520 4146
rect 252468 4082 252520 4088
rect 252652 4140 252704 4146
rect 252652 4082 252704 4088
rect 251180 3732 251232 3738
rect 251180 3674 251232 3680
rect 250352 3392 250404 3398
rect 250352 3334 250404 3340
rect 251088 3392 251140 3398
rect 251088 3334 251140 3340
rect 250364 480 250392 3334
rect 251468 480 251496 4082
rect 252664 480 252692 4082
rect 253676 4078 253704 9658
rect 253860 4146 253888 118186
rect 253952 118182 253980 120006
rect 254596 118454 254624 120006
rect 255332 118522 255360 120006
rect 255320 118516 255372 118522
rect 255320 118458 255372 118464
rect 254584 118448 254636 118454
rect 254584 118390 254636 118396
rect 255792 118318 255820 120006
rect 256758 119762 256786 120020
rect 256712 119734 256786 119762
rect 256988 120006 257324 120034
rect 257632 120006 257968 120034
rect 258276 120006 258520 120034
rect 258828 120006 259164 120034
rect 259472 120006 259808 120034
rect 260024 120006 260360 120034
rect 260852 120006 261004 120034
rect 261312 120006 261648 120034
rect 256712 118386 256740 119734
rect 256988 118590 257016 120006
rect 256976 118584 257028 118590
rect 256976 118526 257028 118532
rect 256700 118380 256752 118386
rect 256700 118322 256752 118328
rect 255780 118312 255832 118318
rect 255780 118254 255832 118260
rect 256608 118312 256660 118318
rect 256608 118254 256660 118260
rect 253940 118176 253992 118182
rect 253940 118118 253992 118124
rect 255228 118108 255280 118114
rect 255228 118050 255280 118056
rect 253940 115932 253992 115938
rect 253940 115874 253992 115880
rect 253952 106350 253980 115874
rect 253940 106344 253992 106350
rect 253940 106286 253992 106292
rect 253848 4140 253900 4146
rect 253848 4082 253900 4088
rect 253664 4072 253716 4078
rect 253664 4014 253716 4020
rect 253848 4004 253900 4010
rect 253848 3946 253900 3952
rect 253860 480 253888 3946
rect 255240 3346 255268 118050
rect 256620 3346 256648 118254
rect 257632 117910 257660 120006
rect 258276 118658 258304 120006
rect 258264 118652 258316 118658
rect 258264 118594 258316 118600
rect 257988 118176 258040 118182
rect 257988 118118 258040 118124
rect 257620 117904 257672 117910
rect 257620 117846 257672 117852
rect 258000 3534 258028 118118
rect 258828 117638 258856 120006
rect 259472 117706 259500 120006
rect 260024 117842 260052 120006
rect 260748 118380 260800 118386
rect 260748 118322 260800 118328
rect 260012 117836 260064 117842
rect 260012 117778 260064 117784
rect 259460 117700 259512 117706
rect 259460 117642 259512 117648
rect 258816 117632 258868 117638
rect 258816 117574 258868 117580
rect 259276 117632 259328 117638
rect 259276 117574 259328 117580
rect 259288 117366 259316 117574
rect 259276 117360 259328 117366
rect 259276 117302 259328 117308
rect 259368 117360 259420 117366
rect 259368 117302 259420 117308
rect 257436 3528 257488 3534
rect 257436 3470 257488 3476
rect 257988 3528 258040 3534
rect 257988 3470 258040 3476
rect 255056 3318 255268 3346
rect 256252 3318 256648 3346
rect 255056 480 255084 3318
rect 256252 480 256280 3318
rect 257448 480 257476 3470
rect 259380 3126 259408 117302
rect 260760 3534 260788 118322
rect 260852 117774 260880 120006
rect 260840 117768 260892 117774
rect 260840 117710 260892 117716
rect 261312 117570 261340 120006
rect 262186 119762 262214 120020
rect 262508 120006 262844 120034
rect 263152 120006 263488 120034
rect 263704 120006 264040 120034
rect 264348 120006 264684 120034
rect 264992 120006 265328 120034
rect 265544 120006 265880 120034
rect 266372 120006 266524 120034
rect 266832 120006 267168 120034
rect 262186 119734 262260 119762
rect 262128 117768 262180 117774
rect 262128 117710 262180 117716
rect 261300 117564 261352 117570
rect 261300 117506 261352 117512
rect 259828 3528 259880 3534
rect 259828 3470 259880 3476
rect 260748 3528 260800 3534
rect 260748 3470 260800 3476
rect 258632 3120 258684 3126
rect 258632 3062 258684 3068
rect 259368 3120 259420 3126
rect 259368 3062 259420 3068
rect 258644 480 258672 3062
rect 259840 480 259868 3470
rect 262140 3262 262168 117710
rect 262232 117502 262260 119734
rect 262508 117978 262536 120006
rect 262496 117972 262548 117978
rect 262496 117914 262548 117920
rect 263152 117638 263180 120006
rect 263704 118250 263732 120006
rect 263692 118244 263744 118250
rect 263692 118186 263744 118192
rect 264348 118046 264376 120006
rect 264992 118114 265020 120006
rect 265544 118318 265572 120006
rect 265532 118312 265584 118318
rect 265532 118254 265584 118260
rect 266372 118182 266400 120006
rect 266360 118176 266412 118182
rect 266360 118118 266412 118124
rect 264980 118108 265032 118114
rect 264980 118050 265032 118056
rect 264336 118040 264388 118046
rect 264336 117982 264388 117988
rect 266268 118040 266320 118046
rect 266268 117982 266320 117988
rect 264888 117972 264940 117978
rect 264888 117914 264940 117920
rect 263508 117904 263560 117910
rect 263508 117846 263560 117852
rect 263416 117836 263468 117842
rect 263416 117778 263468 117784
rect 263140 117632 263192 117638
rect 263140 117574 263192 117580
rect 262220 117496 262272 117502
rect 262220 117438 262272 117444
rect 262220 3528 262272 3534
rect 262220 3470 262272 3476
rect 261024 3256 261076 3262
rect 261024 3198 261076 3204
rect 262128 3256 262180 3262
rect 262128 3198 262180 3204
rect 261036 480 261064 3198
rect 262232 480 262260 3470
rect 263428 480 263456 117778
rect 263520 3534 263548 117846
rect 263508 3528 263560 3534
rect 264900 3482 264928 117914
rect 266280 3534 266308 117982
rect 266832 117366 266860 120006
rect 267706 119762 267734 120020
rect 268028 120006 268364 120034
rect 268672 120006 269008 120034
rect 269224 120006 269560 120034
rect 269868 120006 270204 120034
rect 270512 120006 270848 120034
rect 271064 120006 271400 120034
rect 271892 120006 272044 120034
rect 272352 120006 272688 120034
rect 267706 119734 267780 119762
rect 267752 118386 267780 119734
rect 267740 118380 267792 118386
rect 267740 118322 267792 118328
rect 267648 118176 267700 118182
rect 267648 118118 267700 118124
rect 266820 117360 266872 117366
rect 266820 117302 266872 117308
rect 263508 3470 263560 3476
rect 264624 3454 264928 3482
rect 265808 3528 265860 3534
rect 265808 3470 265860 3476
rect 266268 3528 266320 3534
rect 266268 3470 266320 3476
rect 264624 480 264652 3454
rect 265820 480 265848 3470
rect 267660 3466 267688 118118
rect 268028 117774 268056 120006
rect 268672 117910 268700 120006
rect 268660 117904 268712 117910
rect 268660 117846 268712 117852
rect 269224 117842 269252 120006
rect 269868 117978 269896 120006
rect 270512 118046 270540 120006
rect 271064 118182 271092 120006
rect 271052 118176 271104 118182
rect 271052 118118 271104 118124
rect 270500 118040 270552 118046
rect 270500 117982 270552 117988
rect 269856 117972 269908 117978
rect 269856 117914 269908 117920
rect 269212 117836 269264 117842
rect 269212 117778 269264 117784
rect 268016 117768 268068 117774
rect 268016 117710 268068 117716
rect 271788 117496 271840 117502
rect 271788 117438 271840 117444
rect 269028 117428 269080 117434
rect 269028 117370 269080 117376
rect 269040 3534 269068 117370
rect 271144 117360 271196 117366
rect 271144 117302 271196 117308
rect 268108 3528 268160 3534
rect 268108 3470 268160 3476
rect 269028 3528 269080 3534
rect 269028 3470 269080 3476
rect 267004 3460 267056 3466
rect 267004 3402 267056 3408
rect 267648 3460 267700 3466
rect 267648 3402 267700 3408
rect 267016 480 267044 3402
rect 268120 480 268148 3470
rect 270500 3460 270552 3466
rect 270500 3402 270552 3408
rect 269304 3052 269356 3058
rect 269304 2994 269356 3000
rect 269316 480 269344 2994
rect 270512 480 270540 3402
rect 271156 3058 271184 117302
rect 271696 3528 271748 3534
rect 271696 3470 271748 3476
rect 271144 3052 271196 3058
rect 271144 2994 271196 3000
rect 271708 480 271736 3470
rect 271800 3466 271828 117438
rect 271892 117434 271920 120006
rect 271880 117428 271932 117434
rect 271880 117370 271932 117376
rect 272352 117366 272380 120006
rect 273226 119762 273254 120020
rect 273548 120006 273884 120034
rect 274192 120006 274528 120034
rect 274652 120006 275080 120034
rect 273226 119734 273300 119762
rect 273272 117502 273300 119734
rect 273260 117496 273312 117502
rect 273260 117438 273312 117444
rect 273548 117434 273576 120006
rect 272524 117428 272576 117434
rect 272524 117370 272576 117376
rect 273536 117428 273588 117434
rect 273536 117370 273588 117376
rect 272340 117360 272392 117366
rect 272340 117302 272392 117308
rect 272536 3534 272564 117370
rect 274192 117366 274220 120006
rect 273168 117360 273220 117366
rect 273168 117302 273220 117308
rect 274180 117360 274232 117366
rect 274652 117314 274680 120006
rect 274180 117302 274232 117308
rect 272524 3528 272576 3534
rect 273180 3482 273208 117302
rect 274560 117286 274680 117314
rect 274456 96620 274508 96626
rect 274456 96562 274508 96568
rect 274468 87009 274496 96562
rect 274454 87000 274510 87009
rect 274454 86935 274510 86944
rect 274560 4146 274588 117286
rect 275204 109154 275232 120142
rect 276262 119762 276290 120020
rect 276920 120006 277348 120034
rect 277564 120006 277900 120034
rect 278116 120006 278636 120034
rect 278760 120006 279096 120034
rect 279404 120006 279740 120034
rect 276216 119734 276290 119762
rect 276216 114578 276244 119734
rect 276112 114572 276164 114578
rect 276112 114514 276164 114520
rect 276204 114572 276256 114578
rect 276204 114514 276256 114520
rect 274928 109126 275232 109154
rect 274928 109018 274956 109126
rect 274836 108990 274956 109018
rect 274836 99498 274864 108990
rect 276124 104854 276152 114514
rect 275928 104848 275980 104854
rect 275928 104790 275980 104796
rect 276112 104848 276164 104854
rect 276112 104790 276164 104796
rect 274836 99470 274956 99498
rect 274928 96801 274956 99470
rect 274914 96792 274970 96801
rect 274914 96727 274970 96736
rect 274730 96656 274786 96665
rect 274730 96591 274732 96600
rect 274784 96591 274786 96600
rect 274732 96562 274784 96568
rect 275940 95266 275968 104790
rect 275928 95260 275980 95266
rect 275928 95202 275980 95208
rect 276020 95260 276072 95266
rect 276020 95202 276072 95208
rect 276032 95130 276060 95202
rect 276020 95124 276072 95130
rect 276020 95066 276072 95072
rect 276296 95124 276348 95130
rect 276296 95066 276348 95072
rect 274638 87000 274694 87009
rect 274638 86935 274640 86944
rect 274692 86935 274694 86944
rect 274824 86964 274876 86970
rect 274640 86906 274692 86912
rect 274824 86906 274876 86912
rect 274836 79914 274864 86906
rect 276308 85649 276336 95066
rect 276110 85640 276166 85649
rect 276110 85575 276166 85584
rect 276294 85640 276350 85649
rect 276294 85575 276350 85584
rect 276124 85542 276152 85575
rect 276112 85536 276164 85542
rect 276112 85478 276164 85484
rect 276204 85536 276256 85542
rect 276204 85478 276256 85484
rect 276216 84182 276244 85478
rect 276020 84176 276072 84182
rect 276020 84118 276072 84124
rect 276204 84176 276256 84182
rect 276204 84118 276256 84124
rect 274744 79886 274864 79914
rect 274744 72486 274772 79886
rect 276032 74594 276060 84118
rect 275928 74588 275980 74594
rect 275928 74530 275980 74536
rect 276020 74588 276072 74594
rect 276020 74530 276072 74536
rect 274732 72480 274784 72486
rect 274732 72422 274784 72428
rect 275100 72480 275152 72486
rect 275100 72422 275152 72428
rect 275112 67658 275140 72422
rect 274916 67652 274968 67658
rect 274916 67594 274968 67600
rect 275100 67652 275152 67658
rect 275100 67594 275152 67600
rect 274928 60738 274956 67594
rect 275940 67402 275968 74530
rect 275940 67374 276152 67402
rect 274744 60710 274956 60738
rect 274744 53174 274772 60710
rect 276124 57934 276152 67374
rect 276112 57928 276164 57934
rect 276112 57870 276164 57876
rect 276204 57928 276256 57934
rect 276204 57870 276256 57876
rect 274732 53168 274784 53174
rect 274732 53110 274784 53116
rect 275100 53168 275152 53174
rect 275100 53110 275152 53116
rect 275112 48346 275140 53110
rect 276216 48414 276244 57870
rect 276112 48408 276164 48414
rect 276112 48350 276164 48356
rect 276204 48408 276256 48414
rect 276204 48350 276256 48356
rect 274916 48340 274968 48346
rect 274916 48282 274968 48288
rect 275100 48340 275152 48346
rect 275100 48282 275152 48288
rect 274928 41426 274956 48282
rect 276124 46918 276152 48350
rect 276112 46912 276164 46918
rect 276112 46854 276164 46860
rect 276204 46912 276256 46918
rect 276204 46854 276256 46860
rect 274744 41398 274956 41426
rect 274744 38622 274772 41398
rect 274732 38616 274784 38622
rect 274732 38558 274784 38564
rect 275100 38616 275152 38622
rect 275100 38558 275152 38564
rect 275112 29034 275140 38558
rect 276216 29102 276244 46854
rect 276112 29096 276164 29102
rect 276112 29038 276164 29044
rect 276204 29096 276256 29102
rect 276204 29038 276256 29044
rect 274916 29028 274968 29034
rect 274916 28970 274968 28976
rect 275100 29028 275152 29034
rect 275100 28970 275152 28976
rect 274928 22114 274956 28970
rect 276124 27606 276152 29038
rect 275928 27600 275980 27606
rect 275928 27542 275980 27548
rect 276112 27600 276164 27606
rect 276112 27542 276164 27548
rect 274744 22086 274956 22114
rect 274744 14634 274772 22086
rect 275940 18018 275968 27542
rect 275928 18012 275980 18018
rect 275928 17954 275980 17960
rect 276112 18012 276164 18018
rect 276112 17954 276164 17960
rect 274744 14606 275048 14634
rect 275020 9722 275048 14606
rect 276124 12510 276152 17954
rect 276112 12504 276164 12510
rect 276112 12446 276164 12452
rect 276480 12368 276532 12374
rect 276480 12310 276532 12316
rect 275008 9716 275060 9722
rect 275008 9658 275060 9664
rect 275284 9716 275336 9722
rect 275284 9658 275336 9664
rect 275296 9602 275324 9658
rect 275296 9574 275416 9602
rect 274088 4140 274140 4146
rect 274088 4082 274140 4088
rect 274548 4140 274600 4146
rect 274548 4082 274600 4088
rect 272524 3470 272576 3476
rect 271788 3460 271840 3466
rect 271788 3402 271840 3408
rect 272904 3454 273208 3482
rect 272904 480 272932 3454
rect 274100 480 274128 4082
rect 275388 610 275416 9574
rect 275284 604 275336 610
rect 275284 546 275336 552
rect 275376 604 275428 610
rect 275376 546 275428 552
rect 275296 480 275324 546
rect 276492 480 276520 12310
rect 277320 4146 277348 120006
rect 277872 117774 277900 120006
rect 277860 117768 277912 117774
rect 277860 117710 277912 117716
rect 278608 4146 278636 120006
rect 279068 117978 279096 120006
rect 279056 117972 279108 117978
rect 279056 117914 279108 117920
rect 278688 117768 278740 117774
rect 278688 117710 278740 117716
rect 278700 4162 278728 117710
rect 279712 117366 279740 120006
rect 279942 119762 279970 120020
rect 280600 120006 280936 120034
rect 281244 120006 281396 120034
rect 281796 120006 282132 120034
rect 282440 120006 282776 120034
rect 283084 120006 283420 120034
rect 283636 120006 284156 120034
rect 284280 120006 284616 120034
rect 284924 120006 285260 120034
rect 279942 119734 280016 119762
rect 279700 117360 279752 117366
rect 279700 117302 279752 117308
rect 279988 11370 280016 119734
rect 280908 117978 280936 120006
rect 280344 117972 280396 117978
rect 280344 117914 280396 117920
rect 280896 117972 280948 117978
rect 280896 117914 280948 117920
rect 280068 117360 280120 117366
rect 280068 117302 280120 117308
rect 279804 11342 280016 11370
rect 277308 4140 277360 4146
rect 277308 4082 277360 4088
rect 277676 4140 277728 4146
rect 277676 4082 277728 4088
rect 278596 4140 278648 4146
rect 278700 4134 278912 4162
rect 278596 4082 278648 4088
rect 277688 480 277716 4082
rect 278884 480 278912 4134
rect 279804 3602 279832 11342
rect 280080 11234 280108 117302
rect 279988 11206 280108 11234
rect 279988 4078 280016 11206
rect 280068 4140 280120 4146
rect 280068 4082 280120 4088
rect 279976 4072 280028 4078
rect 279976 4014 280028 4020
rect 279792 3596 279844 3602
rect 279792 3538 279844 3544
rect 280080 480 280108 4082
rect 280356 610 280384 117914
rect 281368 3194 281396 120006
rect 281448 117972 281500 117978
rect 281448 117914 281500 117920
rect 281460 3534 281488 117914
rect 282104 117366 282132 120006
rect 282092 117360 282144 117366
rect 282092 117302 282144 117308
rect 282460 4072 282512 4078
rect 282460 4014 282512 4020
rect 281448 3528 281500 3534
rect 281448 3470 281500 3476
rect 281356 3188 281408 3194
rect 281356 3130 281408 3136
rect 280344 604 280396 610
rect 280344 546 280396 552
rect 281264 604 281316 610
rect 281264 546 281316 552
rect 281276 480 281304 546
rect 282472 480 282500 4014
rect 282748 3330 282776 120006
rect 283392 117366 283420 120006
rect 282828 117360 282880 117366
rect 282828 117302 282880 117308
rect 283380 117360 283432 117366
rect 283380 117302 283432 117308
rect 284024 117360 284076 117366
rect 284024 117302 284076 117308
rect 282840 3398 282868 117302
rect 284036 116498 284064 117302
rect 284128 116634 284156 120006
rect 284588 117434 284616 120006
rect 284576 117428 284628 117434
rect 284576 117370 284628 117376
rect 285232 117366 285260 120006
rect 285462 119762 285490 120020
rect 286120 120006 286456 120034
rect 286764 120006 286916 120034
rect 287316 120006 287652 120034
rect 287960 120006 288296 120034
rect 288604 120006 288940 120034
rect 289156 120006 289676 120034
rect 289800 120006 290136 120034
rect 290444 120006 290872 120034
rect 290996 120006 291148 120034
rect 291640 120006 291976 120034
rect 292284 120006 292528 120034
rect 292836 120006 293172 120034
rect 293480 120006 293908 120034
rect 294032 120006 294368 120034
rect 294676 120006 295012 120034
rect 295320 120006 295656 120034
rect 295872 120006 296208 120034
rect 285416 119734 285490 119762
rect 285220 117360 285272 117366
rect 285220 117302 285272 117308
rect 284128 116606 284248 116634
rect 284036 116470 284156 116498
rect 284128 4146 284156 116470
rect 284116 4140 284168 4146
rect 284116 4082 284168 4088
rect 284220 3670 284248 116606
rect 284208 3664 284260 3670
rect 284208 3606 284260 3612
rect 283656 3596 283708 3602
rect 283656 3538 283708 3544
rect 282828 3392 282880 3398
rect 282828 3334 282880 3340
rect 282736 3324 282788 3330
rect 282736 3266 282788 3272
rect 283668 480 283696 3538
rect 285416 3534 285444 119734
rect 285496 117428 285548 117434
rect 285496 117370 285548 117376
rect 284760 3528 284812 3534
rect 284760 3470 284812 3476
rect 285404 3528 285456 3534
rect 285404 3470 285456 3476
rect 284772 480 284800 3470
rect 285508 3466 285536 117370
rect 286428 117366 286456 120006
rect 285588 117360 285640 117366
rect 285588 117302 285640 117308
rect 286416 117360 286468 117366
rect 286416 117302 286468 117308
rect 285600 3874 285628 117302
rect 285588 3868 285640 3874
rect 285588 3810 285640 3816
rect 286888 3602 286916 120006
rect 287624 117366 287652 120006
rect 286968 117360 287020 117366
rect 286968 117302 287020 117308
rect 287612 117360 287664 117366
rect 287612 117302 287664 117308
rect 286980 4010 287008 117302
rect 286968 4004 287020 4010
rect 286968 3946 287020 3952
rect 288268 3806 288296 120006
rect 288912 117366 288940 120006
rect 288348 117360 288400 117366
rect 288348 117302 288400 117308
rect 288900 117360 288952 117366
rect 288900 117302 288952 117308
rect 289544 117360 289596 117366
rect 289544 117302 289596 117308
rect 288256 3800 288308 3806
rect 288256 3742 288308 3748
rect 286876 3596 286928 3602
rect 286876 3538 286928 3544
rect 285496 3460 285548 3466
rect 285496 3402 285548 3408
rect 287152 3392 287204 3398
rect 287152 3334 287204 3340
rect 285956 3188 286008 3194
rect 285956 3130 286008 3136
rect 285968 480 285996 3130
rect 287164 480 287192 3334
rect 288360 3330 288388 117302
rect 289556 116498 289584 117302
rect 289648 116634 289676 120006
rect 290108 117366 290136 120006
rect 290096 117360 290148 117366
rect 290096 117302 290148 117308
rect 290740 117360 290792 117366
rect 290740 117302 290792 117308
rect 289648 116606 289768 116634
rect 289556 116470 289676 116498
rect 289544 4140 289596 4146
rect 289544 4082 289596 4088
rect 288348 3324 288400 3330
rect 288348 3266 288400 3272
rect 288348 3188 288400 3194
rect 288348 3130 288400 3136
rect 288360 480 288388 3130
rect 289556 480 289584 4082
rect 289648 3398 289676 116470
rect 289740 4146 289768 116606
rect 290752 116498 290780 117302
rect 290844 116634 290872 120006
rect 291120 118182 291148 120006
rect 291108 118176 291160 118182
rect 291108 118118 291160 118124
rect 291948 117366 291976 120006
rect 291936 117360 291988 117366
rect 291936 117302 291988 117308
rect 292396 117360 292448 117366
rect 292396 117302 292448 117308
rect 290844 116606 291148 116634
rect 290752 116470 291056 116498
rect 289728 4140 289780 4146
rect 289728 4082 289780 4088
rect 291028 3738 291056 116470
rect 291120 4078 291148 116606
rect 291108 4072 291160 4078
rect 291108 4014 291160 4020
rect 291016 3732 291068 3738
rect 291016 3674 291068 3680
rect 292408 3670 292436 117302
rect 290740 3664 290792 3670
rect 290740 3606 290792 3612
rect 292396 3664 292448 3670
rect 292396 3606 292448 3612
rect 289636 3392 289688 3398
rect 289636 3334 289688 3340
rect 290752 480 290780 3606
rect 292500 3466 292528 120006
rect 293144 118114 293172 120006
rect 293132 118108 293184 118114
rect 293132 118050 293184 118056
rect 293880 3942 293908 120006
rect 294340 117366 294368 120006
rect 294984 118046 295012 120006
rect 294972 118040 295024 118046
rect 294972 117982 295024 117988
rect 295628 117366 295656 120006
rect 296180 117842 296208 120006
rect 296502 119762 296530 120020
rect 297160 120006 297496 120034
rect 297712 120006 298048 120034
rect 298356 120006 298692 120034
rect 299000 120006 299336 120034
rect 299552 120006 299888 120034
rect 300196 120006 300532 120034
rect 300840 120006 301176 120034
rect 301392 120006 301728 120034
rect 302036 120006 302188 120034
rect 302680 120006 303016 120034
rect 303232 120006 303476 120034
rect 303876 120006 304212 120034
rect 304520 120006 304948 120034
rect 305072 120006 305408 120034
rect 305716 120006 306052 120034
rect 306360 120006 306696 120034
rect 306912 120006 307248 120034
rect 307556 120006 307708 120034
rect 308200 120006 308536 120034
rect 308752 120006 309088 120034
rect 309396 120006 309732 120034
rect 310040 120006 310468 120034
rect 310592 120006 310928 120034
rect 311236 120006 311572 120034
rect 296502 119734 296576 119762
rect 296548 117910 296576 119734
rect 296536 117904 296588 117910
rect 296536 117846 296588 117852
rect 296168 117836 296220 117842
rect 296168 117778 296220 117784
rect 297468 117366 297496 120006
rect 294328 117360 294380 117366
rect 294328 117302 294380 117308
rect 295248 117360 295300 117366
rect 295248 117302 295300 117308
rect 295616 117360 295668 117366
rect 295616 117302 295668 117308
rect 296628 117360 296680 117366
rect 296628 117302 296680 117308
rect 297456 117360 297508 117366
rect 297456 117302 297508 117308
rect 297916 117360 297968 117366
rect 297916 117302 297968 117308
rect 293868 3936 293920 3942
rect 293868 3878 293920 3884
rect 295260 3874 295288 117302
rect 295524 4004 295576 4010
rect 295524 3946 295576 3952
rect 293132 3868 293184 3874
rect 293132 3810 293184 3816
rect 295248 3868 295300 3874
rect 295248 3810 295300 3816
rect 291936 3460 291988 3466
rect 291936 3402 291988 3408
rect 292488 3460 292540 3466
rect 292488 3402 292540 3408
rect 291948 480 291976 3402
rect 293144 480 293172 3810
rect 294328 3528 294380 3534
rect 294328 3470 294380 3476
rect 294340 480 294368 3470
rect 295536 480 295564 3946
rect 296640 3534 296668 117302
rect 297928 4010 297956 117302
rect 297916 4004 297968 4010
rect 297916 3946 297968 3952
rect 298020 3602 298048 120006
rect 298664 118658 298692 120006
rect 298652 118652 298704 118658
rect 298652 118594 298704 118600
rect 299308 118522 299336 120006
rect 299296 118516 299348 118522
rect 299296 118458 299348 118464
rect 299860 117366 299888 120006
rect 300504 118250 300532 120006
rect 301148 118590 301176 120006
rect 301136 118584 301188 118590
rect 301136 118526 301188 118532
rect 300492 118244 300544 118250
rect 300492 118186 300544 118192
rect 301700 117366 301728 120006
rect 302160 118454 302188 120006
rect 302148 118448 302200 118454
rect 302148 118390 302200 118396
rect 302988 117366 303016 120006
rect 303448 117434 303476 120006
rect 304184 118386 304212 120006
rect 304172 118380 304224 118386
rect 304172 118322 304224 118328
rect 303436 117428 303488 117434
rect 303436 117370 303488 117376
rect 299848 117360 299900 117366
rect 299848 117302 299900 117308
rect 300768 117360 300820 117366
rect 300768 117302 300820 117308
rect 301688 117360 301740 117366
rect 301688 117302 301740 117308
rect 302884 117360 302936 117366
rect 302884 117302 302936 117308
rect 302976 117360 303028 117366
rect 302976 117302 303028 117308
rect 303528 117360 303580 117366
rect 303528 117302 303580 117308
rect 299112 3800 299164 3806
rect 299112 3742 299164 3748
rect 296720 3596 296772 3602
rect 296720 3538 296772 3544
rect 298008 3596 298060 3602
rect 298008 3538 298060 3544
rect 296628 3528 296680 3534
rect 296628 3470 296680 3476
rect 296732 480 296760 3538
rect 297916 3324 297968 3330
rect 297916 3266 297968 3272
rect 297928 480 297956 3266
rect 299124 480 299152 3742
rect 300780 3398 300808 117302
rect 301412 4140 301464 4146
rect 301412 4082 301464 4088
rect 300308 3392 300360 3398
rect 300308 3334 300360 3340
rect 300768 3392 300820 3398
rect 300768 3334 300820 3340
rect 300320 480 300348 3334
rect 301424 480 301452 4082
rect 302896 3806 302924 117302
rect 303540 5234 303568 117302
rect 303528 5228 303580 5234
rect 303528 5170 303580 5176
rect 304920 5098 304948 120006
rect 305184 118176 305236 118182
rect 305184 118118 305236 118124
rect 304908 5092 304960 5098
rect 304908 5034 304960 5040
rect 303804 4072 303856 4078
rect 303804 4014 303856 4020
rect 302884 3800 302936 3806
rect 302884 3742 302936 3748
rect 302608 3732 302660 3738
rect 302608 3674 302660 3680
rect 302620 480 302648 3674
rect 303816 480 303844 4014
rect 305196 610 305224 118118
rect 305380 117706 305408 120006
rect 306024 118318 306052 120006
rect 306012 118312 306064 118318
rect 306012 118254 306064 118260
rect 305368 117700 305420 117706
rect 305368 117642 305420 117648
rect 305644 117428 305696 117434
rect 305644 117370 305696 117376
rect 305656 3670 305684 117370
rect 306668 117366 306696 120006
rect 307220 117570 307248 120006
rect 307680 118250 307708 120006
rect 307668 118244 307720 118250
rect 307668 118186 307720 118192
rect 307944 118108 307996 118114
rect 307944 118050 307996 118056
rect 307208 117564 307260 117570
rect 307208 117506 307260 117512
rect 306656 117360 306708 117366
rect 306656 117302 306708 117308
rect 307668 117360 307720 117366
rect 307668 117302 307720 117308
rect 307680 5166 307708 117302
rect 307668 5160 307720 5166
rect 307668 5102 307720 5108
rect 306196 3732 306248 3738
rect 306196 3674 306248 3680
rect 305644 3664 305696 3670
rect 305644 3606 305696 3612
rect 305000 604 305052 610
rect 305000 546 305052 552
rect 305184 604 305236 610
rect 305184 546 305236 552
rect 305012 480 305040 546
rect 306208 480 306236 3674
rect 307392 3460 307444 3466
rect 307392 3402 307444 3408
rect 307404 480 307432 3402
rect 307956 610 307984 118050
rect 308508 117638 308536 120006
rect 308496 117632 308548 117638
rect 308496 117574 308548 117580
rect 308956 117632 309008 117638
rect 308956 117574 309008 117580
rect 308968 5030 308996 117574
rect 308956 5024 309008 5030
rect 308956 4966 309008 4972
rect 309060 3262 309088 120006
rect 309704 117570 309732 120006
rect 309692 117564 309744 117570
rect 309692 117506 309744 117512
rect 310440 4962 310468 120006
rect 310900 117434 310928 120006
rect 311544 117638 311572 120006
rect 311774 119762 311802 120020
rect 312432 120006 312768 120034
rect 313076 120006 313228 120034
rect 313628 120006 313964 120034
rect 314272 120006 314608 120034
rect 314916 120006 315252 120034
rect 315468 120006 315896 120034
rect 316112 120006 316448 120034
rect 311774 119734 311848 119762
rect 311532 117632 311584 117638
rect 311532 117574 311584 117580
rect 310888 117428 310940 117434
rect 310888 117370 310940 117376
rect 310428 4956 310480 4962
rect 310428 4898 310480 4904
rect 311820 4894 311848 119734
rect 311900 117904 311952 117910
rect 311900 117846 311952 117852
rect 311808 4888 311860 4894
rect 311808 4830 311860 4836
rect 309784 3936 309836 3942
rect 309784 3878 309836 3884
rect 309600 3800 309652 3806
rect 309600 3742 309652 3748
rect 309612 3398 309640 3742
rect 309600 3392 309652 3398
rect 309600 3334 309652 3340
rect 309048 3256 309100 3262
rect 309048 3198 309100 3204
rect 307944 604 307996 610
rect 307944 546 307996 552
rect 308588 604 308640 610
rect 308588 546 308640 552
rect 308600 480 308628 546
rect 309796 480 309824 3878
rect 310980 3868 311032 3874
rect 310980 3810 311032 3816
rect 310992 480 311020 3810
rect 311912 626 311940 117846
rect 312740 117706 312768 120006
rect 313200 118046 313228 120006
rect 313188 118040 313240 118046
rect 313188 117982 313240 117988
rect 312636 117700 312688 117706
rect 312636 117642 312688 117648
rect 312728 117700 312780 117706
rect 312728 117642 312780 117648
rect 312544 117360 312596 117366
rect 312544 117302 312596 117308
rect 312556 4146 312584 117302
rect 312544 4140 312596 4146
rect 312544 4082 312596 4088
rect 312648 3942 312676 117642
rect 313936 117366 313964 120006
rect 314580 117910 314608 120006
rect 314568 117904 314620 117910
rect 314568 117846 314620 117852
rect 315224 117774 315252 120006
rect 314660 117768 314712 117774
rect 314660 117710 314712 117716
rect 315212 117768 315264 117774
rect 315212 117710 315264 117716
rect 314108 117496 314160 117502
rect 314108 117438 314160 117444
rect 313924 117360 313976 117366
rect 313924 117302 313976 117308
rect 314120 115954 314148 117438
rect 314568 117360 314620 117366
rect 314568 117302 314620 117308
rect 314028 115938 314148 115954
rect 314016 115932 314160 115938
rect 314068 115926 314108 115932
rect 314016 115874 314068 115880
rect 314108 115874 314160 115880
rect 314028 115843 314056 115874
rect 314120 109070 314148 115874
rect 314108 109064 314160 109070
rect 314108 109006 314160 109012
rect 314016 108996 314068 109002
rect 314016 108938 314068 108944
rect 314028 106298 314056 108938
rect 314028 106270 314148 106298
rect 314120 99414 314148 106270
rect 313924 99408 313976 99414
rect 313924 99350 313976 99356
rect 314108 99408 314160 99414
rect 314108 99350 314160 99356
rect 313936 85542 313964 99350
rect 313924 85536 313976 85542
rect 313924 85478 313976 85484
rect 314016 85536 314068 85542
rect 314016 85478 314068 85484
rect 314028 84182 314056 85478
rect 314016 84176 314068 84182
rect 314016 84118 314068 84124
rect 314200 84176 314252 84182
rect 314200 84118 314252 84124
rect 314212 67402 314240 84118
rect 314028 67374 314240 67402
rect 314028 58002 314056 67374
rect 314016 57996 314068 58002
rect 314016 57938 314068 57944
rect 314016 57860 314068 57866
rect 314016 57802 314068 57808
rect 314028 51134 314056 57802
rect 314016 51128 314068 51134
rect 314016 51070 314068 51076
rect 314016 50992 314068 50998
rect 314016 50934 314068 50940
rect 314028 43518 314056 50934
rect 313740 43512 313792 43518
rect 313740 43454 313792 43460
rect 314016 43512 314068 43518
rect 314016 43454 314068 43460
rect 313752 38690 313780 43454
rect 313740 38684 313792 38690
rect 313740 38626 313792 38632
rect 313924 38684 313976 38690
rect 313924 38626 313976 38632
rect 313936 28898 313964 38626
rect 313648 28892 313700 28898
rect 313648 28834 313700 28840
rect 313924 28892 313976 28898
rect 313924 28834 313976 28840
rect 313660 19378 313688 28834
rect 313648 19372 313700 19378
rect 313648 19314 313700 19320
rect 313924 19372 313976 19378
rect 313924 19314 313976 19320
rect 312636 3936 312688 3942
rect 312636 3878 312688 3884
rect 313936 3874 313964 19314
rect 314580 4826 314608 117302
rect 314672 12442 314700 117710
rect 315304 117428 315356 117434
rect 315304 117370 315356 117376
rect 314660 12436 314712 12442
rect 314660 12378 314712 12384
rect 314568 4820 314620 4826
rect 314568 4762 314620 4768
rect 314568 4140 314620 4146
rect 314568 4082 314620 4088
rect 313924 3868 313976 3874
rect 313924 3810 313976 3816
rect 313372 3460 313424 3466
rect 313372 3402 313424 3408
rect 311912 598 312216 626
rect 312188 480 312216 598
rect 313384 480 313412 3402
rect 314580 480 314608 4082
rect 315316 3534 315344 117370
rect 315764 12436 315816 12442
rect 315764 12378 315816 12384
rect 315304 3528 315356 3534
rect 315304 3470 315356 3476
rect 315776 480 315804 12378
rect 315868 5846 315896 120006
rect 316420 117842 316448 120006
rect 316684 118176 316736 118182
rect 316684 118118 316736 118124
rect 316592 118108 316644 118114
rect 316592 118050 316644 118056
rect 316408 117836 316460 117842
rect 316408 117778 316460 117784
rect 315948 117768 316000 117774
rect 315948 117710 316000 117716
rect 315960 6594 315988 117710
rect 316604 117638 316632 118050
rect 316592 117632 316644 117638
rect 316592 117574 316644 117580
rect 316696 117570 316724 118118
rect 316684 117564 316736 117570
rect 316684 117506 316736 117512
rect 317064 111058 317092 120142
rect 317294 119762 317322 120020
rect 317952 120006 318288 120034
rect 317294 119734 317368 119762
rect 317064 111030 317276 111058
rect 317248 106418 317276 111030
rect 317052 106412 317104 106418
rect 317052 106354 317104 106360
rect 317236 106412 317288 106418
rect 317236 106354 317288 106360
rect 317064 104854 317092 106354
rect 316868 104848 316920 104854
rect 316868 104790 316920 104796
rect 317052 104848 317104 104854
rect 317052 104790 317104 104796
rect 316880 95266 316908 104790
rect 316868 95260 316920 95266
rect 316868 95202 316920 95208
rect 317052 95260 317104 95266
rect 317052 95202 317104 95208
rect 317064 86986 317092 95202
rect 317064 86970 317184 86986
rect 316960 86964 317012 86970
rect 317064 86964 317196 86970
rect 317064 86958 317144 86964
rect 316960 86906 317012 86912
rect 317144 86906 317196 86912
rect 316972 77314 317000 86906
rect 316960 77308 317012 77314
rect 316960 77250 317012 77256
rect 317236 77308 317288 77314
rect 317236 77250 317288 77256
rect 317248 70394 317276 77250
rect 317156 70366 317276 70394
rect 317156 60738 317184 70366
rect 317156 60710 317276 60738
rect 317248 48346 317276 60710
rect 317144 48340 317196 48346
rect 317144 48282 317196 48288
rect 317236 48340 317288 48346
rect 317236 48282 317288 48288
rect 317156 41426 317184 48282
rect 317156 41398 317276 41426
rect 317248 29034 317276 41398
rect 317144 29028 317196 29034
rect 317144 28970 317196 28976
rect 317236 29028 317288 29034
rect 317236 28970 317288 28976
rect 317156 22114 317184 28970
rect 317156 22086 317276 22114
rect 317248 12458 317276 22086
rect 317064 12430 317276 12458
rect 315948 6588 316000 6594
rect 315948 6530 316000 6536
rect 317064 5914 317092 12430
rect 317340 6050 317368 119734
rect 318260 117366 318288 120006
rect 318582 119762 318610 120020
rect 319148 120006 319484 120034
rect 319792 120006 320128 120034
rect 320436 120006 320772 120034
rect 320988 120006 321508 120034
rect 321632 120006 321968 120034
rect 322276 120006 322612 120034
rect 318582 119734 318656 119762
rect 318248 117360 318300 117366
rect 318248 117302 318300 117308
rect 318628 6118 318656 119734
rect 318984 118652 319036 118658
rect 318984 118594 319036 118600
rect 318708 117360 318760 117366
rect 318708 117302 318760 117308
rect 318616 6112 318668 6118
rect 318616 6054 318668 6060
rect 317328 6044 317380 6050
rect 317328 5986 317380 5992
rect 317052 5908 317104 5914
rect 317052 5850 317104 5856
rect 315856 5840 315908 5846
rect 315856 5782 315908 5788
rect 316960 4004 317012 4010
rect 316960 3946 317012 3952
rect 316972 480 317000 3946
rect 318720 3602 318748 117302
rect 318064 3596 318116 3602
rect 318064 3538 318116 3544
rect 318708 3596 318760 3602
rect 318708 3538 318760 3544
rect 318076 480 318104 3538
rect 318996 592 319024 118594
rect 319352 117700 319404 117706
rect 319352 117642 319404 117648
rect 319364 117178 319392 117642
rect 319456 117366 319484 120006
rect 320100 117706 320128 120006
rect 320364 118516 320416 118522
rect 320364 118458 320416 118464
rect 320088 117700 320140 117706
rect 320088 117642 320140 117648
rect 319444 117360 319496 117366
rect 319444 117302 319496 117308
rect 320088 117360 320140 117366
rect 320088 117302 320140 117308
rect 319364 117150 319484 117178
rect 319456 3262 319484 117150
rect 320100 5982 320128 117302
rect 320088 5976 320140 5982
rect 320088 5918 320140 5924
rect 319444 3256 319496 3262
rect 319444 3198 319496 3204
rect 320376 592 320404 118458
rect 320744 117774 320772 120006
rect 320732 117768 320784 117774
rect 320732 117710 320784 117716
rect 321376 117768 321428 117774
rect 321376 117710 321428 117716
rect 321388 6866 321416 117710
rect 321376 6860 321428 6866
rect 321376 6802 321428 6808
rect 321480 6798 321508 120006
rect 321744 117972 321796 117978
rect 321744 117914 321796 117920
rect 321468 6792 321520 6798
rect 321468 6734 321520 6740
rect 321652 3800 321704 3806
rect 321652 3742 321704 3748
rect 318996 564 319300 592
rect 320376 564 320496 592
rect 319272 480 319300 564
rect 320468 480 320496 564
rect 321664 480 321692 3742
rect 321756 2802 321784 117914
rect 321940 117774 321968 120006
rect 322204 117904 322256 117910
rect 322204 117846 322256 117852
rect 321928 117768 321980 117774
rect 321928 117710 321980 117716
rect 322216 3194 322244 117846
rect 322584 117366 322612 120006
rect 322814 119762 322842 120020
rect 323472 120006 323808 120034
rect 322768 119734 322842 119762
rect 322572 117360 322624 117366
rect 322572 117302 322624 117308
rect 322768 6662 322796 119734
rect 323124 118584 323176 118590
rect 323124 118526 323176 118532
rect 322848 117360 322900 117366
rect 322848 117302 322900 117308
rect 322756 6656 322808 6662
rect 322756 6598 322808 6604
rect 322860 4282 322888 117302
rect 322848 4276 322900 4282
rect 322848 4218 322900 4224
rect 322204 3188 322256 3194
rect 322204 3130 322256 3136
rect 321756 2774 322888 2802
rect 322860 480 322888 2774
rect 323136 610 323164 118526
rect 323780 117366 323808 120006
rect 324102 119762 324130 120020
rect 324668 120006 325004 120034
rect 325312 120006 325648 120034
rect 325956 120006 326292 120034
rect 326508 120006 326936 120034
rect 327152 120006 327488 120034
rect 327796 120006 328132 120034
rect 324102 119734 324176 119762
rect 323768 117360 323820 117366
rect 323768 117302 323820 117308
rect 324148 4350 324176 119734
rect 324976 117366 325004 120006
rect 324228 117360 324280 117366
rect 324228 117302 324280 117308
rect 324964 117360 325016 117366
rect 324964 117302 325016 117308
rect 325516 117360 325568 117366
rect 325516 117302 325568 117308
rect 324136 4344 324188 4350
rect 324136 4286 324188 4292
rect 324240 4146 324268 117302
rect 325528 6526 325556 117302
rect 325516 6520 325568 6526
rect 325516 6462 325568 6468
rect 324228 4140 324280 4146
rect 324228 4082 324280 4088
rect 325620 4078 325648 120006
rect 325884 118448 325936 118454
rect 325884 118390 325936 118396
rect 325608 4072 325660 4078
rect 325608 4014 325660 4020
rect 325240 3732 325292 3738
rect 325240 3674 325292 3680
rect 323124 604 323176 610
rect 323124 546 323176 552
rect 324044 604 324096 610
rect 324044 546 324096 552
rect 324056 480 324084 546
rect 325252 480 325280 3674
rect 325896 610 325924 118390
rect 326264 117366 326292 120006
rect 326252 117360 326304 117366
rect 326252 117302 326304 117308
rect 326908 6458 326936 120006
rect 327460 117502 327488 120006
rect 327448 117496 327500 117502
rect 327448 117438 327500 117444
rect 328104 117366 328132 120006
rect 328334 119762 328362 120020
rect 328992 120006 329328 120034
rect 329544 120006 329696 120034
rect 330188 120006 330524 120034
rect 330832 120006 331168 120034
rect 331384 120006 331720 120034
rect 332028 120006 332456 120034
rect 332672 120006 333008 120034
rect 333224 120006 333560 120034
rect 328288 119734 328362 119762
rect 326988 117360 327040 117366
rect 326988 117302 327040 117308
rect 328092 117360 328144 117366
rect 328092 117302 328144 117308
rect 326896 6452 326948 6458
rect 326896 6394 326948 6400
rect 327000 4418 327028 117302
rect 328288 6390 328316 119734
rect 329300 117366 329328 120006
rect 328368 117360 328420 117366
rect 328368 117302 328420 117308
rect 329288 117360 329340 117366
rect 329288 117302 329340 117308
rect 328276 6384 328328 6390
rect 328276 6326 328328 6332
rect 327632 5228 327684 5234
rect 327632 5170 327684 5176
rect 326988 4412 327040 4418
rect 326988 4354 327040 4360
rect 325884 604 325936 610
rect 325884 546 325936 552
rect 326436 604 326488 610
rect 326436 546 326488 552
rect 326448 480 326476 546
rect 327644 480 327672 5170
rect 328380 4486 328408 117302
rect 329668 4622 329696 120006
rect 330024 118380 330076 118386
rect 330024 118322 330076 118328
rect 329748 117360 329800 117366
rect 329748 117302 329800 117308
rect 329656 4616 329708 4622
rect 329656 4558 329708 4564
rect 328368 4480 328420 4486
rect 328368 4422 328420 4428
rect 329760 4010 329788 117302
rect 329748 4004 329800 4010
rect 329748 3946 329800 3952
rect 328828 3664 328880 3670
rect 328828 3606 328880 3612
rect 328840 480 328868 3606
rect 330036 480 330064 118322
rect 330496 117366 330524 120006
rect 331140 117842 331168 120006
rect 331128 117836 331180 117842
rect 331128 117778 331180 117784
rect 331692 117366 331720 120006
rect 331864 117904 331916 117910
rect 331864 117846 331916 117852
rect 330484 117360 330536 117366
rect 330484 117302 330536 117308
rect 331128 117360 331180 117366
rect 331128 117302 331180 117308
rect 331680 117360 331732 117366
rect 331680 117302 331732 117308
rect 331140 6322 331168 117302
rect 331128 6316 331180 6322
rect 331128 6258 331180 6264
rect 331220 5092 331272 5098
rect 331220 5034 331272 5040
rect 331232 480 331260 5034
rect 331876 3126 331904 117846
rect 331956 117632 332008 117638
rect 331956 117574 332008 117580
rect 331968 3330 331996 117574
rect 332428 6254 332456 120006
rect 332876 118312 332928 118318
rect 332876 118254 332928 118260
rect 332508 117360 332560 117366
rect 332508 117302 332560 117308
rect 332416 6248 332468 6254
rect 332416 6190 332468 6196
rect 332520 4554 332548 117302
rect 332508 4548 332560 4554
rect 332508 4490 332560 4496
rect 332416 3936 332468 3942
rect 332416 3878 332468 3884
rect 331956 3324 332008 3330
rect 331956 3266 332008 3272
rect 331864 3120 331916 3126
rect 331864 3062 331916 3068
rect 332428 480 332456 3878
rect 332888 610 332916 118254
rect 332980 117434 333008 120006
rect 332968 117428 333020 117434
rect 332968 117370 333020 117376
rect 333532 117366 333560 120006
rect 333716 120006 333868 120034
rect 334512 120006 334848 120034
rect 335064 120006 335308 120034
rect 335708 120006 336044 120034
rect 336352 120006 336688 120034
rect 336904 120006 337240 120034
rect 337548 120006 337884 120034
rect 338192 120006 338528 120034
rect 333520 117360 333572 117366
rect 333520 117302 333572 117308
rect 333716 6186 333744 120006
rect 334624 117496 334676 117502
rect 334624 117438 334676 117444
rect 333888 117428 333940 117434
rect 333888 117370 333940 117376
rect 333796 117360 333848 117366
rect 333796 117302 333848 117308
rect 333704 6180 333756 6186
rect 333704 6122 333756 6128
rect 333808 4690 333836 117302
rect 333796 4684 333848 4690
rect 333796 4626 333848 4632
rect 333900 3806 333928 117370
rect 333888 3800 333940 3806
rect 333888 3742 333940 3748
rect 334636 3398 334664 117438
rect 334820 117434 334848 120006
rect 334808 117428 334860 117434
rect 334808 117370 334860 117376
rect 335280 5506 335308 120006
rect 336016 118454 336044 120006
rect 336004 118448 336056 118454
rect 336004 118390 336056 118396
rect 336660 117502 336688 120006
rect 336924 118244 336976 118250
rect 336924 118186 336976 118192
rect 336648 117496 336700 117502
rect 336648 117438 336700 117444
rect 335268 5500 335320 5506
rect 335268 5442 335320 5448
rect 334716 5160 334768 5166
rect 334716 5102 334768 5108
rect 334624 3392 334676 3398
rect 334624 3334 334676 3340
rect 332876 604 332928 610
rect 332876 546 332928 552
rect 333612 604 333664 610
rect 333612 546 333664 552
rect 333624 480 333652 546
rect 334728 480 334756 5102
rect 335912 3868 335964 3874
rect 335912 3810 335964 3816
rect 335924 480 335952 3810
rect 336936 2854 336964 118186
rect 337212 117366 337240 120006
rect 337856 118318 337884 120006
rect 338500 118386 338528 120006
rect 338730 119762 338758 120020
rect 338684 119734 338758 119762
rect 339374 119762 339402 120020
rect 340032 120006 340368 120034
rect 340584 120006 340828 120034
rect 341228 120006 341564 120034
rect 341872 120006 342208 120034
rect 342424 120006 342760 120034
rect 343068 120006 343496 120034
rect 343712 120006 344048 120034
rect 344264 120006 344600 120034
rect 339374 119734 339448 119762
rect 338488 118380 338540 118386
rect 338488 118322 338540 118328
rect 337844 118312 337896 118318
rect 337844 118254 337896 118260
rect 337384 117836 337436 117842
rect 337384 117778 337436 117784
rect 337200 117360 337252 117366
rect 337200 117302 337252 117308
rect 337396 3058 337424 117778
rect 338028 117360 338080 117366
rect 338028 117302 338080 117308
rect 338040 4758 338068 117302
rect 338684 115977 338712 119734
rect 339420 118250 339448 119734
rect 339408 118244 339460 118250
rect 339408 118186 339460 118192
rect 339684 118176 339736 118182
rect 339684 118118 339736 118124
rect 338764 117428 338816 117434
rect 338764 117370 338816 117376
rect 338670 115968 338726 115977
rect 338670 115903 338726 115912
rect 338304 5024 338356 5030
rect 338304 4966 338356 4972
rect 338028 4752 338080 4758
rect 338028 4694 338080 4700
rect 337384 3052 337436 3058
rect 337384 2994 337436 3000
rect 336924 2848 336976 2854
rect 336924 2790 336976 2796
rect 337016 2780 337068 2786
rect 337016 2722 337068 2728
rect 337028 610 337056 2722
rect 337016 604 337068 610
rect 337016 546 337068 552
rect 337108 604 337160 610
rect 337108 546 337160 552
rect 337120 480 337148 546
rect 338316 480 338344 4966
rect 338776 3942 338804 117370
rect 339038 115968 339094 115977
rect 339696 115938 339724 118118
rect 340340 117434 340368 120006
rect 340328 117428 340380 117434
rect 340328 117370 340380 117376
rect 339038 115903 339094 115912
rect 339684 115932 339736 115938
rect 339052 109018 339080 115903
rect 339684 115874 339736 115880
rect 339868 115932 339920 115938
rect 339868 115874 339920 115880
rect 339052 108990 339356 109018
rect 339328 96642 339356 108990
rect 339880 106350 339908 115874
rect 339684 106344 339736 106350
rect 339684 106286 339736 106292
rect 339868 106344 339920 106350
rect 339868 106286 339920 106292
rect 339328 96614 339448 96642
rect 339420 85626 339448 96614
rect 339236 85598 339448 85626
rect 339236 85542 339264 85598
rect 339132 85536 339184 85542
rect 339132 85478 339184 85484
rect 339224 85536 339276 85542
rect 339224 85478 339276 85484
rect 339144 84182 339172 85478
rect 338948 84176 339000 84182
rect 338948 84118 339000 84124
rect 339132 84176 339184 84182
rect 339132 84118 339184 84124
rect 338960 75290 338988 84118
rect 338960 75262 339172 75290
rect 339144 67810 339172 75262
rect 339144 67782 339356 67810
rect 339328 66366 339356 67782
rect 339224 66360 339276 66366
rect 339144 66308 339224 66314
rect 339144 66302 339276 66308
rect 339316 66360 339368 66366
rect 339316 66302 339368 66308
rect 339144 66286 339264 66302
rect 339144 64870 339172 66286
rect 339132 64864 339184 64870
rect 339132 64806 339184 64812
rect 339500 64864 339552 64870
rect 339500 64806 339552 64812
rect 339512 45626 339540 64806
rect 339224 45620 339276 45626
rect 339224 45562 339276 45568
rect 339500 45620 339552 45626
rect 339500 45562 339552 45568
rect 339236 37398 339264 45562
rect 339224 37392 339276 37398
rect 339224 37334 339276 37340
rect 339132 37256 339184 37262
rect 339132 37198 339184 37204
rect 339144 29050 339172 37198
rect 339052 29022 339172 29050
rect 339052 28778 339080 29022
rect 339052 28750 339264 28778
rect 339236 27554 339264 28750
rect 339236 27526 339356 27554
rect 339328 18018 339356 27526
rect 339316 18012 339368 18018
rect 339316 17954 339368 17960
rect 339408 18012 339460 18018
rect 339408 17954 339460 17960
rect 339420 9722 339448 17954
rect 339132 9716 339184 9722
rect 339132 9658 339184 9664
rect 339408 9716 339460 9722
rect 339408 9658 339460 9664
rect 339144 9586 339172 9658
rect 339132 9580 339184 9586
rect 339132 9522 339184 9528
rect 338764 3936 338816 3942
rect 338764 3878 338816 3884
rect 339500 3460 339552 3466
rect 339500 3402 339552 3408
rect 339512 480 339540 3402
rect 339696 2854 339724 106286
rect 340800 5370 340828 120006
rect 341156 117496 341208 117502
rect 341156 117438 341208 117444
rect 341168 116090 341196 117438
rect 341536 117366 341564 120006
rect 342180 118522 342208 120006
rect 342168 118516 342220 118522
rect 342168 118458 342220 118464
rect 342732 117366 342760 120006
rect 342904 117428 342956 117434
rect 342904 117370 342956 117376
rect 341524 117360 341576 117366
rect 341524 117302 341576 117308
rect 342168 117360 342220 117366
rect 342168 117302 342220 117308
rect 342720 117360 342772 117366
rect 342720 117302 342772 117308
rect 341168 116062 341242 116090
rect 341214 115954 341242 116062
rect 341214 115938 341288 115954
rect 341214 115932 341300 115938
rect 341214 115926 341248 115932
rect 341248 115874 341300 115880
rect 341432 115932 341484 115938
rect 341432 115874 341484 115880
rect 341260 115843 341288 115874
rect 341444 106282 341472 115874
rect 341432 106276 341484 106282
rect 341432 106218 341484 106224
rect 341524 106276 341576 106282
rect 341524 106218 341576 106224
rect 341536 96694 341564 106218
rect 341524 96688 341576 96694
rect 341524 96630 341576 96636
rect 341432 96620 341484 96626
rect 341432 96562 341484 96568
rect 341444 95266 341472 96562
rect 341432 95260 341484 95266
rect 341432 95202 341484 95208
rect 341524 95260 341576 95266
rect 341524 95202 341576 95208
rect 341536 89758 341564 95202
rect 341340 89752 341392 89758
rect 341524 89752 341576 89758
rect 341392 89700 341524 89706
rect 341340 89694 341576 89700
rect 341352 89678 341564 89694
rect 341536 80730 341564 89678
rect 341536 80702 341748 80730
rect 341720 75954 341748 80702
rect 341708 75948 341760 75954
rect 341708 75890 341760 75896
rect 341892 75948 341944 75954
rect 341892 75890 341944 75896
rect 341904 67658 341932 75890
rect 341524 67652 341576 67658
rect 341524 67594 341576 67600
rect 341892 67652 341944 67658
rect 341892 67594 341944 67600
rect 341536 60738 341564 67594
rect 341352 60710 341564 60738
rect 341352 46986 341380 60710
rect 341248 46980 341300 46986
rect 341248 46922 341300 46928
rect 341340 46980 341392 46986
rect 341340 46922 341392 46928
rect 341260 46850 341288 46922
rect 341248 46844 341300 46850
rect 341248 46786 341300 46792
rect 341432 46844 341484 46850
rect 341432 46786 341484 46792
rect 341444 22114 341472 46786
rect 341444 22098 341564 22114
rect 341444 22092 341576 22098
rect 341444 22086 341524 22092
rect 341524 22034 341576 22040
rect 341708 22092 341760 22098
rect 341708 22034 341760 22040
rect 341720 12050 341748 22034
rect 341720 12022 341840 12050
rect 341812 11778 341840 12022
rect 341720 11750 341840 11778
rect 340788 5364 340840 5370
rect 340788 5306 340840 5312
rect 341720 3874 341748 11750
rect 342180 8022 342208 117302
rect 342168 8016 342220 8022
rect 342168 7958 342220 7964
rect 341892 4956 341944 4962
rect 341892 4898 341944 4904
rect 341708 3868 341760 3874
rect 341708 3810 341760 3816
rect 339684 2848 339736 2854
rect 339684 2790 339736 2796
rect 340144 2780 340196 2786
rect 340144 2722 340196 2728
rect 340156 610 340184 2722
rect 340144 604 340196 610
rect 340144 546 340196 552
rect 340696 604 340748 610
rect 340696 546 340748 552
rect 340708 480 340736 546
rect 341904 480 341932 4898
rect 342916 3738 342944 117370
rect 343088 9580 343140 9586
rect 343088 9522 343140 9528
rect 343100 5438 343128 9522
rect 343468 7954 343496 120006
rect 343916 118108 343968 118114
rect 343916 118050 343968 118056
rect 343548 117360 343600 117366
rect 343548 117302 343600 117308
rect 343456 7948 343508 7954
rect 343456 7890 343508 7896
rect 343088 5432 343140 5438
rect 343088 5374 343140 5380
rect 343560 5302 343588 117302
rect 343928 115938 343956 118050
rect 344020 117434 344048 120006
rect 344008 117428 344060 117434
rect 344008 117370 344060 117376
rect 344572 117366 344600 120006
rect 344894 119762 344922 120020
rect 345552 120006 345888 120034
rect 346104 120006 346348 120034
rect 346748 120006 347084 120034
rect 347300 120006 347636 120034
rect 347944 120006 348280 120034
rect 348588 120006 349016 120034
rect 349140 120006 349476 120034
rect 349784 120006 350120 120034
rect 344848 119734 344922 119762
rect 344560 117360 344612 117366
rect 344560 117302 344612 117308
rect 343916 115932 343968 115938
rect 343916 115874 343968 115880
rect 344100 115932 344152 115938
rect 344100 115874 344152 115880
rect 344112 106350 344140 115874
rect 343916 106344 343968 106350
rect 343916 106286 343968 106292
rect 344100 106344 344152 106350
rect 344100 106286 344152 106292
rect 343928 96626 343956 106286
rect 343916 96620 343968 96626
rect 343916 96562 343968 96568
rect 344100 96620 344152 96626
rect 344100 96562 344152 96568
rect 344112 87038 344140 96562
rect 343916 87032 343968 87038
rect 343916 86974 343968 86980
rect 344100 87032 344152 87038
rect 344100 86974 344152 86980
rect 343548 5296 343600 5302
rect 343548 5238 343600 5244
rect 342904 3732 342956 3738
rect 342904 3674 342956 3680
rect 343088 3528 343140 3534
rect 343088 3470 343140 3476
rect 343100 480 343128 3470
rect 343928 2854 343956 86974
rect 344848 7886 344876 119734
rect 345860 117910 345888 120006
rect 345848 117904 345900 117910
rect 345848 117846 345900 117852
rect 345664 117428 345716 117434
rect 345664 117370 345716 117376
rect 344928 117360 344980 117366
rect 344928 117302 344980 117308
rect 344836 7880 344888 7886
rect 344836 7822 344888 7828
rect 344940 5234 344968 117302
rect 344928 5228 344980 5234
rect 344928 5170 344980 5176
rect 345480 4888 345532 4894
rect 345480 4830 345532 4836
rect 343916 2848 343968 2854
rect 343916 2790 343968 2796
rect 344008 2780 344060 2786
rect 344008 2722 344060 2728
rect 344020 610 344048 2722
rect 344008 604 344060 610
rect 344008 546 344060 552
rect 344284 604 344336 610
rect 344284 546 344336 552
rect 344296 480 344324 546
rect 345492 480 345520 4830
rect 345676 3670 345704 117370
rect 346320 5166 346348 120006
rect 347056 117366 347084 120006
rect 347608 117434 347636 120006
rect 347964 118040 348016 118046
rect 347964 117982 348016 117988
rect 347596 117428 347648 117434
rect 347596 117370 347648 117376
rect 347044 117360 347096 117366
rect 347044 117302 347096 117308
rect 347688 117360 347740 117366
rect 347688 117302 347740 117308
rect 347700 7818 347728 117302
rect 347688 7812 347740 7818
rect 347688 7754 347740 7760
rect 346308 5160 346360 5166
rect 346308 5102 346360 5108
rect 345664 3664 345716 3670
rect 345664 3606 345716 3612
rect 346676 3256 346728 3262
rect 346676 3198 346728 3204
rect 346688 480 346716 3198
rect 347976 626 348004 117982
rect 348252 117366 348280 120006
rect 348424 118448 348476 118454
rect 348424 118390 348476 118396
rect 348240 117360 348292 117366
rect 348240 117302 348292 117308
rect 348436 5778 348464 118390
rect 348988 7750 349016 120006
rect 349448 118658 349476 120006
rect 349436 118652 349488 118658
rect 349436 118594 349488 118600
rect 349804 117428 349856 117434
rect 349804 117370 349856 117376
rect 349068 117360 349120 117366
rect 349068 117302 349120 117308
rect 348976 7744 349028 7750
rect 348976 7686 349028 7692
rect 348424 5772 348476 5778
rect 348424 5714 348476 5720
rect 349080 5098 349108 117302
rect 349068 5092 349120 5098
rect 349068 5034 349120 5040
rect 349068 4820 349120 4826
rect 349068 4762 349120 4768
rect 347884 598 348004 626
rect 347884 480 347912 598
rect 349080 480 349108 4762
rect 349816 3534 349844 117370
rect 350092 117366 350120 120006
rect 350414 119762 350442 120020
rect 350980 120006 351316 120034
rect 351624 120006 351868 120034
rect 352268 120006 352604 120034
rect 352820 120006 353156 120034
rect 353464 120006 353800 120034
rect 354108 120006 354536 120034
rect 354660 120006 354996 120034
rect 355304 120006 355640 120034
rect 350368 119734 350442 119762
rect 350080 117360 350132 117366
rect 350080 117302 350132 117308
rect 350368 7682 350396 119734
rect 351184 118312 351236 118318
rect 351184 118254 351236 118260
rect 350448 117360 350500 117366
rect 350448 117302 350500 117308
rect 350356 7676 350408 7682
rect 350356 7618 350408 7624
rect 350460 5030 350488 117302
rect 351196 6594 351224 118254
rect 351288 117366 351316 120006
rect 351276 117360 351328 117366
rect 351276 117302 351328 117308
rect 351092 6588 351144 6594
rect 351092 6530 351144 6536
rect 351184 6588 351236 6594
rect 351184 6530 351236 6536
rect 351104 6474 351132 6530
rect 351104 6446 351408 6474
rect 350448 5024 350500 5030
rect 350448 4966 350500 4972
rect 349804 3528 349856 3534
rect 349804 3470 349856 3476
rect 350264 3188 350316 3194
rect 350264 3130 350316 3136
rect 350276 480 350304 3130
rect 351380 480 351408 6446
rect 351840 4962 351868 120006
rect 352576 117366 352604 120006
rect 353128 117638 353156 120006
rect 353116 117632 353168 117638
rect 353116 117574 353168 117580
rect 353772 117366 353800 120006
rect 353944 118244 353996 118250
rect 353944 118186 353996 118192
rect 352472 117360 352524 117366
rect 352472 117302 352524 117308
rect 352564 117360 352616 117366
rect 352564 117302 352616 117308
rect 353208 117360 353260 117366
rect 353208 117302 353260 117308
rect 353760 117360 353812 117366
rect 353760 117302 353812 117308
rect 352484 117178 352512 117302
rect 352484 117150 352604 117178
rect 352576 5930 352604 117150
rect 353220 7614 353248 117302
rect 353208 7608 353260 7614
rect 353208 7550 353260 7556
rect 352484 5902 352604 5930
rect 351828 4956 351880 4962
rect 351828 4898 351880 4904
rect 352484 3466 352512 5902
rect 352564 5840 352616 5846
rect 352564 5782 352616 5788
rect 352472 3460 352524 3466
rect 352472 3402 352524 3408
rect 352576 480 352604 5782
rect 353956 5574 353984 118186
rect 354508 9042 354536 120006
rect 354968 118114 354996 120006
rect 354956 118108 355008 118114
rect 354956 118050 355008 118056
rect 355612 117366 355640 120006
rect 355934 119762 355962 120020
rect 356500 120006 356836 120034
rect 357144 120006 357388 120034
rect 357788 120006 358124 120034
rect 358340 120006 358768 120034
rect 358984 120006 359320 120034
rect 359628 120006 360056 120034
rect 360180 120006 360516 120034
rect 360824 120006 361160 120034
rect 355888 119734 355962 119762
rect 354588 117360 354640 117366
rect 354588 117302 354640 117308
rect 355600 117360 355652 117366
rect 355600 117302 355652 117308
rect 354496 9036 354548 9042
rect 354496 8978 354548 8984
rect 354496 6724 354548 6730
rect 354496 6666 354548 6672
rect 354508 5778 354536 6666
rect 354496 5772 354548 5778
rect 354496 5714 354548 5720
rect 353944 5568 353996 5574
rect 353944 5510 353996 5516
rect 354600 4894 354628 117302
rect 355888 8974 355916 119734
rect 356808 118250 356836 120006
rect 356796 118244 356848 118250
rect 356796 118186 356848 118192
rect 355968 117360 356020 117366
rect 355968 117302 356020 117308
rect 355876 8968 355928 8974
rect 355876 8910 355928 8916
rect 354956 5908 355008 5914
rect 354956 5850 355008 5856
rect 354588 4888 354640 4894
rect 354588 4830 354640 4836
rect 353760 3120 353812 3126
rect 353760 3062 353812 3068
rect 353772 480 353800 3062
rect 354968 480 354996 5850
rect 355980 4826 356008 117302
rect 357360 7342 357388 120006
rect 357992 117768 358044 117774
rect 357992 117710 358044 117716
rect 358004 117178 358032 117710
rect 358096 117366 358124 120006
rect 358084 117360 358136 117366
rect 358084 117302 358136 117308
rect 358636 117360 358688 117366
rect 358636 117302 358688 117308
rect 358004 117150 358124 117178
rect 357348 7336 357400 7342
rect 357348 7278 357400 7284
rect 356152 6044 356204 6050
rect 356152 5986 356204 5992
rect 355968 4820 356020 4826
rect 355968 4762 356020 4768
rect 356164 480 356192 5986
rect 358096 3602 358124 117150
rect 358648 9994 358676 117302
rect 358636 9988 358688 9994
rect 358636 9930 358688 9936
rect 358740 7274 358768 120006
rect 359292 118182 359320 120006
rect 359280 118176 359332 118182
rect 359280 118118 359332 118124
rect 360028 10062 360056 120006
rect 360108 118176 360160 118182
rect 360108 118118 360160 118124
rect 360016 10056 360068 10062
rect 360016 9998 360068 10004
rect 360120 8634 360148 118118
rect 360488 117706 360516 120006
rect 360476 117700 360528 117706
rect 360476 117642 360528 117648
rect 361132 117366 361160 120006
rect 361454 119762 361482 120020
rect 362020 120006 362356 120034
rect 362664 120006 362908 120034
rect 363308 120006 363644 120034
rect 363860 120006 364104 120034
rect 364504 120006 364840 120034
rect 365056 120006 365576 120034
rect 365700 120006 366036 120034
rect 366344 120006 366680 120034
rect 361408 119734 361482 119762
rect 361120 117360 361172 117366
rect 361120 117302 361172 117308
rect 361408 10198 361436 119734
rect 362328 118318 362356 120006
rect 362316 118312 362368 118318
rect 362316 118254 362368 118260
rect 361488 117360 361540 117366
rect 361488 117302 361540 117308
rect 361396 10192 361448 10198
rect 361396 10134 361448 10140
rect 361500 8702 361528 117302
rect 362880 8770 362908 120006
rect 363616 117366 363644 120006
rect 364076 118590 364104 120006
rect 364064 118584 364116 118590
rect 364064 118526 364116 118532
rect 364812 117366 364840 120006
rect 364984 118108 365036 118114
rect 364984 118050 365036 118056
rect 363604 117360 363656 117366
rect 363604 117302 363656 117308
rect 364248 117360 364300 117366
rect 364248 117302 364300 117308
rect 364800 117360 364852 117366
rect 364800 117302 364852 117308
rect 364260 10130 364288 117302
rect 364248 10124 364300 10130
rect 364248 10066 364300 10072
rect 362868 8764 362920 8770
rect 362868 8706 362920 8712
rect 361488 8696 361540 8702
rect 361488 8638 361540 8644
rect 360108 8628 360160 8634
rect 360108 8570 360160 8576
rect 358728 7268 358780 7274
rect 358728 7210 358780 7216
rect 360200 6928 360252 6934
rect 360200 6870 360252 6876
rect 360212 6730 360240 6870
rect 362132 6860 362184 6866
rect 362132 6802 362184 6808
rect 360200 6724 360252 6730
rect 360200 6666 360252 6672
rect 358544 6112 358596 6118
rect 358544 6054 358596 6060
rect 357348 3596 357400 3602
rect 357348 3538 357400 3544
rect 358084 3596 358136 3602
rect 358084 3538 358136 3544
rect 357360 480 357388 3538
rect 358556 480 358584 6054
rect 359740 5976 359792 5982
rect 359740 5918 359792 5924
rect 359752 480 359780 5918
rect 360936 3324 360988 3330
rect 360936 3266 360988 3272
rect 360948 480 360976 3266
rect 362144 480 362172 6802
rect 363328 6792 363380 6798
rect 363328 6734 363380 6740
rect 363340 480 363368 6734
rect 364996 3602 365024 118050
rect 365548 10266 365576 120006
rect 366008 118250 366036 120006
rect 365996 118244 366048 118250
rect 365996 118186 366048 118192
rect 366652 117366 366680 120006
rect 366882 119762 366910 120020
rect 367540 120006 367876 120034
rect 368184 120006 368428 120034
rect 368736 120006 369072 120034
rect 369380 120006 369716 120034
rect 370024 120006 370360 120034
rect 370576 120006 371096 120034
rect 371220 120006 371556 120034
rect 371864 120006 372200 120034
rect 366882 119734 366956 119762
rect 365628 117360 365680 117366
rect 365628 117302 365680 117308
rect 366640 117360 366692 117366
rect 366640 117302 366692 117308
rect 365536 10260 365588 10266
rect 365536 10202 365588 10208
rect 365640 8838 365668 117302
rect 366928 11014 366956 119734
rect 367848 117434 367876 120006
rect 367836 117428 367888 117434
rect 367836 117370 367888 117376
rect 367008 117360 367060 117366
rect 367008 117302 367060 117308
rect 366916 11008 366968 11014
rect 366916 10950 366968 10956
rect 367020 8906 367048 117302
rect 368400 9654 368428 120006
rect 369044 117366 369072 120006
rect 369688 118454 369716 120006
rect 369676 118448 369728 118454
rect 369676 118390 369728 118396
rect 369124 117428 369176 117434
rect 369124 117370 369176 117376
rect 369032 117360 369084 117366
rect 369032 117302 369084 117308
rect 368388 9648 368440 9654
rect 368388 9590 368440 9596
rect 367008 8900 367060 8906
rect 367008 8842 367060 8848
rect 365628 8832 365680 8838
rect 365628 8774 365680 8780
rect 366916 6656 366968 6662
rect 366916 6598 366968 6604
rect 365720 4276 365772 4282
rect 365720 4218 365772 4224
rect 364524 3596 364576 3602
rect 364524 3538 364576 3544
rect 364984 3596 365036 3602
rect 364984 3538 365036 3544
rect 364536 480 364564 3538
rect 365732 480 365760 4218
rect 366928 480 366956 6598
rect 368020 4140 368072 4146
rect 368020 4082 368072 4088
rect 368032 480 368060 4082
rect 369136 3330 369164 117370
rect 370332 117366 370360 120006
rect 369768 117360 369820 117366
rect 369768 117302 369820 117308
rect 370320 117360 370372 117366
rect 370320 117302 370372 117308
rect 369780 10946 369808 117302
rect 369768 10940 369820 10946
rect 369768 10882 369820 10888
rect 371068 10878 371096 120006
rect 371528 117434 371556 120006
rect 371516 117428 371568 117434
rect 371516 117370 371568 117376
rect 372172 117366 372200 120006
rect 372402 119762 372430 120020
rect 373060 120006 373396 120034
rect 373704 120006 373948 120034
rect 374256 120006 374592 120034
rect 374900 120006 375328 120034
rect 375544 120006 375880 120034
rect 376096 120006 376616 120034
rect 376740 120006 377076 120034
rect 377384 120006 377720 120034
rect 372402 119734 372476 119762
rect 371148 117360 371200 117366
rect 371148 117302 371200 117308
rect 372160 117360 372212 117366
rect 372160 117302 372212 117308
rect 371056 10872 371108 10878
rect 371056 10814 371108 10820
rect 371160 9586 371188 117302
rect 372448 10810 372476 119734
rect 373368 118114 373396 120006
rect 373356 118108 373408 118114
rect 373356 118050 373408 118056
rect 372528 117360 372580 117366
rect 372528 117302 372580 117308
rect 372436 10804 372488 10810
rect 372436 10746 372488 10752
rect 371148 9580 371200 9586
rect 371148 9522 371200 9528
rect 372540 9518 372568 117302
rect 372528 9512 372580 9518
rect 372528 9454 372580 9460
rect 370412 6520 370464 6526
rect 370412 6462 370464 6468
rect 369216 4344 369268 4350
rect 369216 4286 369268 4292
rect 369124 3324 369176 3330
rect 369124 3266 369176 3272
rect 369228 480 369256 4286
rect 370424 480 370452 6462
rect 373920 5710 373948 120006
rect 374564 117366 374592 120006
rect 374644 118448 374696 118454
rect 374644 118390 374696 118396
rect 374656 118182 374684 118390
rect 374644 118176 374696 118182
rect 374644 118118 374696 118124
rect 374644 118040 374696 118046
rect 374644 117982 374696 117988
rect 374552 117360 374604 117366
rect 374552 117302 374604 117308
rect 374000 6452 374052 6458
rect 374000 6394 374052 6400
rect 373908 5704 373960 5710
rect 373908 5646 373960 5652
rect 372804 4412 372856 4418
rect 372804 4354 372856 4360
rect 371608 4072 371660 4078
rect 371608 4014 371660 4020
rect 371620 480 371648 4014
rect 372816 480 372844 4354
rect 374012 480 374040 6394
rect 374656 3126 374684 117982
rect 375196 117360 375248 117366
rect 375196 117302 375248 117308
rect 375208 10742 375236 117302
rect 375196 10736 375248 10742
rect 375196 10678 375248 10684
rect 375300 3398 375328 120006
rect 375852 117366 375880 120006
rect 375840 117360 375892 117366
rect 375840 117302 375892 117308
rect 376588 10674 376616 120006
rect 377048 118046 377076 120006
rect 377036 118040 377088 118046
rect 377036 117982 377088 117988
rect 377404 117428 377456 117434
rect 377404 117370 377456 117376
rect 376668 117360 376720 117366
rect 376668 117302 376720 117308
rect 376576 10668 376628 10674
rect 376576 10610 376628 10616
rect 376680 7546 376708 117302
rect 376392 7540 376444 7546
rect 376392 7482 376444 7488
rect 376668 7540 376720 7546
rect 376668 7482 376720 7488
rect 376404 5642 376432 7482
rect 376760 6928 376812 6934
rect 376758 6896 376760 6905
rect 376812 6896 376814 6905
rect 376758 6831 376814 6840
rect 376392 5636 376444 5642
rect 376392 5578 376444 5584
rect 376392 4480 376444 4486
rect 376392 4422 376444 4428
rect 375196 3392 375248 3398
rect 375196 3334 375248 3340
rect 375288 3392 375340 3398
rect 375288 3334 375340 3340
rect 374644 3120 374696 3126
rect 374644 3062 374696 3068
rect 375208 480 375236 3334
rect 376404 480 376432 4422
rect 377416 3262 377444 117370
rect 377692 117366 377720 120006
rect 377922 119762 377950 120020
rect 378580 120006 378916 120034
rect 379224 120006 379376 120034
rect 379776 120006 380112 120034
rect 380420 120006 380756 120034
rect 381064 120006 381400 120034
rect 381616 120006 382136 120034
rect 382260 120006 382596 120034
rect 382812 120006 382964 120034
rect 377922 119734 377996 119762
rect 377680 117360 377732 117366
rect 377680 117302 377732 117308
rect 377968 10606 377996 119734
rect 378888 117366 378916 120006
rect 378048 117360 378100 117366
rect 378048 117302 378100 117308
rect 378876 117360 378928 117366
rect 378876 117302 378928 117308
rect 377956 10600 378008 10606
rect 377956 10542 378008 10548
rect 377588 6384 377640 6390
rect 377588 6326 377640 6332
rect 377404 3256 377456 3262
rect 377404 3198 377456 3204
rect 377600 480 377628 6326
rect 378060 5778 378088 117302
rect 379348 5914 379376 120006
rect 380084 117366 380112 120006
rect 380164 118584 380216 118590
rect 380164 118526 380216 118532
rect 379428 117360 379480 117366
rect 379428 117302 379480 117308
rect 380072 117360 380124 117366
rect 380072 117302 380124 117308
rect 379336 5908 379388 5914
rect 379336 5850 379388 5856
rect 378048 5772 378100 5778
rect 378048 5714 378100 5720
rect 379440 4146 379468 117302
rect 379610 6896 379666 6905
rect 379610 6831 379666 6840
rect 379624 6798 379652 6831
rect 379612 6792 379664 6798
rect 379612 6734 379664 6740
rect 379980 4616 380032 4622
rect 379980 4558 380032 4564
rect 379428 4140 379480 4146
rect 379428 4082 379480 4088
rect 378784 4004 378836 4010
rect 378784 3946 378836 3952
rect 378796 480 378824 3946
rect 379992 480 380020 4558
rect 380176 3194 380204 118526
rect 380728 117978 380756 120006
rect 380716 117972 380768 117978
rect 380716 117914 380768 117920
rect 380256 117700 380308 117706
rect 380256 117642 380308 117648
rect 380268 117502 380296 117642
rect 380256 117496 380308 117502
rect 380256 117438 380308 117444
rect 381372 117366 381400 120006
rect 380808 117360 380860 117366
rect 380808 117302 380860 117308
rect 381360 117360 381412 117366
rect 381360 117302 381412 117308
rect 380820 10538 380848 117302
rect 380808 10532 380860 10538
rect 380808 10474 380860 10480
rect 382108 10470 382136 120006
rect 382568 117366 382596 120006
rect 382188 117360 382240 117366
rect 382188 117302 382240 117308
rect 382556 117360 382608 117366
rect 382556 117302 382608 117308
rect 382096 10464 382148 10470
rect 382096 10406 382148 10412
rect 381176 6316 381228 6322
rect 381176 6258 381228 6264
rect 380164 3188 380216 3194
rect 380164 3130 380216 3136
rect 381188 480 381216 6258
rect 382200 5846 382228 117302
rect 382936 114578 382964 120006
rect 383442 119762 383470 120020
rect 384100 120006 384436 120034
rect 384652 120006 384804 120034
rect 385296 120006 385632 120034
rect 385940 120006 386276 120034
rect 386492 120006 386828 120034
rect 387136 120006 387656 120034
rect 387780 120006 388116 120034
rect 388332 120006 388852 120034
rect 388976 120006 389128 120034
rect 389620 120006 389956 120034
rect 390172 120006 390508 120034
rect 390816 120006 391152 120034
rect 391460 120006 391796 120034
rect 392012 120006 392348 120034
rect 392656 120006 393176 120034
rect 393300 120006 393636 120034
rect 393852 120006 394372 120034
rect 394496 120006 394648 120034
rect 395140 120006 395476 120034
rect 395692 120006 396028 120034
rect 396336 120006 396672 120034
rect 396980 120006 397316 120034
rect 397532 120006 397868 120034
rect 398176 120006 398696 120034
rect 398820 120006 399156 120034
rect 399372 120006 399708 120034
rect 383442 119734 383516 119762
rect 382924 114572 382976 114578
rect 382924 114514 382976 114520
rect 383108 114572 383160 114578
rect 383108 114514 383160 114520
rect 383120 109138 383148 114514
rect 383108 109132 383160 109138
rect 383108 109074 383160 109080
rect 383108 108996 383160 109002
rect 383108 108938 383160 108944
rect 383120 106321 383148 108938
rect 383106 106312 383162 106321
rect 383106 106247 383162 106256
rect 383290 106312 383346 106321
rect 383290 106247 383346 106256
rect 383304 99482 383332 106247
rect 383292 99476 383344 99482
rect 383292 99418 383344 99424
rect 383200 99340 383252 99346
rect 383200 99282 383252 99288
rect 383212 96626 383240 99282
rect 382924 96620 382976 96626
rect 382924 96562 382976 96568
rect 383200 96620 383252 96626
rect 383200 96562 383252 96568
rect 382936 87038 382964 96562
rect 382924 87032 382976 87038
rect 382924 86974 382976 86980
rect 383108 87032 383160 87038
rect 383108 86974 383160 86980
rect 383120 79914 383148 86974
rect 383120 79886 383240 79914
rect 383212 77217 383240 79886
rect 383198 77208 383254 77217
rect 383198 77143 383254 77152
rect 383292 67652 383344 67658
rect 383292 67594 383344 67600
rect 383304 60858 383332 67594
rect 383292 60852 383344 60858
rect 383292 60794 383344 60800
rect 383200 60716 383252 60722
rect 383200 60658 383252 60664
rect 383212 57934 383240 60658
rect 383016 57928 383068 57934
rect 383016 57870 383068 57876
rect 383200 57928 383252 57934
rect 383200 57870 383252 57876
rect 383028 48346 383056 57870
rect 383016 48340 383068 48346
rect 383016 48282 383068 48288
rect 383292 48340 383344 48346
rect 383292 48282 383344 48288
rect 383304 43466 383332 48282
rect 383212 43438 383332 43466
rect 383212 38622 383240 43438
rect 383016 38616 383068 38622
rect 383016 38558 383068 38564
rect 383200 38616 383252 38622
rect 383200 38558 383252 38564
rect 383028 29034 383056 38558
rect 383016 29028 383068 29034
rect 383016 28970 383068 28976
rect 383292 29028 383344 29034
rect 383292 28970 383344 28976
rect 383304 28937 383332 28970
rect 383290 28928 383346 28937
rect 383290 28863 383346 28872
rect 383382 21992 383438 22001
rect 383382 21927 383438 21936
rect 383396 7410 383424 21927
rect 383384 7404 383436 7410
rect 383384 7346 383436 7352
rect 383488 6050 383516 119734
rect 383660 117496 383712 117502
rect 383658 117464 383660 117473
rect 383712 117464 383714 117473
rect 383658 117399 383714 117408
rect 384408 117366 384436 120006
rect 384776 117450 384804 120006
rect 384776 117422 384988 117450
rect 383568 117360 383620 117366
rect 383568 117302 383620 117308
rect 384396 117360 384448 117366
rect 384396 117302 384448 117308
rect 384856 117360 384908 117366
rect 384856 117302 384908 117308
rect 383476 6044 383528 6050
rect 383476 5986 383528 5992
rect 383580 5930 383608 117302
rect 383658 77208 383714 77217
rect 383658 77143 383714 77152
rect 383672 67658 383700 77143
rect 383660 67652 383712 67658
rect 383660 67594 383712 67600
rect 384868 10402 384896 117302
rect 384856 10396 384908 10402
rect 384856 10338 384908 10344
rect 384960 7478 384988 117422
rect 385604 117366 385632 120006
rect 385592 117360 385644 117366
rect 385592 117302 385644 117308
rect 386248 12238 386276 120006
rect 386800 117366 386828 120006
rect 387628 117450 387656 120006
rect 387628 117422 387748 117450
rect 386328 117360 386380 117366
rect 386328 117302 386380 117308
rect 386788 117360 386840 117366
rect 386788 117302 386840 117308
rect 387616 117360 387668 117366
rect 387616 117302 387668 117308
rect 386236 12232 386288 12238
rect 386236 12174 386288 12180
rect 384948 7472 385000 7478
rect 384948 7414 385000 7420
rect 384672 6248 384724 6254
rect 384672 6190 384724 6196
rect 383488 5902 383608 5930
rect 382188 5840 382240 5846
rect 382188 5782 382240 5788
rect 383488 4078 383516 5902
rect 383568 4548 383620 4554
rect 383568 4490 383620 4496
rect 383476 4072 383528 4078
rect 383476 4014 383528 4020
rect 382372 3052 382424 3058
rect 382372 2994 382424 3000
rect 382384 480 382412 2994
rect 383580 480 383608 4490
rect 384684 480 384712 6190
rect 386340 5982 386368 117302
rect 387628 7546 387656 117302
rect 387616 7540 387668 7546
rect 387616 7482 387668 7488
rect 387248 6792 387300 6798
rect 387248 6734 387300 6740
rect 387260 6526 387288 6734
rect 387248 6520 387300 6526
rect 387248 6462 387300 6468
rect 387720 6118 387748 117422
rect 388088 117366 388116 120006
rect 388076 117360 388128 117366
rect 388076 117302 388128 117308
rect 388824 109070 388852 120006
rect 388904 117360 388956 117366
rect 388904 117302 388956 117308
rect 388812 109064 388864 109070
rect 388812 109006 388864 109012
rect 388916 12170 388944 117302
rect 388996 109064 389048 109070
rect 388996 109006 389048 109012
rect 388904 12164 388956 12170
rect 388904 12106 388956 12112
rect 389008 8294 389036 109006
rect 388996 8288 389048 8294
rect 388996 8230 389048 8236
rect 389100 6866 389128 120006
rect 389928 117366 389956 120006
rect 389916 117360 389968 117366
rect 389916 117302 389968 117308
rect 390376 117360 390428 117366
rect 390376 117302 390428 117308
rect 390388 12102 390416 117302
rect 390376 12096 390428 12102
rect 390376 12038 390428 12044
rect 390480 8226 390508 120006
rect 391124 117366 391152 120006
rect 391112 117360 391164 117366
rect 391112 117302 391164 117308
rect 391768 12034 391796 120006
rect 392320 117366 392348 120006
rect 393148 117450 393176 120006
rect 393228 117700 393280 117706
rect 393228 117642 393280 117648
rect 393240 117609 393268 117642
rect 393226 117600 393282 117609
rect 393226 117535 393282 117544
rect 393148 117422 393268 117450
rect 391848 117360 391900 117366
rect 391848 117302 391900 117308
rect 392308 117360 392360 117366
rect 392308 117302 392360 117308
rect 393136 117360 393188 117366
rect 393136 117302 393188 117308
rect 391756 12028 391808 12034
rect 391756 11970 391808 11976
rect 391860 10282 391888 117302
rect 391768 10254 391888 10282
rect 390468 8220 390520 8226
rect 390468 8162 390520 8168
rect 389088 6860 389140 6866
rect 389088 6802 389140 6808
rect 391768 6730 391796 10254
rect 393148 9450 393176 117302
rect 393136 9444 393188 9450
rect 393136 9386 393188 9392
rect 393240 6730 393268 117422
rect 393608 117366 393636 120006
rect 393596 117360 393648 117366
rect 393596 117302 393648 117308
rect 394344 109070 394372 120006
rect 394424 117360 394476 117366
rect 394424 117302 394476 117308
rect 394332 109064 394384 109070
rect 394332 109006 394384 109012
rect 394436 11966 394464 117302
rect 394516 109064 394568 109070
rect 394516 109006 394568 109012
rect 394424 11960 394476 11966
rect 394424 11902 394476 11908
rect 394528 9382 394556 109006
rect 394516 9376 394568 9382
rect 394516 9318 394568 9324
rect 391756 6724 391808 6730
rect 391756 6666 391808 6672
rect 393228 6724 393280 6730
rect 393228 6666 393280 6672
rect 394620 6662 394648 120006
rect 394700 117768 394752 117774
rect 394884 117768 394936 117774
rect 394752 117716 394884 117722
rect 394700 117710 394936 117716
rect 394712 117694 394924 117710
rect 395448 117366 395476 120006
rect 395436 117360 395488 117366
rect 395436 117302 395488 117308
rect 395896 117360 395948 117366
rect 395896 117302 395948 117308
rect 395908 11898 395936 117302
rect 395896 11892 395948 11898
rect 395896 11834 395948 11840
rect 396000 9314 396028 120006
rect 396264 118380 396316 118386
rect 396264 118322 396316 118328
rect 395988 9308 396040 9314
rect 395988 9250 396040 9256
rect 394608 6656 394660 6662
rect 394608 6598 394660 6604
rect 395436 6588 395488 6594
rect 395436 6530 395488 6536
rect 391848 6520 391900 6526
rect 391848 6462 391900 6468
rect 388260 6180 388312 6186
rect 388260 6122 388312 6128
rect 387708 6112 387760 6118
rect 387708 6054 387760 6060
rect 386328 5976 386380 5982
rect 386328 5918 386380 5924
rect 387064 4684 387116 4690
rect 387064 4626 387116 4632
rect 385868 3800 385920 3806
rect 385868 3742 385920 3748
rect 385880 480 385908 3742
rect 387076 480 387104 4626
rect 388272 480 388300 6122
rect 390652 5500 390704 5506
rect 390652 5442 390704 5448
rect 389456 3936 389508 3942
rect 389456 3878 389508 3884
rect 389468 480 389496 3878
rect 390664 480 390692 5442
rect 391860 480 391888 6462
rect 394240 4752 394292 4758
rect 394240 4694 394292 4700
rect 393044 3868 393096 3874
rect 393044 3810 393096 3816
rect 393056 480 393084 3810
rect 394252 480 394280 4694
rect 395448 480 395476 6530
rect 396276 626 396304 118322
rect 396644 117366 396672 120006
rect 396632 117360 396684 117366
rect 396632 117302 396684 117308
rect 397288 11830 397316 120006
rect 397840 117366 397868 120006
rect 398668 117450 398696 120006
rect 398668 117422 398788 117450
rect 397368 117360 397420 117366
rect 397368 117302 397420 117308
rect 397828 117360 397880 117366
rect 397828 117302 397880 117308
rect 398656 117360 398708 117366
rect 398656 117302 398708 117308
rect 397276 11824 397328 11830
rect 397276 11766 397328 11772
rect 397380 6594 397408 117302
rect 398668 9246 398696 117302
rect 398656 9240 398708 9246
rect 398656 9182 398708 9188
rect 397368 6588 397420 6594
rect 397368 6530 397420 6536
rect 398760 6526 398788 117422
rect 399128 117366 399156 120006
rect 399680 117434 399708 120006
rect 400002 119762 400030 120020
rect 400568 120006 400904 120034
rect 401212 120006 401548 120034
rect 401856 120006 402192 120034
rect 402408 120006 402928 120034
rect 403052 120006 403388 120034
rect 400002 119734 400076 119762
rect 399668 117428 399720 117434
rect 399668 117370 399720 117376
rect 399116 117360 399168 117366
rect 399116 117302 399168 117308
rect 399944 117360 399996 117366
rect 399944 117302 399996 117308
rect 399956 11762 399984 117302
rect 399944 11756 399996 11762
rect 399944 11698 399996 11704
rect 398748 6520 398800 6526
rect 398748 6462 398800 6468
rect 400048 6458 400076 119734
rect 400876 118386 400904 120006
rect 400956 118516 401008 118522
rect 400956 118458 401008 118464
rect 400864 118380 400916 118386
rect 400864 118322 400916 118328
rect 400128 117428 400180 117434
rect 400128 117370 400180 117376
rect 400036 6452 400088 6458
rect 400036 6394 400088 6400
rect 399024 5568 399076 5574
rect 399024 5510 399076 5516
rect 397828 5432 397880 5438
rect 397828 5374 397880 5380
rect 396276 598 396672 626
rect 396644 480 396672 598
rect 397840 480 397868 5374
rect 399036 480 399064 5510
rect 400140 4282 400168 117370
rect 400968 109018 400996 118458
rect 400876 108990 400996 109018
rect 400876 106282 400904 108990
rect 400588 106276 400640 106282
rect 400588 106218 400640 106224
rect 400864 106276 400916 106282
rect 400864 106218 400916 106224
rect 400600 96694 400628 106218
rect 400588 96688 400640 96694
rect 400588 96630 400640 96636
rect 400772 96688 400824 96694
rect 400772 96630 400824 96636
rect 400784 91798 400812 96630
rect 400772 91792 400824 91798
rect 400772 91734 400824 91740
rect 401048 91792 401100 91798
rect 401048 91734 401100 91740
rect 401060 86986 401088 91734
rect 400968 86958 401088 86986
rect 400968 85542 400996 86958
rect 400772 85536 400824 85542
rect 400772 85478 400824 85484
rect 400956 85536 401008 85542
rect 400956 85478 401008 85484
rect 400784 77058 400812 85478
rect 400784 77030 400996 77058
rect 400968 70446 400996 77030
rect 400956 70440 401008 70446
rect 400956 70382 401008 70388
rect 401048 70372 401100 70378
rect 401048 70314 401100 70320
rect 401060 67658 401088 70314
rect 400956 67652 401008 67658
rect 400956 67594 401008 67600
rect 401048 67652 401100 67658
rect 401048 67594 401100 67600
rect 400968 56642 400996 67594
rect 400772 56636 400824 56642
rect 400772 56578 400824 56584
rect 400956 56636 401008 56642
rect 400956 56578 401008 56584
rect 400784 38622 400812 56578
rect 400588 38616 400640 38622
rect 400588 38558 400640 38564
rect 400772 38616 400824 38622
rect 400772 38558 400824 38564
rect 400600 29034 400628 38558
rect 400588 29028 400640 29034
rect 400588 28970 400640 28976
rect 400864 29028 400916 29034
rect 400864 28970 400916 28976
rect 400876 22114 400904 28970
rect 400876 22086 401088 22114
rect 401060 19310 401088 22086
rect 400772 19304 400824 19310
rect 400772 19246 400824 19252
rect 401048 19304 401100 19310
rect 401048 19246 401100 19252
rect 400784 9722 400812 19246
rect 400772 9716 400824 9722
rect 400772 9658 400824 9664
rect 400956 9716 401008 9722
rect 400956 9658 401008 9664
rect 400128 4276 400180 4282
rect 400128 4218 400180 4224
rect 400220 3732 400272 3738
rect 400220 3674 400272 3680
rect 400232 480 400260 3674
rect 400968 814 400996 9658
rect 401324 5364 401376 5370
rect 401324 5306 401376 5312
rect 400956 808 401008 814
rect 400956 750 401008 756
rect 401336 480 401364 5306
rect 401520 4350 401548 120006
rect 402164 117366 402192 120006
rect 402152 117360 402204 117366
rect 402152 117302 402204 117308
rect 402796 117360 402848 117366
rect 402796 117302 402848 117308
rect 402520 8016 402572 8022
rect 402520 7958 402572 7964
rect 401508 4344 401560 4350
rect 401508 4286 401560 4292
rect 402532 480 402560 7958
rect 402808 6390 402836 117302
rect 402796 6384 402848 6390
rect 402796 6326 402848 6332
rect 402900 3942 402928 120006
rect 403360 117366 403388 120006
rect 403682 119762 403710 120020
rect 404234 119762 404262 120020
rect 404892 120006 405228 120034
rect 403682 119734 403756 119762
rect 404234 119734 404308 119762
rect 403348 117360 403400 117366
rect 403348 117302 403400 117308
rect 403728 114578 403756 119734
rect 404280 118522 404308 119734
rect 404268 118516 404320 118522
rect 404268 118458 404320 118464
rect 404360 117700 404412 117706
rect 404360 117642 404412 117648
rect 404268 117360 404320 117366
rect 404268 117302 404320 117308
rect 403716 114572 403768 114578
rect 403716 114514 403768 114520
rect 403900 114572 403952 114578
rect 403900 114514 403952 114520
rect 403912 109070 403940 114514
rect 403900 109064 403952 109070
rect 403900 109006 403952 109012
rect 403992 108996 404044 109002
rect 403992 108938 404044 108944
rect 404004 106282 404032 108938
rect 403992 106276 404044 106282
rect 403992 106218 404044 106224
rect 404084 106276 404136 106282
rect 404084 106218 404136 106224
rect 404096 99362 404124 106218
rect 403912 99334 404124 99362
rect 403912 96642 403940 99334
rect 403912 96626 404032 96642
rect 403716 96620 403768 96626
rect 403912 96620 404044 96626
rect 403912 96614 403992 96620
rect 403716 96562 403768 96568
rect 403992 96562 404044 96568
rect 403728 87038 403756 96562
rect 404004 96531 404032 96562
rect 403716 87032 403768 87038
rect 403716 86974 403768 86980
rect 403900 87032 403952 87038
rect 403900 86974 403952 86980
rect 403912 86902 403940 86974
rect 403900 86896 403952 86902
rect 403900 86838 403952 86844
rect 403992 86896 404044 86902
rect 403992 86838 404044 86844
rect 404004 71210 404032 86838
rect 403820 71182 404032 71210
rect 403820 66298 403848 71182
rect 403808 66292 403860 66298
rect 403808 66234 403860 66240
rect 404084 66292 404136 66298
rect 404084 66234 404136 66240
rect 404096 66178 404124 66234
rect 404096 66150 404216 66178
rect 404188 60602 404216 66150
rect 404004 60574 404216 60602
rect 404004 56574 404032 60574
rect 403808 56568 403860 56574
rect 403808 56510 403860 56516
rect 403992 56568 404044 56574
rect 403992 56510 404044 56516
rect 403820 46986 403848 56510
rect 403808 46980 403860 46986
rect 403808 46922 403860 46928
rect 404084 46980 404136 46986
rect 404084 46922 404136 46928
rect 404096 43602 404124 46922
rect 404004 43574 404124 43602
rect 404004 42106 404032 43574
rect 404004 42078 404124 42106
rect 404096 31822 404124 42078
rect 404084 31816 404136 31822
rect 404084 31758 404136 31764
rect 404084 31680 404136 31686
rect 404084 31622 404136 31628
rect 404096 21978 404124 31622
rect 404096 21950 404216 21978
rect 404188 6322 404216 21950
rect 404176 6316 404228 6322
rect 404176 6258 404228 6264
rect 404280 4418 404308 117302
rect 404372 117230 404400 117642
rect 405200 117366 405228 120006
rect 405522 119762 405550 120020
rect 406088 120006 406424 120034
rect 406732 120006 406976 120034
rect 407376 120006 407712 120034
rect 407928 120006 408264 120034
rect 408572 120006 408908 120034
rect 409216 120006 409368 120034
rect 405522 119734 405596 119762
rect 405188 117360 405240 117366
rect 405188 117302 405240 117308
rect 404360 117224 404412 117230
rect 404360 117166 404412 117172
rect 405568 6186 405596 119734
rect 406396 117366 406424 120006
rect 405648 117360 405700 117366
rect 405648 117302 405700 117308
rect 406384 117360 406436 117366
rect 406384 117302 406436 117308
rect 405556 6180 405608 6186
rect 405556 6122 405608 6128
rect 404912 5296 404964 5302
rect 404912 5238 404964 5244
rect 404268 4412 404320 4418
rect 404268 4354 404320 4360
rect 402888 3936 402940 3942
rect 402888 3878 402940 3884
rect 403716 808 403768 814
rect 403716 750 403768 756
rect 403728 480 403756 750
rect 404924 480 404952 5238
rect 405660 4486 405688 117302
rect 406108 7948 406160 7954
rect 406108 7890 406160 7896
rect 405648 4480 405700 4486
rect 405648 4422 405700 4428
rect 406120 480 406148 7890
rect 406948 4554 406976 120006
rect 407684 117366 407712 120006
rect 408236 118590 408264 120006
rect 408224 118584 408276 118590
rect 408224 118526 408276 118532
rect 407764 117904 407816 117910
rect 407764 117846 407816 117852
rect 407028 117360 407080 117366
rect 407028 117302 407080 117308
rect 407672 117360 407724 117366
rect 407672 117302 407724 117308
rect 406936 4548 406988 4554
rect 406936 4490 406988 4496
rect 407040 3942 407068 117302
rect 407028 3936 407080 3942
rect 407028 3878 407080 3884
rect 407776 3670 407804 117846
rect 408880 117366 408908 120006
rect 408408 117360 408460 117366
rect 408408 117302 408460 117308
rect 408868 117360 408920 117366
rect 408868 117302 408920 117308
rect 408420 6254 408448 117302
rect 409340 114646 409368 120006
rect 409754 119762 409782 120020
rect 410412 120006 410748 120034
rect 409754 119734 409828 119762
rect 409696 117360 409748 117366
rect 409696 117302 409748 117308
rect 409328 114640 409380 114646
rect 409328 114582 409380 114588
rect 409604 114640 409656 114646
rect 409604 114582 409656 114588
rect 409616 114510 409644 114582
rect 409420 114504 409472 114510
rect 409420 114446 409472 114452
rect 409604 114504 409656 114510
rect 409604 114446 409656 114452
rect 409432 104922 409460 114446
rect 409328 104916 409380 104922
rect 409328 104858 409380 104864
rect 409420 104916 409472 104922
rect 409420 104858 409472 104864
rect 409340 95266 409368 104858
rect 409328 95260 409380 95266
rect 409328 95202 409380 95208
rect 409604 95260 409656 95266
rect 409604 95202 409656 95208
rect 409616 95146 409644 95202
rect 409524 95118 409644 95146
rect 409524 89758 409552 95118
rect 409512 89752 409564 89758
rect 409512 89694 409564 89700
rect 409604 89684 409656 89690
rect 409604 89626 409656 89632
rect 409616 67658 409644 89626
rect 409512 67652 409564 67658
rect 409512 67594 409564 67600
rect 409604 67652 409656 67658
rect 409604 67594 409656 67600
rect 409524 66230 409552 67594
rect 409420 66224 409472 66230
rect 409420 66166 409472 66172
rect 409512 66224 409564 66230
rect 409512 66166 409564 66172
rect 409432 56642 409460 66166
rect 409328 56636 409380 56642
rect 409328 56578 409380 56584
rect 409420 56636 409472 56642
rect 409420 56578 409472 56584
rect 409340 51066 409368 56578
rect 409328 51060 409380 51066
rect 409328 51002 409380 51008
rect 409512 51060 409564 51066
rect 409512 51002 409564 51008
rect 409524 41290 409552 51002
rect 409524 41262 409644 41290
rect 409616 38622 409644 41262
rect 409328 38616 409380 38622
rect 409328 38558 409380 38564
rect 409604 38616 409656 38622
rect 409604 38558 409656 38564
rect 409340 29034 409368 38558
rect 409328 29028 409380 29034
rect 409328 28970 409380 28976
rect 409420 29028 409472 29034
rect 409420 28970 409472 28976
rect 409432 19378 409460 28970
rect 409420 19372 409472 19378
rect 409420 19314 409472 19320
rect 409604 19372 409656 19378
rect 409604 19314 409656 19320
rect 409512 9104 409564 9110
rect 409512 9046 409564 9052
rect 408408 6248 408460 6254
rect 408408 6190 408460 6196
rect 408500 5228 408552 5234
rect 408500 5170 408552 5176
rect 407304 3664 407356 3670
rect 407304 3606 407356 3612
rect 407764 3664 407816 3670
rect 407764 3606 407816 3612
rect 407316 480 407344 3606
rect 408512 480 408540 5170
rect 409524 3874 409552 9046
rect 409616 8158 409644 19314
rect 409708 8514 409736 117302
rect 409800 9110 409828 119734
rect 410720 117366 410748 120006
rect 411042 119762 411070 120020
rect 411608 120006 411944 120034
rect 412252 120006 412588 120034
rect 412896 120006 413232 120034
rect 413448 120006 413784 120034
rect 414092 120006 414428 120034
rect 411042 119734 411116 119762
rect 410708 117360 410760 117366
rect 410708 117302 410760 117308
rect 410524 117224 410576 117230
rect 410524 117166 410576 117172
rect 409788 9104 409840 9110
rect 409788 9046 409840 9052
rect 409708 8486 409828 8514
rect 409604 8152 409656 8158
rect 409604 8094 409656 8100
rect 409696 7880 409748 7886
rect 409696 7822 409748 7828
rect 409512 3868 409564 3874
rect 409512 3810 409564 3816
rect 409708 480 409736 7822
rect 409800 4622 409828 8486
rect 409788 4616 409840 4622
rect 409788 4558 409840 4564
rect 410536 3058 410564 117166
rect 411088 8090 411116 119734
rect 411916 117774 411944 120006
rect 411904 117768 411956 117774
rect 411904 117710 411956 117716
rect 411168 117360 411220 117366
rect 411168 117302 411220 117308
rect 411076 8084 411128 8090
rect 411076 8026 411128 8032
rect 411180 4690 411208 117302
rect 412088 5160 412140 5166
rect 412088 5102 412140 5108
rect 411168 4684 411220 4690
rect 411168 4626 411220 4632
rect 410892 3664 410944 3670
rect 410892 3606 410944 3612
rect 410524 3052 410576 3058
rect 410524 2994 410576 3000
rect 410904 480 410932 3606
rect 412100 480 412128 5102
rect 412560 4758 412588 120006
rect 413204 117366 413232 120006
rect 413756 117502 413784 120006
rect 413744 117496 413796 117502
rect 413744 117438 413796 117444
rect 414400 117366 414428 120006
rect 414722 119762 414750 120020
rect 415274 119762 415302 120020
rect 415932 120006 416268 120034
rect 414722 119734 414796 119762
rect 415274 119734 415348 119762
rect 414664 117496 414716 117502
rect 414664 117438 414716 117444
rect 413192 117360 413244 117366
rect 413192 117302 413244 117308
rect 413928 117360 413980 117366
rect 413928 117302 413980 117308
rect 414388 117360 414440 117366
rect 414388 117302 414440 117308
rect 413940 8022 413968 117302
rect 413928 8016 413980 8022
rect 413928 7958 413980 7964
rect 413284 7812 413336 7818
rect 413284 7754 413336 7760
rect 412548 4752 412600 4758
rect 412548 4694 412600 4700
rect 413296 480 413324 7754
rect 414676 3806 414704 117438
rect 414768 113218 414796 119734
rect 415320 117706 415348 119734
rect 415308 117700 415360 117706
rect 415308 117642 415360 117648
rect 416240 117366 416268 120006
rect 416562 119762 416590 120020
rect 417128 120006 417464 120034
rect 417772 120006 418108 120034
rect 418324 120006 418660 120034
rect 418968 120006 419304 120034
rect 419612 120006 419948 120034
rect 420164 120006 420316 120034
rect 416562 119734 416636 119762
rect 415308 117360 415360 117366
rect 415308 117302 415360 117308
rect 416228 117360 416280 117366
rect 416228 117302 416280 117308
rect 414756 113212 414808 113218
rect 414756 113154 414808 113160
rect 415216 113212 415268 113218
rect 415216 113154 415268 113160
rect 415228 106350 415256 113154
rect 415216 106344 415268 106350
rect 415216 106286 415268 106292
rect 415216 106208 415268 106214
rect 415216 106150 415268 106156
rect 415228 104802 415256 106150
rect 415136 104774 415256 104802
rect 415136 103494 415164 104774
rect 414940 103488 414992 103494
rect 414940 103430 414992 103436
rect 415124 103488 415176 103494
rect 415124 103430 415176 103436
rect 414952 94602 414980 103430
rect 414952 94574 415164 94602
rect 415136 89758 415164 94574
rect 415124 89752 415176 89758
rect 415124 89694 415176 89700
rect 415124 89616 415176 89622
rect 415124 89558 415176 89564
rect 415136 84182 415164 89558
rect 415032 84176 415084 84182
rect 415032 84118 415084 84124
rect 415124 84176 415176 84182
rect 415124 84118 415176 84124
rect 415044 74594 415072 84118
rect 414940 74588 414992 74594
rect 414940 74530 414992 74536
rect 415032 74588 415084 74594
rect 415032 74530 415084 74536
rect 414952 66230 414980 74530
rect 414756 66224 414808 66230
rect 414756 66166 414808 66172
rect 414940 66224 414992 66230
rect 414940 66166 414992 66172
rect 414768 56642 414796 66166
rect 414756 56636 414808 56642
rect 414756 56578 414808 56584
rect 415216 56636 415268 56642
rect 415216 56578 415268 56584
rect 415228 48346 415256 56578
rect 414940 48340 414992 48346
rect 414940 48282 414992 48288
rect 415216 48340 415268 48346
rect 415216 48282 415268 48288
rect 414952 43466 414980 48282
rect 414952 43438 415164 43466
rect 415136 31822 415164 43438
rect 415124 31816 415176 31822
rect 415124 31758 415176 31764
rect 415032 31748 415084 31754
rect 415032 31690 415084 31696
rect 415044 29034 415072 31690
rect 415032 29028 415084 29034
rect 415032 28970 415084 28976
rect 415216 29028 415268 29034
rect 415216 28970 415268 28976
rect 415228 12458 415256 28970
rect 415136 12430 415256 12458
rect 415136 7954 415164 12430
rect 415124 7948 415176 7954
rect 415124 7890 415176 7896
rect 415320 5506 415348 117302
rect 416608 7886 416636 119734
rect 416964 118652 417016 118658
rect 416964 118594 417016 118600
rect 416688 117360 416740 117366
rect 416688 117302 416740 117308
rect 416596 7880 416648 7886
rect 416596 7822 416648 7828
rect 415308 5500 415360 5506
rect 415308 5442 415360 5448
rect 416700 5438 416728 117302
rect 416872 7744 416924 7750
rect 416872 7686 416924 7692
rect 416688 5432 416740 5438
rect 416688 5374 416740 5380
rect 415676 5092 415728 5098
rect 415676 5034 415728 5040
rect 414664 3800 414716 3806
rect 414664 3742 414716 3748
rect 414480 3528 414532 3534
rect 414480 3470 414532 3476
rect 414492 480 414520 3470
rect 415688 480 415716 5034
rect 416884 480 416912 7686
rect 416976 610 417004 118594
rect 417436 118454 417464 120006
rect 417424 118448 417476 118454
rect 417424 118390 417476 118396
rect 418080 5370 418108 120006
rect 418632 117366 418660 120006
rect 419276 117570 419304 120006
rect 419264 117564 419316 117570
rect 419264 117506 419316 117512
rect 419920 117366 419948 120006
rect 420184 117564 420236 117570
rect 420184 117506 420236 117512
rect 418620 117360 418672 117366
rect 418620 117302 418672 117308
rect 419448 117360 419500 117366
rect 419448 117302 419500 117308
rect 419908 117360 419960 117366
rect 419908 117302 419960 117308
rect 419460 7818 419488 117302
rect 419448 7812 419500 7818
rect 419448 7754 419500 7760
rect 418068 5364 418120 5370
rect 418068 5306 418120 5312
rect 419172 5024 419224 5030
rect 419172 4966 419224 4972
rect 416964 604 417016 610
rect 416964 546 417016 552
rect 417976 604 418028 610
rect 417976 546 418028 552
rect 417988 480 418016 546
rect 419184 480 419212 4966
rect 420196 3738 420224 117506
rect 420288 116006 420316 120006
rect 420794 119762 420822 120020
rect 421452 120006 421788 120034
rect 422004 120006 422156 120034
rect 422648 120006 422984 120034
rect 423292 120006 423536 120034
rect 423844 120006 424180 120034
rect 424488 120006 424824 120034
rect 425132 120006 425468 120034
rect 425684 120006 426020 120034
rect 420794 119734 420868 119762
rect 420840 117910 420868 119734
rect 420828 117904 420880 117910
rect 420828 117846 420880 117852
rect 421760 117434 421788 120006
rect 421748 117428 421800 117434
rect 421748 117370 421800 117376
rect 420828 117360 420880 117366
rect 420828 117302 420880 117308
rect 420276 116000 420328 116006
rect 420276 115942 420328 115948
rect 420460 116000 420512 116006
rect 420460 115942 420512 115948
rect 420472 109018 420500 115942
rect 420472 108990 420684 109018
rect 420656 104854 420684 108990
rect 420552 104848 420604 104854
rect 420552 104790 420604 104796
rect 420644 104848 420696 104854
rect 420644 104790 420696 104796
rect 420564 95266 420592 104790
rect 420552 95260 420604 95266
rect 420552 95202 420604 95208
rect 420736 95260 420788 95266
rect 420736 95202 420788 95208
rect 420748 86986 420776 95202
rect 420656 86970 420776 86986
rect 420552 86964 420604 86970
rect 420552 86906 420604 86912
rect 420644 86964 420776 86970
rect 420696 86958 420776 86964
rect 420644 86906 420696 86912
rect 420564 77382 420592 86906
rect 420552 77376 420604 77382
rect 420552 77318 420604 77324
rect 420736 77376 420788 77382
rect 420736 77318 420788 77324
rect 420748 77217 420776 77318
rect 420734 77208 420790 77217
rect 420734 77143 420790 77152
rect 420644 67652 420696 67658
rect 420644 67594 420696 67600
rect 420656 67538 420684 67594
rect 420656 67510 420776 67538
rect 420748 60790 420776 67510
rect 420736 60784 420788 60790
rect 420736 60726 420788 60732
rect 420644 60716 420696 60722
rect 420644 60658 420696 60664
rect 420656 58018 420684 60658
rect 420656 57990 420776 58018
rect 420748 57934 420776 57990
rect 420460 57928 420512 57934
rect 420460 57870 420512 57876
rect 420736 57928 420788 57934
rect 420736 57870 420788 57876
rect 420472 48385 420500 57870
rect 420458 48376 420514 48385
rect 420458 48311 420514 48320
rect 420642 48376 420698 48385
rect 420642 48311 420698 48320
rect 420656 48278 420684 48311
rect 420552 48272 420604 48278
rect 420552 48214 420604 48220
rect 420644 48272 420696 48278
rect 420644 48214 420696 48220
rect 420564 41290 420592 48214
rect 420564 41262 420684 41290
rect 420656 33862 420684 41262
rect 420460 33856 420512 33862
rect 420460 33798 420512 33804
rect 420644 33856 420696 33862
rect 420644 33798 420696 33804
rect 420472 29073 420500 33798
rect 420458 29064 420514 29073
rect 420458 28999 420514 29008
rect 420642 29030 420698 29039
rect 420552 28960 420604 28966
rect 420642 28965 420698 28974
rect 420552 28902 420604 28908
rect 420644 28960 420696 28965
rect 420644 28902 420696 28908
rect 420564 21978 420592 28902
rect 420564 21950 420684 21978
rect 420656 14550 420684 21950
rect 420460 14544 420512 14550
rect 420460 14486 420512 14492
rect 420644 14544 420696 14550
rect 420644 14486 420696 14492
rect 420472 9722 420500 14486
rect 420460 9716 420512 9722
rect 420460 9658 420512 9664
rect 420644 9716 420696 9722
rect 420644 9658 420696 9664
rect 420656 7750 420684 9658
rect 420644 7744 420696 7750
rect 420644 7686 420696 7692
rect 420368 7676 420420 7682
rect 420368 7618 420420 7624
rect 420184 3732 420236 3738
rect 420184 3674 420236 3680
rect 420380 480 420408 7618
rect 420840 5302 420868 117302
rect 421010 77208 421066 77217
rect 421010 77143 421066 77152
rect 421024 67658 421052 77143
rect 421012 67652 421064 67658
rect 421012 67594 421064 67600
rect 422128 7682 422156 120006
rect 422852 118448 422904 118454
rect 422852 118390 422904 118396
rect 422864 117842 422892 118390
rect 422852 117836 422904 117842
rect 422852 117778 422904 117784
rect 422208 117428 422260 117434
rect 422208 117370 422260 117376
rect 422116 7676 422168 7682
rect 422116 7618 422168 7624
rect 420828 5296 420880 5302
rect 420828 5238 420880 5244
rect 422220 5234 422248 117370
rect 422956 117366 422984 120006
rect 422944 117360 422996 117366
rect 422944 117302 422996 117308
rect 422208 5228 422260 5234
rect 422208 5170 422260 5176
rect 423508 5098 423536 120006
rect 424152 117366 424180 120006
rect 424796 118658 424824 120006
rect 424784 118652 424836 118658
rect 424784 118594 424836 118600
rect 425336 117632 425388 117638
rect 425336 117574 425388 117580
rect 423588 117360 423640 117366
rect 423588 117302 423640 117308
rect 424140 117360 424192 117366
rect 424140 117302 424192 117308
rect 424968 117360 425020 117366
rect 424968 117302 425020 117308
rect 423496 5092 423548 5098
rect 423496 5034 423548 5040
rect 422760 4956 422812 4962
rect 422760 4898 422812 4904
rect 421564 3460 421616 3466
rect 421564 3402 421616 3408
rect 421576 480 421604 3402
rect 422772 480 422800 4898
rect 423600 3670 423628 117302
rect 424980 7614 425008 117302
rect 423956 7608 424008 7614
rect 423956 7550 424008 7556
rect 424968 7608 425020 7614
rect 424968 7550 425020 7556
rect 423588 3664 423640 3670
rect 423588 3606 423640 3612
rect 423968 480 423996 7550
rect 425348 610 425376 117574
rect 425440 117366 425468 120006
rect 425428 117360 425480 117366
rect 425428 117302 425480 117308
rect 425992 114510 426020 120006
rect 426314 119762 426342 120020
rect 426972 120006 427308 120034
rect 427524 120006 427676 120034
rect 428168 120006 428504 120034
rect 428812 120006 429148 120034
rect 429364 120006 429700 120034
rect 430008 120006 430344 120034
rect 430652 120006 430988 120034
rect 431204 120006 431356 120034
rect 426314 119734 426388 119762
rect 426360 117502 426388 119734
rect 426348 117496 426400 117502
rect 426348 117438 426400 117444
rect 427280 117366 427308 120006
rect 426348 117360 426400 117366
rect 426348 117302 426400 117308
rect 427268 117360 427320 117366
rect 427268 117302 427320 117308
rect 425980 114504 426032 114510
rect 425980 114446 426032 114452
rect 426164 114436 426216 114442
rect 426164 114378 426216 114384
rect 426176 104854 426204 114378
rect 425980 104848 426032 104854
rect 425980 104790 426032 104796
rect 426164 104848 426216 104854
rect 426164 104790 426216 104796
rect 425992 87009 426020 104790
rect 425978 87000 426034 87009
rect 425978 86935 426034 86944
rect 426162 87000 426218 87009
rect 426162 86935 426218 86944
rect 426176 80714 426204 86935
rect 426072 80708 426124 80714
rect 426072 80650 426124 80656
rect 426164 80708 426216 80714
rect 426164 80650 426216 80656
rect 426084 74526 426112 80650
rect 426072 74520 426124 74526
rect 426072 74462 426124 74468
rect 426070 64968 426126 64977
rect 426070 64903 426126 64912
rect 426084 64870 426112 64903
rect 425980 64864 426032 64870
rect 425980 64806 426032 64812
rect 426072 64864 426124 64870
rect 426072 64806 426124 64812
rect 425992 55350 426020 64806
rect 425980 55344 426032 55350
rect 425980 55286 426032 55292
rect 426072 55344 426124 55350
rect 426072 55286 426124 55292
rect 426084 55214 426112 55286
rect 425796 55208 425848 55214
rect 425796 55150 425848 55156
rect 426072 55208 426124 55214
rect 426072 55150 426124 55156
rect 425808 45626 425836 55150
rect 425796 45620 425848 45626
rect 425796 45562 425848 45568
rect 425980 45620 426032 45626
rect 425980 45562 426032 45568
rect 425992 45490 426020 45562
rect 425796 45484 425848 45490
rect 425796 45426 425848 45432
rect 425980 45484 426032 45490
rect 425980 45426 426032 45432
rect 425808 44169 425836 45426
rect 425794 44160 425850 44169
rect 425794 44095 425850 44104
rect 425978 44160 426034 44169
rect 425978 44095 426034 44104
rect 425992 34542 426020 44095
rect 425980 34536 426032 34542
rect 425980 34478 426032 34484
rect 426072 34536 426124 34542
rect 426072 34478 426124 34484
rect 426084 24818 426112 34478
rect 426072 24812 426124 24818
rect 426072 24754 426124 24760
rect 426164 24812 426216 24818
rect 426164 24754 426216 24760
rect 426176 9178 426204 24754
rect 426164 9172 426216 9178
rect 426164 9114 426216 9120
rect 426360 5166 426388 117302
rect 426440 74520 426492 74526
rect 426440 74462 426492 74468
rect 426452 64977 426480 74462
rect 426438 64968 426494 64977
rect 426438 64903 426494 64912
rect 427648 9042 427676 120006
rect 428476 117638 428504 120006
rect 428464 117632 428516 117638
rect 428464 117574 428516 117580
rect 427728 117360 427780 117366
rect 427728 117302 427780 117308
rect 427544 9036 427596 9042
rect 427544 8978 427596 8984
rect 427636 9036 427688 9042
rect 427636 8978 427688 8984
rect 426348 5160 426400 5166
rect 426348 5102 426400 5108
rect 426348 4888 426400 4894
rect 426348 4830 426400 4836
rect 425152 604 425204 610
rect 425152 546 425204 552
rect 425336 604 425388 610
rect 425336 546 425388 552
rect 425164 480 425192 546
rect 426360 480 426388 4830
rect 427556 480 427584 8978
rect 427740 5030 427768 117302
rect 427728 5024 427780 5030
rect 427728 4966 427780 4972
rect 429120 4962 429148 120006
rect 429672 117366 429700 120006
rect 430316 117570 430344 120006
rect 430304 117564 430356 117570
rect 430304 117506 430356 117512
rect 429844 117496 429896 117502
rect 429844 117438 429896 117444
rect 429660 117360 429712 117366
rect 429660 117302 429712 117308
rect 429108 4956 429160 4962
rect 429108 4898 429160 4904
rect 429856 3602 429884 117438
rect 430960 117366 430988 120006
rect 431224 117564 431276 117570
rect 431224 117506 431276 117512
rect 430488 117360 430540 117366
rect 430488 117302 430540 117308
rect 430948 117360 431000 117366
rect 430948 117302 431000 117308
rect 430500 9110 430528 117302
rect 430488 9104 430540 9110
rect 430488 9046 430540 9052
rect 431132 8968 431184 8974
rect 431132 8910 431184 8916
rect 429936 4820 429988 4826
rect 429936 4762 429988 4768
rect 428740 3596 428792 3602
rect 428740 3538 428792 3544
rect 429844 3596 429896 3602
rect 429844 3538 429896 3544
rect 428752 480 428780 3538
rect 429948 480 429976 4762
rect 431144 480 431172 8910
rect 431236 3466 431264 117506
rect 431328 114753 431356 120006
rect 431834 119762 431862 120020
rect 432492 120006 432828 120034
rect 433044 120006 433196 120034
rect 433688 120006 434024 120034
rect 431788 119734 431862 119762
rect 431788 118454 431816 119734
rect 431776 118448 431828 118454
rect 431776 118390 431828 118396
rect 432800 117366 432828 120006
rect 431868 117360 431920 117366
rect 431868 117302 431920 117308
rect 432788 117360 432840 117366
rect 432788 117302 432840 117308
rect 431314 114744 431370 114753
rect 431314 114679 431370 114688
rect 431590 114608 431646 114617
rect 431590 114543 431646 114552
rect 431604 114510 431632 114543
rect 431592 114504 431644 114510
rect 431592 114446 431644 114452
rect 431684 114504 431736 114510
rect 431684 114446 431736 114452
rect 431696 106350 431724 114446
rect 431684 106344 431736 106350
rect 431684 106286 431736 106292
rect 431592 106276 431644 106282
rect 431592 106218 431644 106224
rect 431604 104938 431632 106218
rect 431604 104910 431724 104938
rect 431696 104854 431724 104910
rect 431408 104848 431460 104854
rect 431408 104790 431460 104796
rect 431684 104848 431736 104854
rect 431684 104790 431736 104796
rect 431420 95198 431448 104790
rect 431408 95192 431460 95198
rect 431408 95134 431460 95140
rect 431500 95192 431552 95198
rect 431500 95134 431552 95140
rect 431512 85610 431540 95134
rect 431500 85604 431552 85610
rect 431500 85546 431552 85552
rect 431592 85604 431644 85610
rect 431592 85546 431644 85552
rect 431604 80102 431632 85546
rect 431788 80102 431816 80133
rect 431592 80096 431644 80102
rect 431776 80096 431828 80102
rect 431644 80044 431776 80050
rect 431592 80038 431828 80044
rect 431604 80022 431816 80038
rect 431604 75886 431632 80022
rect 431592 75880 431644 75886
rect 431592 75822 431644 75828
rect 431776 75880 431828 75886
rect 431776 75822 431828 75828
rect 431788 66337 431816 75822
rect 431590 66328 431646 66337
rect 431590 66263 431646 66272
rect 431774 66328 431830 66337
rect 431774 66263 431830 66272
rect 431604 64870 431632 66263
rect 431408 64864 431460 64870
rect 431408 64806 431460 64812
rect 431592 64864 431644 64870
rect 431592 64806 431644 64812
rect 431420 55282 431448 64806
rect 431408 55276 431460 55282
rect 431408 55218 431460 55224
rect 431592 55276 431644 55282
rect 431592 55218 431644 55224
rect 431604 45558 431632 55218
rect 431500 45552 431552 45558
rect 431500 45494 431552 45500
rect 431592 45552 431644 45558
rect 431592 45494 431644 45500
rect 431512 35970 431540 45494
rect 431408 35964 431460 35970
rect 431408 35906 431460 35912
rect 431500 35964 431552 35970
rect 431500 35906 431552 35912
rect 431420 27674 431448 35906
rect 431408 27668 431460 27674
rect 431408 27610 431460 27616
rect 431684 27668 431736 27674
rect 431684 27610 431736 27616
rect 431696 22114 431724 27610
rect 431696 22086 431816 22114
rect 431788 12458 431816 22086
rect 431696 12430 431816 12458
rect 431696 8974 431724 12430
rect 431684 8968 431736 8974
rect 431684 8910 431736 8916
rect 431880 4894 431908 117302
rect 433168 10334 433196 120006
rect 433996 117366 434024 120006
rect 433248 117360 433300 117366
rect 433248 117302 433300 117308
rect 433984 117360 434036 117366
rect 433984 117302 434036 117308
rect 433156 10328 433208 10334
rect 433156 10270 433208 10276
rect 431868 4888 431920 4894
rect 431868 4830 431920 4836
rect 433260 4826 433288 117302
rect 436296 35902 436324 192918
rect 436388 80034 436416 196143
rect 436466 194032 436522 194041
rect 436466 193967 436522 193976
rect 436480 120630 436508 193967
rect 436572 176225 436600 201078
rect 436664 177993 436692 201146
rect 436744 201068 436796 201074
rect 436744 201010 436796 201016
rect 436756 182073 436784 201010
rect 436834 198928 436890 198937
rect 436834 198863 436890 198872
rect 436848 192982 436876 198863
rect 436836 192976 436888 192982
rect 436836 192918 436888 192924
rect 436742 182064 436798 182073
rect 436742 181999 436798 182008
rect 436650 177984 436706 177993
rect 436650 177919 436706 177928
rect 436558 176216 436614 176225
rect 436558 176151 436614 176160
rect 438136 155650 438164 700606
rect 462332 700602 462360 703520
rect 462320 700596 462372 700602
rect 462320 700538 462372 700544
rect 478524 700534 478552 703520
rect 494808 700670 494836 703520
rect 494796 700664 494848 700670
rect 494796 700606 494848 700612
rect 478512 700528 478564 700534
rect 478512 700470 478564 700476
rect 442264 700460 442316 700466
rect 442264 700402 442316 700408
rect 440884 673532 440936 673538
rect 440884 673474 440936 673480
rect 439504 626612 439556 626618
rect 439504 626554 439556 626560
rect 438216 579692 438268 579698
rect 438216 579634 438268 579640
rect 438124 155644 438176 155650
rect 438124 155586 438176 155592
rect 437386 152280 437442 152289
rect 437386 152215 437442 152224
rect 437400 151978 437428 152215
rect 437388 151972 437440 151978
rect 437388 151914 437440 151920
rect 437020 150340 437072 150346
rect 437020 150282 437072 150288
rect 437032 150249 437060 150282
rect 437018 150240 437074 150249
rect 437018 150175 437074 150184
rect 438228 146266 438256 579634
rect 438308 485852 438360 485858
rect 438308 485794 438360 485800
rect 438216 146260 438268 146266
rect 438216 146202 438268 146208
rect 437388 144900 437440 144906
rect 437388 144842 437440 144848
rect 437400 144537 437428 144842
rect 437386 144528 437442 144537
rect 437386 144463 437442 144472
rect 438320 142118 438348 485794
rect 439516 148918 439544 626554
rect 440896 150346 440924 673474
rect 442276 151978 442304 700402
rect 527192 700398 527220 703520
rect 527180 700392 527232 700398
rect 527180 700334 527232 700340
rect 543476 700330 543504 703520
rect 559668 700466 559696 703520
rect 559656 700460 559708 700466
rect 559656 700402 559708 700408
rect 543464 700324 543516 700330
rect 543464 700266 543516 700272
rect 580170 698048 580226 698057
rect 580170 697983 580226 697992
rect 580184 696998 580212 697983
rect 580172 696992 580224 696998
rect 580172 696934 580224 696940
rect 580170 686352 580226 686361
rect 580170 686287 580226 686296
rect 580184 685914 580212 686287
rect 580172 685908 580224 685914
rect 580172 685850 580224 685856
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 580170 651128 580226 651137
rect 580170 651063 580226 651072
rect 580184 650078 580212 651063
rect 580172 650072 580224 650078
rect 580172 650014 580224 650020
rect 580170 639432 580226 639441
rect 580170 639367 580226 639376
rect 580184 638994 580212 639367
rect 580172 638988 580224 638994
rect 580172 638930 580224 638936
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 580170 604208 580226 604217
rect 580170 604143 580226 604152
rect 580184 603158 580212 604143
rect 580172 603152 580224 603158
rect 580172 603094 580224 603100
rect 580170 592512 580226 592521
rect 580170 592447 580226 592456
rect 580184 592074 580212 592447
rect 580172 592068 580224 592074
rect 580172 592010 580224 592016
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 579698 580212 580751
rect 580172 579692 580224 579698
rect 580172 579634 580224 579640
rect 580446 557288 580502 557297
rect 580446 557223 580502 557232
rect 511264 556300 511316 556306
rect 511264 556242 511316 556248
rect 484400 556232 484452 556238
rect 484400 556174 484452 556180
rect 484412 554676 484440 556174
rect 511276 554676 511304 556242
rect 580354 545592 580410 545601
rect 580354 545527 580410 545536
rect 580262 533896 580318 533905
rect 580262 533831 580318 533840
rect 478892 520118 480010 520146
rect 478892 498846 478920 520118
rect 506860 517546 506888 520132
rect 505744 517540 505796 517546
rect 505744 517482 505796 517488
rect 506848 517540 506900 517546
rect 506848 517482 506900 517488
rect 478880 498840 478932 498846
rect 478880 498782 478932 498788
rect 458824 389428 458876 389434
rect 458824 389370 458876 389376
rect 475844 389428 475896 389434
rect 475844 389370 475896 389376
rect 456798 375184 456854 375193
rect 456798 375119 456854 375128
rect 456812 374066 456840 375119
rect 456800 374060 456852 374066
rect 456800 374002 456852 374008
rect 457442 358048 457498 358057
rect 457442 357983 457498 357992
rect 457456 201958 457484 357983
rect 458836 202774 458864 389370
rect 464252 389360 464304 389366
rect 464252 389302 464304 389308
rect 464264 387532 464292 389302
rect 475856 387532 475884 389370
rect 487436 389292 487488 389298
rect 487436 389234 487488 389240
rect 487448 387532 487476 389234
rect 499028 389224 499080 389230
rect 499028 389166 499080 389172
rect 499040 387532 499068 389166
rect 504730 378448 504786 378457
rect 503732 378406 504730 378434
rect 503732 361434 503760 378406
rect 504730 378383 504786 378392
rect 503640 361406 503760 361434
rect 503640 360074 503668 361406
rect 504730 360496 504786 360505
rect 504376 360454 504730 360482
rect 503640 360046 503760 360074
rect 503732 359938 503760 360046
rect 503732 359910 503852 359938
rect 503824 350554 503852 359910
rect 504376 351914 504404 360454
rect 504730 360431 504786 360440
rect 504100 351886 504404 351914
rect 504100 350554 504128 351886
rect 503824 350526 504036 350554
rect 504100 350526 504220 350554
rect 504008 344978 504036 350526
rect 503916 344950 504036 344978
rect 503812 342032 503864 342038
rect 503812 341974 503864 341980
rect 503718 340912 503774 340921
rect 503718 340847 503774 340856
rect 460584 337618 460612 340068
rect 460572 337612 460624 337618
rect 460572 337554 460624 337560
rect 472176 337550 472204 340068
rect 472164 337544 472216 337550
rect 472164 337486 472216 337492
rect 483768 337482 483796 340068
rect 483756 337476 483808 337482
rect 483756 337418 483808 337424
rect 495360 337414 495388 340068
rect 495348 337408 495400 337414
rect 495348 337350 495400 337356
rect 503732 331378 503760 340847
rect 503640 331350 503760 331378
rect 503640 331226 503668 331350
rect 503628 331220 503680 331226
rect 503628 331162 503680 331168
rect 503824 331106 503852 341974
rect 503916 340921 503944 344950
rect 504192 342038 504220 350526
rect 504824 345092 504876 345098
rect 504824 345034 504876 345040
rect 504730 343632 504786 343641
rect 504730 343567 504786 343576
rect 504180 342032 504232 342038
rect 504180 341974 504232 341980
rect 503902 340912 503958 340921
rect 504744 340882 504772 343567
rect 503902 340847 503958 340856
rect 504732 340876 504784 340882
rect 504732 340818 504784 340824
rect 503904 340808 503956 340814
rect 503904 340750 503956 340756
rect 503732 331078 503852 331106
rect 503732 328438 503760 331078
rect 503536 328432 503588 328438
rect 503536 328374 503588 328380
rect 503720 328432 503772 328438
rect 503720 328374 503772 328380
rect 503548 318850 503576 328374
rect 503916 321745 503944 340750
rect 504836 332602 504864 345034
rect 504468 332574 504864 332602
rect 504468 331242 504496 332574
rect 503996 331220 504048 331226
rect 503996 331162 504048 331168
rect 504376 331214 504496 331242
rect 504008 323610 504036 331162
rect 503996 323604 504048 323610
rect 503996 323546 504048 323552
rect 504180 323604 504232 323610
rect 504180 323546 504232 323552
rect 503902 321736 503958 321745
rect 503902 321671 503958 321680
rect 503902 321464 503958 321473
rect 503902 321399 503958 321408
rect 503536 318844 503588 318850
rect 503536 318786 503588 318792
rect 503720 318844 503772 318850
rect 503720 318786 503772 318792
rect 503732 313954 503760 318786
rect 503444 313948 503496 313954
rect 503444 313890 503496 313896
rect 503720 313948 503772 313954
rect 503720 313890 503772 313896
rect 503456 309194 503484 313890
rect 503628 311908 503680 311914
rect 503628 311850 503680 311856
rect 503640 311778 503668 311850
rect 503628 311772 503680 311778
rect 503628 311714 503680 311720
rect 503444 309188 503496 309194
rect 503444 309130 503496 309136
rect 503812 309188 503864 309194
rect 503812 309130 503864 309136
rect 503824 292482 503852 309130
rect 503732 292454 503852 292482
rect 503732 283082 503760 292454
rect 503720 283076 503772 283082
rect 503720 283018 503772 283024
rect 503812 283008 503864 283014
rect 503812 282950 503864 282956
rect 503628 273352 503680 273358
rect 503628 273294 503680 273300
rect 503640 273222 503668 273294
rect 503628 273216 503680 273222
rect 503628 273158 503680 273164
rect 503720 263696 503772 263702
rect 503720 263638 503772 263644
rect 503732 263566 503760 263638
rect 503720 263560 503772 263566
rect 503720 263502 503772 263508
rect 503628 254040 503680 254046
rect 503628 253982 503680 253988
rect 503640 253910 503668 253982
rect 503628 253904 503680 253910
rect 503824 253858 503852 282950
rect 503628 253846 503680 253852
rect 503732 253830 503852 253858
rect 503732 244458 503760 253830
rect 503720 244452 503772 244458
rect 503720 244394 503772 244400
rect 503812 244384 503864 244390
rect 503812 244326 503864 244332
rect 503628 234728 503680 234734
rect 503628 234670 503680 234676
rect 503640 234598 503668 234670
rect 503628 234592 503680 234598
rect 503824 234546 503852 244326
rect 503628 234534 503680 234540
rect 503732 234518 503852 234546
rect 503732 225146 503760 234518
rect 503720 225140 503772 225146
rect 503720 225082 503772 225088
rect 503812 225072 503864 225078
rect 503812 225014 503864 225020
rect 503628 215416 503680 215422
rect 503628 215358 503680 215364
rect 503640 215286 503668 215358
rect 503628 215280 503680 215286
rect 503824 215234 503852 225014
rect 503628 215222 503680 215228
rect 503732 215206 503852 215234
rect 503732 205834 503760 215206
rect 503720 205828 503772 205834
rect 503720 205770 503772 205776
rect 503812 205760 503864 205766
rect 503812 205702 503864 205708
rect 503720 205692 503772 205698
rect 503720 205634 503772 205640
rect 458824 202768 458876 202774
rect 458824 202710 458876 202716
rect 503732 202230 503760 205634
rect 503824 202298 503852 205702
rect 503916 202366 503944 321399
rect 504192 318850 504220 323546
rect 503996 318844 504048 318850
rect 503996 318786 504048 318792
rect 504180 318844 504232 318850
rect 504180 318786 504232 318792
rect 504008 311914 504036 318786
rect 504376 318782 504404 331214
rect 504364 318776 504416 318782
rect 504364 318718 504416 318724
rect 504456 318776 504508 318782
rect 504456 318718 504508 318724
rect 503996 311908 504048 311914
rect 503996 311850 504048 311856
rect 503996 311772 504048 311778
rect 503996 311714 504048 311720
rect 504008 273358 504036 311714
rect 504468 309262 504496 318718
rect 504364 309256 504416 309262
rect 504364 309198 504416 309204
rect 504456 309256 504508 309262
rect 504456 309198 504508 309204
rect 504376 309126 504404 309198
rect 504180 309120 504232 309126
rect 504180 309062 504232 309068
rect 504364 309120 504416 309126
rect 504364 309062 504416 309068
rect 504192 299538 504220 309062
rect 504180 299532 504232 299538
rect 504180 299474 504232 299480
rect 504456 299532 504508 299538
rect 504456 299474 504508 299480
rect 504468 298110 504496 299474
rect 504456 298104 504508 298110
rect 504456 298046 504508 298052
rect 504732 298104 504784 298110
rect 504732 298046 504784 298052
rect 504744 288454 504772 298046
rect 504548 288448 504600 288454
rect 504548 288390 504600 288396
rect 504732 288448 504784 288454
rect 504732 288390 504784 288396
rect 504560 280242 504588 288390
rect 504468 280214 504588 280242
rect 504468 278730 504496 280214
rect 504456 278724 504508 278730
rect 504456 278666 504508 278672
rect 504548 278724 504600 278730
rect 504548 278666 504600 278672
rect 503996 273352 504048 273358
rect 503996 273294 504048 273300
rect 503996 273216 504048 273222
rect 503996 273158 504048 273164
rect 504008 263702 504036 273158
rect 503996 263696 504048 263702
rect 503996 263638 504048 263644
rect 503996 263560 504048 263566
rect 503996 263502 504048 263508
rect 504008 254046 504036 263502
rect 504560 260953 504588 278666
rect 504270 260944 504326 260953
rect 504270 260879 504326 260888
rect 504546 260944 504602 260953
rect 504546 260879 504602 260888
rect 504284 260846 504312 260879
rect 504272 260840 504324 260846
rect 504272 260782 504324 260788
rect 504548 260840 504600 260846
rect 504548 260782 504600 260788
rect 503996 254040 504048 254046
rect 503996 253982 504048 253988
rect 503996 253904 504048 253910
rect 503996 253846 504048 253852
rect 504008 234734 504036 253846
rect 504560 253842 504588 260782
rect 504272 253836 504324 253842
rect 504272 253778 504324 253784
rect 504548 253836 504600 253842
rect 504548 253778 504600 253784
rect 504284 251190 504312 253778
rect 504088 251184 504140 251190
rect 504088 251126 504140 251132
rect 504272 251184 504324 251190
rect 504272 251126 504324 251132
rect 504100 241534 504128 251126
rect 504088 241528 504140 241534
rect 504088 241470 504140 241476
rect 504456 241528 504508 241534
rect 504456 241470 504508 241476
rect 504468 234734 504496 241470
rect 503996 234728 504048 234734
rect 503996 234670 504048 234676
rect 504456 234728 504508 234734
rect 504456 234670 504508 234676
rect 503996 234592 504048 234598
rect 503996 234534 504048 234540
rect 504364 234592 504416 234598
rect 504364 234534 504416 234540
rect 504008 215422 504036 234534
rect 504376 231810 504404 234534
rect 504180 231804 504232 231810
rect 504180 231746 504232 231752
rect 504364 231804 504416 231810
rect 504364 231746 504416 231752
rect 504192 222222 504220 231746
rect 504180 222216 504232 222222
rect 504180 222158 504232 222164
rect 504456 222216 504508 222222
rect 504456 222158 504508 222164
rect 504468 215422 504496 222158
rect 503996 215416 504048 215422
rect 503996 215358 504048 215364
rect 504456 215416 504508 215422
rect 504456 215358 504508 215364
rect 503996 215280 504048 215286
rect 503996 215222 504048 215228
rect 504272 215280 504324 215286
rect 504272 215222 504324 215228
rect 504008 205698 504036 215222
rect 504284 212514 504312 215222
rect 504192 212486 504312 212514
rect 504192 205698 504220 212486
rect 503996 205692 504048 205698
rect 503996 205634 504048 205640
rect 504180 205692 504232 205698
rect 504180 205634 504232 205640
rect 504272 205624 504324 205630
rect 504272 205566 504324 205572
rect 504284 202910 504312 205566
rect 504180 202904 504232 202910
rect 504180 202846 504232 202852
rect 504272 202904 504324 202910
rect 504272 202846 504324 202852
rect 503904 202360 503956 202366
rect 503904 202302 503956 202308
rect 503812 202292 503864 202298
rect 503812 202234 503864 202240
rect 503720 202224 503772 202230
rect 503720 202166 503772 202172
rect 457444 201952 457496 201958
rect 457444 201894 457496 201900
rect 504192 201278 504220 202846
rect 505756 202162 505784 517482
rect 579894 498672 579950 498681
rect 579894 498607 579950 498616
rect 579908 498234 579936 498607
rect 579896 498228 579948 498234
rect 579896 498170 579948 498176
rect 580170 486840 580226 486849
rect 580170 486775 580226 486784
rect 580184 485858 580212 486775
rect 580172 485852 580224 485858
rect 580172 485794 580224 485800
rect 580170 463448 580226 463457
rect 580170 463383 580226 463392
rect 580184 462398 580212 463383
rect 580172 462392 580224 462398
rect 580172 462334 580224 462340
rect 579894 451752 579950 451761
rect 579894 451687 579950 451696
rect 579908 451314 579936 451687
rect 579896 451308 579948 451314
rect 579896 451250 579948 451256
rect 579802 416528 579858 416537
rect 579802 416463 579858 416472
rect 579816 415478 579844 416463
rect 579804 415472 579856 415478
rect 579804 415414 579856 415420
rect 579986 346080 580042 346089
rect 579986 346015 580042 346024
rect 580000 345098 580028 346015
rect 579988 345092 580040 345098
rect 579988 345034 580040 345040
rect 580170 322688 580226 322697
rect 580170 322623 580226 322632
rect 580184 321638 580212 322623
rect 580172 321632 580224 321638
rect 580172 321574 580224 321580
rect 580170 310856 580226 310865
rect 580170 310791 580226 310800
rect 580184 310554 580212 310791
rect 580172 310548 580224 310554
rect 580172 310490 580224 310496
rect 579986 275768 580042 275777
rect 579986 275703 580042 275712
rect 580000 274718 580028 275703
rect 579988 274712 580040 274718
rect 579988 274654 580040 274660
rect 580170 263936 580226 263945
rect 580170 263871 580226 263880
rect 580184 263634 580212 263871
rect 580172 263628 580224 263634
rect 580172 263570 580224 263576
rect 580170 252240 580226 252249
rect 580170 252175 580226 252184
rect 580078 228848 580134 228857
rect 580078 228783 580134 228792
rect 580092 227798 580120 228783
rect 580080 227792 580132 227798
rect 580080 227734 580132 227740
rect 579802 217016 579858 217025
rect 579802 216951 579858 216960
rect 579816 216714 579844 216951
rect 579804 216708 579856 216714
rect 579804 216650 579856 216656
rect 580078 205320 580134 205329
rect 580078 205255 580134 205264
rect 505744 202156 505796 202162
rect 505744 202098 505796 202104
rect 504180 201272 504232 201278
rect 504180 201214 504232 201220
rect 504456 201272 504508 201278
rect 504456 201214 504508 201220
rect 504468 186266 504496 201214
rect 579988 200184 580040 200190
rect 579988 200126 580040 200132
rect 504376 186238 504496 186266
rect 504376 183569 504404 186238
rect 504362 183560 504418 183569
rect 504362 183495 504418 183504
rect 504638 183560 504694 183569
rect 504638 183495 504694 183504
rect 504652 173942 504680 183495
rect 580000 181937 580028 200126
rect 579986 181928 580042 181937
rect 579986 181863 580042 181872
rect 504456 173936 504508 173942
rect 504456 173878 504508 173884
rect 504640 173936 504692 173942
rect 504640 173878 504692 173884
rect 504468 166954 504496 173878
rect 504376 166926 504496 166954
rect 504376 164218 504404 166926
rect 504180 164212 504232 164218
rect 504180 164154 504232 164160
rect 504364 164212 504416 164218
rect 504364 164154 504416 164160
rect 504192 154601 504220 164154
rect 504178 154592 504234 154601
rect 504178 154527 504234 154536
rect 504454 154592 504510 154601
rect 504454 154527 504510 154536
rect 442264 151972 442316 151978
rect 442264 151914 442316 151920
rect 440884 150340 440936 150346
rect 440884 150282 440936 150288
rect 439504 148912 439556 148918
rect 439504 148854 439556 148860
rect 438308 142112 438360 142118
rect 438308 142054 438360 142060
rect 437388 140752 437440 140758
rect 437388 140694 437440 140700
rect 437400 140321 437428 140694
rect 437386 140312 437442 140321
rect 437386 140247 437442 140256
rect 437388 137964 437440 137970
rect 437388 137906 437440 137912
rect 437400 137873 437428 137906
rect 437386 137864 437442 137873
rect 437386 137799 437442 137808
rect 504468 136610 504496 154527
rect 437020 136604 437072 136610
rect 437020 136546 437072 136552
rect 504456 136604 504508 136610
rect 504456 136546 504508 136552
rect 437032 136105 437060 136546
rect 437018 136096 437074 136105
rect 437018 136031 437074 136040
rect 437388 133884 437440 133890
rect 437388 133826 437440 133832
rect 437400 133657 437428 133826
rect 437386 133648 437442 133657
rect 437386 133583 437442 133592
rect 436836 132456 436888 132462
rect 436836 132398 436888 132404
rect 436848 132025 436876 132398
rect 436834 132016 436890 132025
rect 436834 131951 436890 131960
rect 580092 129742 580120 205255
rect 580184 132462 580212 252175
rect 580276 144906 580304 533831
rect 580368 200938 580396 545527
rect 580460 500342 580488 557223
rect 580538 510368 580594 510377
rect 580538 510303 580594 510312
rect 580448 500336 580500 500342
rect 580448 500278 580500 500284
rect 580552 500274 580580 510303
rect 580540 500268 580592 500274
rect 580540 500210 580592 500216
rect 580446 439920 580502 439929
rect 580446 439855 580502 439864
rect 580356 200932 580408 200938
rect 580356 200874 580408 200880
rect 580354 170096 580410 170105
rect 580354 170031 580410 170040
rect 580264 144900 580316 144906
rect 580264 144842 580316 144848
rect 580262 134872 580318 134881
rect 580262 134807 580318 134816
rect 580172 132456 580224 132462
rect 580172 132398 580224 132404
rect 437388 129736 437440 129742
rect 437388 129678 437440 129684
rect 580080 129736 580132 129742
rect 580080 129678 580132 129684
rect 437400 129577 437428 129678
rect 437386 129568 437442 129577
rect 437386 129503 437442 129512
rect 436926 124536 436982 124545
rect 436926 124471 436982 124480
rect 436834 122904 436890 122913
rect 436834 122839 436890 122848
rect 436468 120624 436520 120630
rect 436468 120566 436520 120572
rect 436742 120456 436798 120465
rect 436742 120391 436798 120400
rect 436376 80028 436428 80034
rect 436376 79970 436428 79976
rect 436284 35896 436336 35902
rect 436284 35838 436336 35844
rect 436756 17950 436784 120391
rect 436848 64870 436876 122839
rect 436940 111790 436968 124471
rect 580276 120698 580304 134807
rect 580368 120766 580396 170031
rect 580460 140758 580488 439855
rect 580630 404832 580686 404841
rect 580630 404767 580686 404776
rect 580538 393000 580594 393009
rect 580538 392935 580594 392944
rect 580448 140752 580500 140758
rect 580448 140694 580500 140700
rect 580552 137970 580580 392935
rect 580644 200870 580672 404767
rect 580722 369608 580778 369617
rect 580722 369543 580778 369552
rect 580736 201006 580764 369543
rect 580906 357912 580962 357921
rect 580906 357847 580962 357856
rect 580814 299160 580870 299169
rect 580814 299095 580870 299104
rect 580724 201000 580776 201006
rect 580724 200942 580776 200948
rect 580632 200864 580684 200870
rect 580632 200806 580684 200812
rect 580630 158400 580686 158409
rect 580630 158335 580686 158344
rect 580540 137964 580592 137970
rect 580540 137906 580592 137912
rect 580644 128314 580672 158335
rect 580828 133890 580856 299095
rect 580920 200802 580948 357847
rect 580908 200796 580960 200802
rect 580908 200738 580960 200744
rect 580816 133884 580868 133890
rect 580816 133826 580868 133832
rect 580632 128308 580684 128314
rect 580632 128250 580684 128256
rect 580906 123176 580962 123185
rect 580906 123111 580962 123120
rect 580920 120834 580948 123111
rect 580908 120828 580960 120834
rect 580908 120770 580960 120776
rect 580356 120760 580408 120766
rect 580356 120702 580408 120708
rect 580264 120692 580316 120698
rect 580264 120634 580316 120640
rect 493324 118652 493376 118658
rect 493324 118594 493376 118600
rect 478144 118584 478196 118590
rect 478144 118526 478196 118532
rect 475384 118516 475436 118522
rect 475384 118458 475436 118464
rect 474004 118380 474056 118386
rect 474004 118322 474056 118328
rect 443000 118312 443052 118318
rect 443000 118254 443052 118260
rect 439504 117360 439556 117366
rect 439504 117302 439556 117308
rect 436928 111784 436980 111790
rect 436928 111726 436980 111732
rect 436836 64864 436888 64870
rect 436836 64806 436888 64812
rect 436744 17944 436796 17950
rect 436744 17886 436796 17892
rect 437480 10056 437532 10062
rect 437480 9998 437532 10004
rect 434628 9988 434680 9994
rect 434628 9930 434680 9936
rect 433524 7336 433576 7342
rect 433524 7278 433576 7284
rect 433248 4820 433300 4826
rect 433248 4762 433300 4768
rect 431224 3460 431276 3466
rect 431224 3402 431276 3408
rect 432328 3120 432380 3126
rect 432328 3062 432380 3068
rect 432340 480 432368 3062
rect 433536 480 433564 7278
rect 434640 480 434668 9930
rect 437020 8628 437072 8634
rect 437020 8570 437072 8576
rect 435824 7268 435876 7274
rect 435824 7210 435876 7216
rect 435836 480 435864 7210
rect 437032 480 437060 8570
rect 437492 626 437520 9998
rect 439516 3534 439544 117302
rect 441620 10192 441672 10198
rect 441620 10134 441672 10140
rect 440608 8696 440660 8702
rect 440608 8638 440660 8644
rect 439504 3528 439556 3534
rect 439504 3470 439556 3476
rect 439412 3052 439464 3058
rect 439412 2994 439464 3000
rect 437492 598 438164 626
rect 438136 592 438164 598
rect 438136 564 438256 592
rect 438228 480 438256 564
rect 439424 480 439452 2994
rect 440620 480 440648 8638
rect 441632 610 441660 10134
rect 441620 604 441672 610
rect 441620 546 441672 552
rect 441804 604 441856 610
rect 441804 546 441856 552
rect 441816 480 441844 546
rect 443012 480 443040 118254
rect 449900 118244 449952 118250
rect 449900 118186 449952 118192
rect 448520 10260 448572 10266
rect 448520 10202 448572 10208
rect 444380 10124 444432 10130
rect 444380 10066 444432 10072
rect 444196 8764 444248 8770
rect 444196 8706 444248 8712
rect 444208 480 444236 8706
rect 444392 610 444420 10066
rect 447784 8832 447836 8838
rect 447784 8774 447836 8780
rect 446588 3188 446640 3194
rect 446588 3130 446640 3136
rect 444380 604 444432 610
rect 444380 546 444432 552
rect 445392 604 445444 610
rect 445392 546 445444 552
rect 445404 480 445432 546
rect 446600 480 446628 3130
rect 447796 480 447824 8774
rect 448532 610 448560 10202
rect 449912 626 449940 118186
rect 456800 118176 456852 118182
rect 456800 118118 456852 118124
rect 451280 11008 451332 11014
rect 451280 10950 451332 10956
rect 451292 3194 451320 10950
rect 455420 10940 455472 10946
rect 455420 10882 455472 10888
rect 454868 9648 454920 9654
rect 454868 9590 454920 9596
rect 451372 8900 451424 8906
rect 451372 8842 451424 8848
rect 451280 3188 451332 3194
rect 451280 3130 451332 3136
rect 451384 1442 451412 8842
rect 453672 3324 453724 3330
rect 453672 3266 453724 3272
rect 452476 3188 452528 3194
rect 452476 3130 452528 3136
rect 451292 1414 451412 1442
rect 448520 604 448572 610
rect 448520 546 448572 552
rect 448980 604 449032 610
rect 449912 598 450216 626
rect 448980 546 449032 552
rect 448992 480 449020 546
rect 450188 480 450216 598
rect 451292 480 451320 1414
rect 452488 480 452516 3130
rect 453684 480 453712 3266
rect 454880 480 454908 9590
rect 455432 610 455460 10882
rect 456812 610 456840 118118
rect 463700 118108 463752 118114
rect 463700 118050 463752 118056
rect 459652 10872 459704 10878
rect 459652 10814 459704 10820
rect 458456 9580 458508 9586
rect 458456 9522 458508 9528
rect 455420 604 455472 610
rect 455420 546 455472 552
rect 456064 604 456116 610
rect 456064 546 456116 552
rect 456800 604 456852 610
rect 456800 546 456852 552
rect 457260 604 457312 610
rect 457260 546 457312 552
rect 456076 480 456104 546
rect 457272 480 457300 546
rect 458468 480 458496 9522
rect 459664 480 459692 10814
rect 462320 10804 462372 10810
rect 462320 10746 462372 10752
rect 462044 9512 462096 9518
rect 462044 9454 462096 9460
rect 460848 3256 460900 3262
rect 460848 3198 460900 3204
rect 460860 480 460888 3198
rect 462056 480 462084 9454
rect 462332 3482 462360 10746
rect 463712 3482 463740 118050
rect 470600 118040 470652 118046
rect 470600 117982 470652 117988
rect 466460 10736 466512 10742
rect 466460 10678 466512 10684
rect 465632 5704 465684 5710
rect 465632 5646 465684 5652
rect 462332 3454 463280 3482
rect 463712 3454 464476 3482
rect 463252 480 463280 3454
rect 464448 480 464476 3454
rect 465644 480 465672 5646
rect 466472 3482 466500 10678
rect 469220 10668 469272 10674
rect 469220 10610 469272 10616
rect 469128 5636 469180 5642
rect 469128 5578 469180 5584
rect 466472 3454 466868 3482
rect 466840 480 466868 3454
rect 467932 3392 467984 3398
rect 467932 3334 467984 3340
rect 467944 480 467972 3334
rect 469140 480 469168 5578
rect 469232 3482 469260 10610
rect 469232 3454 470364 3482
rect 470336 480 470364 3454
rect 470612 3346 470640 117982
rect 473360 10600 473412 10606
rect 473360 10542 473412 10548
rect 472716 5772 472768 5778
rect 472716 5714 472768 5720
rect 470612 3318 471560 3346
rect 471532 480 471560 3318
rect 472728 480 472756 5714
rect 473372 3346 473400 10542
rect 473372 3318 473952 3346
rect 473924 480 473952 3318
rect 474016 2922 474044 118322
rect 475108 4140 475160 4146
rect 475108 4082 475160 4088
rect 474004 2916 474056 2922
rect 474004 2858 474056 2864
rect 475120 480 475148 4082
rect 475396 2990 475424 118458
rect 477500 117972 477552 117978
rect 477500 117914 477552 117920
rect 476304 5908 476356 5914
rect 476304 5850 476356 5856
rect 475384 2984 475436 2990
rect 475384 2926 475436 2932
rect 476316 480 476344 5850
rect 477512 4146 477540 117914
rect 477592 10532 477644 10538
rect 477592 10474 477644 10480
rect 477500 4140 477552 4146
rect 477500 4082 477552 4088
rect 477604 3482 477632 10474
rect 477512 3454 477632 3482
rect 477512 480 477540 3454
rect 478156 3058 478184 118526
rect 489184 117904 489236 117910
rect 489184 117846 489236 117852
rect 486424 117836 486476 117842
rect 486424 117778 486476 117784
rect 480904 117768 480956 117774
rect 480904 117710 480956 117716
rect 480260 10464 480312 10470
rect 480260 10406 480312 10412
rect 479892 5840 479944 5846
rect 479892 5782 479944 5788
rect 478696 4140 478748 4146
rect 478696 4082 478748 4088
rect 478144 3052 478196 3058
rect 478144 2994 478196 3000
rect 478708 480 478736 4082
rect 479904 480 479932 5782
rect 480272 3618 480300 10406
rect 480916 4146 480944 117710
rect 482284 117700 482336 117706
rect 482284 117642 482336 117648
rect 482296 6882 482324 117642
rect 485780 10396 485832 10402
rect 485780 10338 485832 10344
rect 483480 7404 483532 7410
rect 483480 7346 483532 7352
rect 482204 6854 482324 6882
rect 480904 4140 480956 4146
rect 480904 4082 480956 4088
rect 481272 4140 481324 4146
rect 481272 4082 481324 4088
rect 480272 3590 481128 3618
rect 481100 480 481128 3590
rect 481284 3126 481312 4082
rect 482204 3262 482232 6854
rect 482284 4072 482336 4078
rect 482284 4014 482336 4020
rect 482192 3256 482244 3262
rect 482192 3198 482244 3204
rect 481272 3120 481324 3126
rect 481272 3062 481324 3068
rect 482296 480 482324 4014
rect 483492 480 483520 7346
rect 484584 6044 484636 6050
rect 484584 5986 484636 5992
rect 484596 480 484624 5986
rect 485792 480 485820 10338
rect 486436 3194 486464 117778
rect 488540 12232 488592 12238
rect 488540 12174 488592 12180
rect 486976 7472 487028 7478
rect 486976 7414 487028 7420
rect 486424 3188 486476 3194
rect 486424 3130 486476 3136
rect 486988 480 487016 7414
rect 488172 5976 488224 5982
rect 488172 5918 488224 5924
rect 488184 480 488212 5918
rect 488552 3618 488580 12174
rect 489196 4146 489224 117846
rect 492680 12164 492732 12170
rect 492680 12106 492732 12112
rect 490564 7540 490616 7546
rect 490564 7482 490616 7488
rect 489184 4140 489236 4146
rect 489184 4082 489236 4088
rect 489552 4140 489604 4146
rect 489552 4082 489604 4088
rect 488552 3590 489408 3618
rect 489380 480 489408 3590
rect 489564 3330 489592 4082
rect 489552 3324 489604 3330
rect 489552 3266 489604 3272
rect 490576 480 490604 7482
rect 491760 6112 491812 6118
rect 491760 6054 491812 6060
rect 491772 480 491800 6054
rect 492692 3482 492720 12106
rect 492692 3454 492996 3482
rect 492968 480 492996 3454
rect 493336 3398 493364 118594
rect 500224 118448 500276 118454
rect 500224 118390 500276 118396
rect 496084 117632 496136 117638
rect 496084 117574 496136 117580
rect 495440 12096 495492 12102
rect 495440 12038 495492 12044
rect 494152 8288 494204 8294
rect 494152 8230 494204 8236
rect 493324 3392 493376 3398
rect 493324 3334 493376 3340
rect 494164 480 494192 8230
rect 495348 6860 495400 6866
rect 495348 6802 495400 6808
rect 495360 480 495388 6802
rect 495452 3618 495480 12038
rect 496096 4146 496124 117574
rect 499580 12028 499632 12034
rect 499580 11970 499632 11976
rect 497740 8220 497792 8226
rect 497740 8162 497792 8168
rect 496084 4140 496136 4146
rect 496084 4082 496136 4088
rect 495452 3590 496584 3618
rect 496556 480 496584 3590
rect 497752 480 497780 8162
rect 498936 6792 498988 6798
rect 498936 6734 498988 6740
rect 498948 480 498976 6734
rect 499592 610 499620 11970
rect 500236 4078 500264 118390
rect 579804 111784 579856 111790
rect 579804 111726 579856 111732
rect 579816 111489 579844 111726
rect 579802 111480 579858 111489
rect 579802 111415 579858 111424
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 580172 77240 580224 77246
rect 580172 77182 580224 77188
rect 580184 76265 580212 77182
rect 580170 76256 580226 76265
rect 580170 76191 580226 76200
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 580172 30320 580224 30326
rect 580172 30262 580224 30268
rect 580184 29345 580212 30262
rect 580170 29336 580226 29345
rect 580170 29271 580226 29280
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 502340 11960 502392 11966
rect 502340 11902 502392 11908
rect 501236 9444 501288 9450
rect 501236 9386 501288 9392
rect 500224 4072 500276 4078
rect 500224 4014 500276 4020
rect 499580 604 499632 610
rect 499580 546 499632 552
rect 500132 604 500184 610
rect 500132 546 500184 552
rect 500144 480 500172 546
rect 501248 480 501276 9386
rect 502352 2854 502380 11902
rect 506480 11892 506532 11898
rect 506480 11834 506532 11840
rect 504824 9376 504876 9382
rect 504824 9318 504876 9324
rect 502432 6724 502484 6730
rect 502432 6666 502484 6672
rect 502340 2848 502392 2854
rect 502340 2790 502392 2796
rect 502444 480 502472 6666
rect 503548 4146 503852 4162
rect 503536 4140 503864 4146
rect 503588 4134 503812 4140
rect 503536 4082 503588 4088
rect 503812 4082 503864 4088
rect 503628 2848 503680 2854
rect 503628 2790 503680 2796
rect 503640 480 503668 2790
rect 504836 480 504864 9318
rect 506020 6656 506072 6662
rect 506020 6598 506072 6604
rect 506032 480 506060 6598
rect 506492 610 506520 11834
rect 510620 11824 510672 11830
rect 510620 11766 510672 11772
rect 508412 9308 508464 9314
rect 508412 9250 508464 9256
rect 506480 604 506532 610
rect 506480 546 506532 552
rect 507216 604 507268 610
rect 507216 546 507268 552
rect 507228 480 507256 546
rect 508424 480 508452 9250
rect 509608 6588 509660 6594
rect 509608 6530 509660 6536
rect 509620 480 509648 6530
rect 510632 610 510660 11766
rect 513380 11756 513432 11762
rect 513380 11698 513432 11704
rect 512000 9240 512052 9246
rect 512000 9182 512052 9188
rect 510620 604 510672 610
rect 510620 546 510672 552
rect 510804 604 510856 610
rect 510804 546 510856 552
rect 510816 480 510844 546
rect 512012 480 512040 9182
rect 513196 6520 513248 6526
rect 513196 6462 513248 6468
rect 513208 480 513236 6462
rect 513392 610 513420 11698
rect 581092 10328 581144 10334
rect 581092 10270 581144 10276
rect 566740 9172 566792 9178
rect 566740 9114 566792 9120
rect 534540 8152 534592 8158
rect 534540 8094 534592 8100
rect 516784 6452 516836 6458
rect 516784 6394 516836 6400
rect 515588 4276 515640 4282
rect 515588 4218 515640 4224
rect 513380 604 513432 610
rect 513380 546 513432 552
rect 514392 604 514444 610
rect 514392 546 514444 552
rect 514404 480 514432 546
rect 515600 480 515628 4218
rect 516796 480 516824 6394
rect 520280 6384 520332 6390
rect 520280 6326 520332 6332
rect 519084 4344 519136 4350
rect 519084 4286 519136 4292
rect 517888 2916 517940 2922
rect 517888 2858 517940 2864
rect 517900 480 517928 2858
rect 519096 480 519124 4286
rect 520292 480 520320 6326
rect 523868 6316 523920 6322
rect 523868 6258 523920 6264
rect 522672 4412 522724 4418
rect 522672 4354 522724 4360
rect 521476 4004 521528 4010
rect 521476 3946 521528 3952
rect 521488 480 521516 3946
rect 522684 480 522712 4354
rect 523880 480 523908 6258
rect 531044 6248 531096 6254
rect 531044 6190 531096 6196
rect 527456 6180 527508 6186
rect 527456 6122 527508 6128
rect 526260 4480 526312 4486
rect 526260 4422 526312 4428
rect 525064 2984 525116 2990
rect 525064 2926 525116 2932
rect 525076 480 525104 2926
rect 526272 480 526300 4422
rect 527468 480 527496 6122
rect 529848 4548 529900 4554
rect 529848 4490 529900 4496
rect 528652 3936 528704 3942
rect 528652 3878 528704 3884
rect 528664 480 528692 3878
rect 529860 480 529888 4490
rect 531056 480 531084 6190
rect 533436 4616 533488 4622
rect 533436 4558 533488 4564
rect 532240 3052 532292 3058
rect 532240 2994 532292 3000
rect 532252 480 532280 2994
rect 533448 480 533476 4558
rect 534552 480 534580 8094
rect 538128 8084 538180 8090
rect 538128 8026 538180 8032
rect 536932 4684 536984 4690
rect 536932 4626 536984 4632
rect 535736 3868 535788 3874
rect 535736 3810 535788 3816
rect 535748 480 535776 3810
rect 536944 480 536972 4626
rect 538140 480 538168 8026
rect 541716 8016 541768 8022
rect 541716 7958 541768 7964
rect 540520 4752 540572 4758
rect 540520 4694 540572 4700
rect 539324 3120 539376 3126
rect 539324 3062 539376 3068
rect 539336 480 539364 3062
rect 540532 480 540560 4694
rect 541728 480 541756 7958
rect 545304 7948 545356 7954
rect 545304 7890 545356 7896
rect 544108 5500 544160 5506
rect 544108 5442 544160 5448
rect 542912 3800 542964 3806
rect 542912 3742 542964 3748
rect 542924 480 542952 3742
rect 544120 480 544148 5442
rect 545316 480 545344 7890
rect 548892 7880 548944 7886
rect 548892 7822 548944 7828
rect 547696 5432 547748 5438
rect 547696 5374 547748 5380
rect 546500 3256 546552 3262
rect 546500 3198 546552 3204
rect 546512 480 546540 3198
rect 547708 480 547736 5374
rect 548904 480 548932 7822
rect 552388 7812 552440 7818
rect 552388 7754 552440 7760
rect 551192 5364 551244 5370
rect 551192 5306 551244 5312
rect 550088 3188 550140 3194
rect 550088 3130 550140 3136
rect 550100 480 550128 3130
rect 551204 480 551232 5306
rect 552400 480 552428 7754
rect 555976 7744 556028 7750
rect 555976 7686 556028 7692
rect 554780 5296 554832 5302
rect 554780 5238 554832 5244
rect 553584 3732 553636 3738
rect 553584 3674 553636 3680
rect 553596 480 553624 3674
rect 554792 480 554820 5238
rect 555988 480 556016 7686
rect 559564 7676 559616 7682
rect 559564 7618 559616 7624
rect 558368 5228 558420 5234
rect 558368 5170 558420 5176
rect 557172 3324 557224 3330
rect 557172 3266 557224 3272
rect 557184 480 557212 3266
rect 558380 480 558408 5170
rect 559576 480 559604 7618
rect 563152 7608 563204 7614
rect 563152 7550 563204 7556
rect 561956 5092 562008 5098
rect 561956 5034 562008 5040
rect 560760 3664 560812 3670
rect 560760 3606 560812 3612
rect 560772 480 560800 3606
rect 561968 480 561996 5034
rect 563164 480 563192 7550
rect 565544 5160 565596 5166
rect 565544 5102 565596 5108
rect 564348 3392 564400 3398
rect 564348 3334 564400 3340
rect 564360 480 564388 3334
rect 565556 480 565584 5102
rect 566752 480 566780 9114
rect 573824 9104 573876 9110
rect 573824 9046 573876 9052
rect 570236 9036 570288 9042
rect 570236 8978 570288 8984
rect 569040 5024 569092 5030
rect 569040 4966 569092 4972
rect 567844 3596 567896 3602
rect 567844 3538 567896 3544
rect 567856 480 567884 3538
rect 569052 480 569080 4966
rect 570248 480 570276 8978
rect 572628 4956 572680 4962
rect 572628 4898 572680 4904
rect 571432 4140 571484 4146
rect 571432 4082 571484 4088
rect 571444 480 571472 4082
rect 572640 480 572668 4898
rect 573836 480 573864 9046
rect 577412 8968 577464 8974
rect 577412 8910 577464 8916
rect 576216 4888 576268 4894
rect 576216 4830 576268 4836
rect 575020 3460 575072 3466
rect 575020 3402 575072 3408
rect 575032 480 575060 3402
rect 576228 480 576256 4830
rect 577424 480 577452 8910
rect 579804 4820 579856 4826
rect 579804 4762 579856 4768
rect 578608 4072 578660 4078
rect 578608 4014 578660 4020
rect 578620 480 578648 4014
rect 579816 480 579844 4762
rect 581104 626 581132 10270
rect 582196 3528 582248 3534
rect 582196 3470 582248 3476
rect 581012 598 581132 626
rect 581012 480 581040 598
rect 582208 480 582236 3470
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3790 682216 3846 682272
rect 3422 667936 3478 667992
rect 3054 624824 3110 624880
rect 3146 481092 3202 481128
rect 3146 481072 3148 481092
rect 3148 481072 3200 481092
rect 3200 481072 3202 481092
rect 3238 452376 3294 452432
rect 3330 437960 3386 438016
rect 3238 423680 3294 423736
rect 3054 394984 3110 395040
rect 2962 366172 3018 366208
rect 2962 366152 2964 366172
rect 2964 366152 3016 366172
rect 3016 366152 3018 366172
rect 2962 337456 3018 337512
rect 2962 323040 3018 323096
rect 2962 308760 3018 308816
rect 2962 294344 3018 294400
rect 2962 280064 3018 280120
rect 2870 265648 2926 265704
rect 2870 251252 2926 251288
rect 2870 251232 2872 251252
rect 2872 251232 2924 251252
rect 2924 251232 2926 251252
rect 2870 236952 2926 237008
rect 2778 222556 2834 222592
rect 2778 222536 2780 222556
rect 2780 222536 2832 222556
rect 2832 222536 2834 222556
rect 2778 165008 2834 165064
rect 3146 380568 3202 380624
rect 3054 208120 3110 208176
rect 3054 193840 3110 193896
rect 3514 653520 3570 653576
rect 3606 610408 3662 610464
rect 3698 595992 3754 596048
rect 3882 567296 3938 567352
rect 3790 553016 3846 553072
rect 3698 179460 3700 179480
rect 3700 179460 3752 179480
rect 3752 179460 3754 179480
rect 3698 179424 3754 179460
rect 3974 538600 4030 538656
rect 4066 509904 4122 509960
rect 3974 495488 4030 495544
rect 2778 136348 2780 136368
rect 2780 136348 2832 136368
rect 2832 136348 2834 136368
rect 2778 136312 2834 136348
rect 3238 122032 3294 122088
rect 3238 107616 3294 107672
rect 3422 93200 3478 93256
rect 3146 78920 3202 78976
rect 3330 64504 3386 64560
rect 3422 35844 3424 35864
rect 3424 35844 3476 35864
rect 3476 35844 3478 35864
rect 3422 35808 3478 35844
rect 2778 21428 2780 21448
rect 2780 21428 2832 21448
rect 2832 21428 2834 21448
rect 2778 21392 2834 21428
rect 8114 531256 8170 531312
rect 8390 531256 8446 531312
rect 8114 511944 8170 512000
rect 8390 511944 8446 512000
rect 7930 473320 7986 473376
rect 8114 473320 8170 473376
rect 4158 150728 4214 150784
rect 4066 50088 4122 50144
rect 8022 193160 8078 193216
rect 8298 193160 8354 193216
rect 9678 188944 9734 189000
rect 6918 153076 6920 153096
rect 6920 153076 6972 153096
rect 6972 153076 6974 153096
rect 6918 153040 6974 153076
rect 3882 7112 3938 7168
rect 19246 188944 19302 189000
rect 16486 153040 16542 153096
rect 70122 370232 70178 370288
rect 70122 355544 70178 355600
rect 71502 385192 71558 385248
rect 70306 377848 70362 377904
rect 71042 377848 71098 377904
rect 70306 370232 70362 370288
rect 70214 348200 70270 348256
rect 70122 341400 70178 341456
rect 67638 188828 67694 188864
rect 67638 188808 67640 188828
rect 67640 188808 67692 188828
rect 67692 188808 67694 188828
rect 64878 148724 64880 148744
rect 64880 148724 64932 148744
rect 64932 148724 64934 148744
rect 64878 148688 64934 148724
rect 70398 148688 70454 148744
rect 71594 362888 71650 362944
rect 71594 348200 71650 348256
rect 72330 392944 72386 393000
rect 84106 545808 84162 545864
rect 84014 541456 84070 541512
rect 83922 537104 83978 537160
rect 83830 528672 83886 528728
rect 82818 524864 82874 524920
rect 85302 533024 85358 533080
rect 85394 525544 85450 525600
rect 86406 549908 86462 549944
rect 86406 549888 86408 549908
rect 86408 549888 86460 549908
rect 86460 549888 86462 549908
rect 85578 537716 85634 537772
rect 96618 395836 96620 395856
rect 96620 395836 96672 395856
rect 96672 395836 96674 395856
rect 96618 395800 96674 395836
rect 99286 395800 99342 395856
rect 116030 578312 116086 578368
rect 118054 546488 118110 546544
rect 117778 537376 117834 537432
rect 117778 533296 117834 533352
rect 117962 529624 118018 529680
rect 117318 521056 117374 521112
rect 118606 542428 118662 542464
rect 118606 542408 118608 542428
rect 118608 542408 118660 542428
rect 118660 542408 118662 542428
rect 118606 525136 118662 525192
rect 125506 578348 125508 578368
rect 125508 578348 125560 578368
rect 125560 578348 125562 578368
rect 125506 578312 125562 578348
rect 77206 188808 77262 188864
rect 86958 188828 87014 188864
rect 86958 188808 86960 188828
rect 86960 188808 87012 188828
rect 87012 188808 87014 188828
rect 96342 188808 96398 188864
rect 84198 148844 84254 148880
rect 84198 148824 84200 148844
rect 84200 148824 84252 148844
rect 84252 148824 84254 148844
rect 93582 148824 93638 148880
rect 97998 117816 98054 117872
rect 99286 117816 99342 117872
rect 115938 188828 115994 188864
rect 115938 188808 115940 188828
rect 115940 188808 115992 188828
rect 115992 188808 115994 188828
rect 122654 212472 122710 212528
rect 122838 212472 122894 212528
rect 122654 202816 122710 202872
rect 122930 202816 122986 202872
rect 125506 188808 125562 188864
rect 117226 117680 117282 117736
rect 115938 117272 115994 117328
rect 117226 117272 117282 117328
rect 125782 118360 125838 118416
rect 128082 251232 128138 251288
rect 126978 118632 127034 118688
rect 126242 118224 126298 118280
rect 128542 387912 128598 387968
rect 128450 373224 128506 373280
rect 128450 372680 128506 372736
rect 128910 365880 128966 365936
rect 128634 358672 128690 358728
rect 128818 343576 128874 343632
rect 128358 335280 128414 335336
rect 128542 335280 128598 335336
rect 128450 251232 128506 251288
rect 128450 212472 128506 212528
rect 128634 212472 128690 212528
rect 128358 193160 128414 193216
rect 128542 193160 128598 193216
rect 128358 164192 128414 164248
rect 128542 164192 128598 164248
rect 128542 154808 128598 154864
rect 128542 154536 128598 154592
rect 128818 125588 128874 125624
rect 128818 125568 128820 125588
rect 128820 125568 128872 125588
rect 128872 125568 128874 125588
rect 129094 387912 129150 387968
rect 129186 380568 129242 380624
rect 129002 143520 129058 143576
rect 129094 125588 129150 125624
rect 129278 372680 129334 372736
rect 129094 125568 129096 125588
rect 129096 125568 129148 125588
rect 129148 125568 129150 125588
rect 129738 350920 129794 350976
rect 129186 118088 129242 118144
rect 128818 115912 128874 115968
rect 129002 115932 129058 115968
rect 129002 115912 129004 115932
rect 129004 115912 129056 115932
rect 129056 115912 129058 115932
rect 128726 106256 128782 106312
rect 128910 106256 128966 106312
rect 128910 67768 128966 67824
rect 129094 67632 129150 67688
rect 130382 117952 130438 118008
rect 130658 171944 130714 172000
rect 130750 170856 130806 170912
rect 130566 169768 130622 169824
rect 130934 172896 130990 172952
rect 130934 156576 130990 156632
rect 131210 199280 131266 199336
rect 131210 198192 131266 198248
rect 131302 197104 131358 197160
rect 131210 196036 131266 196072
rect 131210 196016 131212 196036
rect 131212 196016 131264 196036
rect 131264 196016 131266 196036
rect 131210 195064 131266 195120
rect 131210 193976 131266 194032
rect 131210 192888 131266 192944
rect 131210 191936 131266 191992
rect 131210 190848 131266 190904
rect 131210 189760 131266 189816
rect 131210 188672 131266 188728
rect 131210 187720 131266 187776
rect 131210 186632 131266 186688
rect 131210 185544 131266 185600
rect 131210 184456 131266 184512
rect 131210 183524 131266 183560
rect 131210 183504 131212 183524
rect 131212 183504 131264 183524
rect 131264 183504 131266 183524
rect 131210 175072 131266 175128
rect 131210 159296 131266 159352
rect 131210 156168 131266 156224
rect 131210 155080 131266 155136
rect 131210 153992 131266 154048
rect 131210 152904 131266 152960
rect 131210 151952 131266 152008
rect 131210 150864 131266 150920
rect 131210 149776 131266 149832
rect 131210 148688 131266 148744
rect 131210 148280 131266 148336
rect 131118 145560 131174 145616
rect 131118 144472 131174 144528
rect 131118 138216 131174 138272
rect 131302 131960 131358 132016
rect 131394 128696 131450 128752
rect 131578 165552 131634 165608
rect 131578 158208 131634 158264
rect 131486 127744 131542 127800
rect 132038 180376 132094 180432
rect 132038 173984 132094 174040
rect 132038 166640 132094 166696
rect 132038 160384 132094 160440
rect 131946 134000 132002 134056
rect 131854 130872 131910 130928
rect 131762 126656 131818 126712
rect 131670 125568 131726 125624
rect 132222 147736 132278 147792
rect 132406 167728 132462 167784
rect 132406 162424 132462 162480
rect 132314 147464 132370 147520
rect 132222 146648 132278 146704
rect 132314 142432 132370 142488
rect 132222 140392 132278 140448
rect 132130 135088 132186 135144
rect 132314 121352 132370 121408
rect 132130 120400 132186 120456
rect 132866 241440 132922 241496
rect 132682 164464 132738 164520
rect 132498 136176 132554 136232
rect 132866 196016 132922 196072
rect 132866 195880 132922 195936
rect 132866 182416 132922 182472
rect 132866 182280 132922 182336
rect 132866 178200 132922 178256
rect 133234 185408 133290 185464
rect 133050 184864 133106 184920
rect 132958 168680 133014 168736
rect 132958 164192 133014 164248
rect 132958 154672 133014 154728
rect 132958 154536 133014 154592
rect 132774 124480 132830 124536
rect 132958 118496 133014 118552
rect 133234 181328 133290 181384
rect 133326 179288 133382 179344
rect 133510 241440 133566 241496
rect 133418 177112 133474 177168
rect 133234 176160 133290 176216
rect 133142 164192 133198 164248
rect 133510 163512 133566 163568
rect 133510 161336 133566 161392
rect 133234 118108 133290 118144
rect 133234 118088 133236 118108
rect 133236 118088 133288 118108
rect 133288 118088 133290 118108
rect 133050 117544 133106 117600
rect 133602 139304 133658 139360
rect 133694 137128 133750 137184
rect 133878 141344 133934 141400
rect 133970 133456 134026 133512
rect 134338 341400 134394 341456
rect 134338 200096 134394 200152
rect 154578 340468 154634 340504
rect 154578 340448 154580 340468
rect 154580 340448 154632 340468
rect 154632 340448 154634 340468
rect 157338 340448 157394 340504
rect 185582 341400 185638 341456
rect 193218 340348 193220 340368
rect 193220 340348 193272 340368
rect 193272 340348 193274 340368
rect 193218 340312 193274 340348
rect 195702 202680 195758 202736
rect 195794 202544 195850 202600
rect 198646 556688 198702 556744
rect 198554 552064 198610 552120
rect 198462 543768 198518 543824
rect 198370 538464 198426 538520
rect 198278 524592 198334 524648
rect 198186 399608 198242 399664
rect 198094 391176 198150 391232
rect 198002 387096 198058 387152
rect 197910 378664 197966 378720
rect 197818 370232 197874 370288
rect 197726 361800 197782 361856
rect 197634 357448 197690 357504
rect 197542 353368 197598 353424
rect 197450 349016 197506 349072
rect 197266 202816 197322 202872
rect 197174 202408 197230 202464
rect 197082 202272 197138 202328
rect 222198 556144 222254 556200
rect 198922 547848 198978 547904
rect 198738 534112 198794 534168
rect 198646 202000 198702 202056
rect 198830 529216 198886 529272
rect 219438 528944 219494 529000
rect 199014 403688 199070 403744
rect 199106 395256 199162 395312
rect 199198 382744 199254 382800
rect 199290 374312 199346 374368
rect 199014 202136 199070 202192
rect 199382 365880 199438 365936
rect 199474 344936 199530 344992
rect 219530 524456 219586 524512
rect 222290 552064 222346 552120
rect 222382 546896 222438 546952
rect 222474 542544 222530 542600
rect 222566 538328 222622 538384
rect 222658 533296 222714 533352
rect 265990 415384 266046 415440
rect 266174 415384 266230 415440
rect 240138 340484 240140 340504
rect 240140 340484 240192 340504
rect 240192 340484 240194 340504
rect 240138 340448 240194 340484
rect 249706 340468 249762 340504
rect 249706 340448 249708 340468
rect 249708 340448 249760 340468
rect 249760 340448 249762 340468
rect 259458 340468 259514 340504
rect 259458 340448 259460 340468
rect 259460 340448 259512 340468
rect 259512 340448 259514 340468
rect 202786 340312 202842 340368
rect 230478 340348 230480 340368
rect 230480 340348 230532 340368
rect 230532 340348 230534 340368
rect 230478 340312 230534 340348
rect 240046 340312 240102 340368
rect 213458 202000 213514 202056
rect 220358 202816 220414 202872
rect 223854 202680 223910 202736
rect 226338 202544 226394 202600
rect 228638 202408 228694 202464
rect 233422 202272 233478 202328
rect 252650 202444 252652 202464
rect 252652 202444 252704 202464
rect 252704 202444 252706 202464
rect 252650 202408 252706 202444
rect 253478 202308 253480 202328
rect 253480 202308 253532 202328
rect 253532 202308 253534 202328
rect 253478 202272 253534 202308
rect 258170 326984 258226 327040
rect 258354 326984 258410 327040
rect 255594 309168 255650 309224
rect 255870 309168 255926 309224
rect 258354 309168 258410 309224
rect 258630 309168 258686 309224
rect 257986 241440 258042 241496
rect 258170 241440 258226 241496
rect 253938 202272 253994 202328
rect 254122 202444 254124 202464
rect 254124 202444 254176 202464
rect 254176 202444 254178 202464
rect 254122 202408 254178 202444
rect 258538 202292 258594 202328
rect 258538 202272 258540 202292
rect 258540 202272 258592 202292
rect 258592 202272 258594 202292
rect 259458 202272 259514 202328
rect 261942 202136 261998 202192
rect 266818 399608 266874 399664
rect 266910 382744 266966 382800
rect 267094 357448 267150 357504
rect 267186 349016 267242 349072
rect 267738 403688 267794 403744
rect 267830 395256 267886 395312
rect 267922 391176 267978 391232
rect 268014 386824 268070 386880
rect 268106 378392 268162 378448
rect 268198 374312 268254 374368
rect 268290 369960 268346 370016
rect 268382 365880 268438 365936
rect 268474 361528 268530 361584
rect 268566 353368 268622 353424
rect 268658 344936 268714 344992
rect 268934 340448 268990 340504
rect 269118 340468 269174 340504
rect 269118 340448 269120 340468
rect 269120 340448 269172 340468
rect 269172 340448 269174 340468
rect 271786 563080 271842 563136
rect 271694 562944 271750 563000
rect 271510 560224 271566 560280
rect 271694 560224 271750 560280
rect 271694 540912 271750 540968
rect 271970 540912 272026 540968
rect 271602 502324 271604 502344
rect 271604 502324 271656 502344
rect 271656 502324 271658 502344
rect 271602 502288 271658 502324
rect 271786 492632 271842 492688
rect 271786 419464 271842 419520
rect 271970 419464 272026 419520
rect 271602 389156 271658 389192
rect 271602 389136 271604 389156
rect 271604 389136 271656 389156
rect 271656 389136 271658 389156
rect 271786 389136 271842 389192
rect 271970 294072 272026 294128
rect 271786 293936 271842 293992
rect 271970 274760 272026 274816
rect 271786 274624 271842 274680
rect 271602 255312 271658 255368
rect 271786 255312 271842 255368
rect 273258 340468 273314 340504
rect 273258 340448 273260 340468
rect 273260 340448 273312 340468
rect 273312 340448 273314 340468
rect 281262 521872 281318 521928
rect 281354 521634 281410 521690
rect 277306 202136 277362 202192
rect 281078 492632 281134 492688
rect 281262 492632 281318 492688
rect 281078 454008 281134 454064
rect 281262 454008 281318 454064
rect 281078 434696 281134 434752
rect 281262 434696 281318 434752
rect 281630 396072 281686 396128
rect 281630 395936 281686 395992
rect 281170 260752 281226 260808
rect 281078 251096 281134 251152
rect 289818 578876 289874 578912
rect 289818 578856 289820 578876
rect 289820 578856 289872 578876
rect 289872 578856 289874 578876
rect 296718 575728 296774 575784
rect 297362 572872 297418 572928
rect 296718 570016 296774 570072
rect 296442 566072 296498 566128
rect 296718 563216 296774 563272
rect 297270 541048 297326 541104
rect 296534 531528 296590 531584
rect 296718 509496 296774 509552
rect 296718 506524 296774 506560
rect 296718 506504 296720 506524
rect 296720 506504 296772 506524
rect 296772 506504 296774 506524
rect 297914 560360 297970 560416
rect 297822 556824 297878 556880
rect 297822 553560 297878 553616
rect 297730 550704 297786 550760
rect 297638 538328 297694 538384
rect 297638 534792 297694 534848
rect 297362 528536 297418 528592
rect 297454 525816 297510 525872
rect 297546 522008 297602 522064
rect 297454 519016 297510 519072
rect 297454 516180 297510 516216
rect 297454 516160 297456 516180
rect 297456 516160 297508 516180
rect 297508 516160 297510 516180
rect 297454 513440 297510 513496
rect 297362 503784 297418 503840
rect 299110 547848 299166 547904
rect 299018 544040 299074 544096
rect 299386 578856 299442 578912
rect 305182 579300 305184 579320
rect 305184 579300 305236 579320
rect 305236 579300 305238 579320
rect 305182 579264 305238 579300
rect 315854 579300 315856 579320
rect 315856 579300 315908 579320
rect 315908 579300 315910 579320
rect 315854 579264 315910 579300
rect 301870 473320 301926 473376
rect 302054 473320 302110 473376
rect 302238 202564 302294 202600
rect 302238 202544 302240 202564
rect 302240 202544 302292 202564
rect 302292 202544 302294 202564
rect 307022 483112 307078 483168
rect 307022 482976 307078 483032
rect 307022 463800 307078 463856
rect 307022 463684 307078 463720
rect 307022 463664 307024 463684
rect 307024 463664 307076 463684
rect 307076 463664 307078 463684
rect 306838 454008 306894 454064
rect 307022 454008 307078 454064
rect 304262 202000 304318 202056
rect 307206 202580 307208 202600
rect 307208 202580 307260 202600
rect 307260 202580 307262 202600
rect 307206 202544 307262 202580
rect 308862 251368 308918 251424
rect 308862 251232 308918 251288
rect 307298 202000 307354 202056
rect 377402 572056 377458 572112
rect 378138 569676 378194 569732
rect 377678 519152 377734 519208
rect 378230 566412 378286 566468
rect 378322 563420 378378 563476
rect 378414 559544 378470 559600
rect 378598 556552 378654 556608
rect 378506 521736 378562 521792
rect 378690 550704 378746 550760
rect 378874 547032 378930 547088
rect 380530 575456 380586 575512
rect 379518 553424 379574 553480
rect 379610 543768 379666 543824
rect 380346 541048 380402 541104
rect 379702 537512 379758 537568
rect 379794 534520 379850 534576
rect 379886 531392 379942 531448
rect 379978 525000 380034 525056
rect 378414 202136 378470 202192
rect 380070 515480 380126 515536
rect 380162 512488 380218 512544
rect 380254 509496 380310 509552
rect 380438 528672 380494 528728
rect 380346 506504 380402 506560
rect 380714 502968 380770 503024
rect 380898 381384 380954 381440
rect 380898 377168 380954 377224
rect 380898 374060 380954 374096
rect 380898 374040 380900 374060
rect 380900 374040 380952 374060
rect 380952 374040 380954 374060
rect 380898 370368 380954 370424
rect 381542 367376 381598 367432
rect 380898 363568 380954 363624
rect 380898 353504 380954 353560
rect 381634 360304 381690 360360
rect 381726 356768 381782 356824
rect 416870 380840 416926 380896
rect 417422 376896 417478 376952
rect 416778 374584 416834 374640
rect 416870 370096 416926 370152
rect 416962 367104 417018 367160
rect 417054 363296 417110 363352
rect 417146 360168 417202 360224
rect 417238 356496 417294 356552
rect 417330 353368 417386 353424
rect 434258 173848 434314 173904
rect 434994 190168 435050 190224
rect 434902 188808 434958 188864
rect 434810 186224 434866 186280
rect 434718 184592 434774 184648
rect 434534 171944 434590 172000
rect 434442 169632 434498 169688
rect 434350 167728 434406 167784
rect 434166 165552 434222 165608
rect 434074 163512 434130 163568
rect 436374 196152 436430 196208
rect 436282 193024 436338 193080
rect 436190 180240 436246 180296
rect 436098 161200 436154 161256
rect 433982 159296 434038 159352
rect 433890 157256 433946 157312
rect 436098 155080 436154 155136
rect 436190 148860 436192 148880
rect 436192 148860 436244 148880
rect 436244 148860 436246 148880
rect 436190 148824 436246 148860
rect 436098 146260 436154 146296
rect 436098 146240 436100 146260
rect 436100 146240 436152 146260
rect 436152 146240 436154 146260
rect 436098 142060 436100 142080
rect 436100 142060 436152 142080
rect 436152 142060 436154 142080
rect 436098 142024 436154 142060
rect 134062 130328 134118 130384
rect 436098 127744 436154 127800
rect 133970 122984 134026 123040
rect 134062 121896 134118 121952
rect 140778 118496 140834 118552
rect 140870 106392 140926 106448
rect 140778 106276 140834 106312
rect 140778 106256 140780 106276
rect 140780 106256 140832 106276
rect 140832 106256 140834 106276
rect 140778 60832 140834 60888
rect 140778 55256 140834 55312
rect 140870 41384 140926 41440
rect 140778 41248 140834 41304
rect 145102 106256 145158 106312
rect 145286 106256 145342 106312
rect 144826 75792 144882 75848
rect 145010 75792 145066 75848
rect 145102 66136 145158 66192
rect 145194 66000 145250 66056
rect 143722 44104 143778 44160
rect 143998 44104 144054 44160
rect 146482 117952 146538 118008
rect 146850 117952 146906 118008
rect 148046 104896 148102 104952
rect 148230 104896 148286 104952
rect 151818 118632 151874 118688
rect 152186 115912 152242 115968
rect 152462 115912 152518 115968
rect 164606 29144 164662 29200
rect 164514 29008 164570 29064
rect 171138 117172 171140 117192
rect 171140 117172 171192 117192
rect 171192 117172 171194 117192
rect 171138 117136 171194 117172
rect 174266 9560 174322 9616
rect 180706 117136 180762 117192
rect 182178 118088 182234 118144
rect 181074 9560 181130 9616
rect 183374 37168 183430 37224
rect 183650 37168 183706 37224
rect 183926 9832 183982 9888
rect 183650 9696 183706 9752
rect 184938 117816 184994 117872
rect 189078 29008 189134 29064
rect 189354 28872 189410 28928
rect 193954 117680 194010 117736
rect 195978 118224 196034 118280
rect 197634 118360 197690 118416
rect 203062 115912 203118 115968
rect 203706 115912 203762 115968
rect 204534 115912 204590 115968
rect 204902 115912 204958 115968
rect 204626 86944 204682 87000
rect 204810 86944 204866 87000
rect 209962 86944 210018 87000
rect 210146 86944 210202 87000
rect 215942 115912 215998 115968
rect 216126 115912 216182 115968
rect 217046 115912 217102 115968
rect 217414 115912 217470 115968
rect 218242 104760 218298 104816
rect 218426 104624 218482 104680
rect 220174 115912 220230 115968
rect 220358 115912 220414 115968
rect 221462 115912 221518 115968
rect 221646 115912 221702 115968
rect 221094 66272 221150 66328
rect 221278 66272 221334 66328
rect 227994 115912 228050 115968
rect 228270 115912 228326 115968
rect 227810 28872 227866 28928
rect 227994 28872 228050 28928
rect 233422 80144 233478 80200
rect 233238 79872 233294 79928
rect 238942 106256 238998 106312
rect 239126 106256 239182 106312
rect 244278 75792 244334 75848
rect 244646 75792 244702 75848
rect 246946 106392 247002 106448
rect 246946 106256 247002 106312
rect 246946 9832 247002 9888
rect 246762 9696 246818 9752
rect 274454 86944 274510 87000
rect 274914 96736 274970 96792
rect 274730 96620 274786 96656
rect 274730 96600 274732 96620
rect 274732 96600 274784 96620
rect 274784 96600 274786 96620
rect 274638 86964 274694 87000
rect 274638 86944 274640 86964
rect 274640 86944 274692 86964
rect 274692 86944 274694 86964
rect 276110 85584 276166 85640
rect 276294 85584 276350 85640
rect 338670 115912 338726 115968
rect 339038 115912 339094 115968
rect 376758 6876 376760 6896
rect 376760 6876 376812 6896
rect 376812 6876 376814 6896
rect 376758 6840 376814 6876
rect 379610 6840 379666 6896
rect 383106 106256 383162 106312
rect 383290 106256 383346 106312
rect 383198 77152 383254 77208
rect 383290 28872 383346 28928
rect 383382 21936 383438 21992
rect 383658 117444 383660 117464
rect 383660 117444 383712 117464
rect 383712 117444 383714 117464
rect 383658 117408 383714 117444
rect 383658 77152 383714 77208
rect 393226 117544 393282 117600
rect 420734 77152 420790 77208
rect 420458 48320 420514 48376
rect 420642 48320 420698 48376
rect 420458 29008 420514 29064
rect 420642 28974 420698 29030
rect 421010 77152 421066 77208
rect 425978 86944 426034 87000
rect 426162 86944 426218 87000
rect 426070 64912 426126 64968
rect 425794 44104 425850 44160
rect 425978 44104 426034 44160
rect 426438 64912 426494 64968
rect 431314 114688 431370 114744
rect 431590 114552 431646 114608
rect 431590 66272 431646 66328
rect 431774 66272 431830 66328
rect 436466 193976 436522 194032
rect 436834 198872 436890 198928
rect 436742 182008 436798 182064
rect 436650 177928 436706 177984
rect 436558 176160 436614 176216
rect 437386 152224 437442 152280
rect 437018 150184 437074 150240
rect 437386 144472 437442 144528
rect 580170 697992 580226 698048
rect 580170 686296 580226 686352
rect 580170 674600 580226 674656
rect 580170 651072 580226 651128
rect 580170 639376 580226 639432
rect 580170 627680 580226 627736
rect 580170 604152 580226 604208
rect 580170 592456 580226 592512
rect 580170 580760 580226 580816
rect 580446 557232 580502 557288
rect 580354 545536 580410 545592
rect 580262 533840 580318 533896
rect 456798 375128 456854 375184
rect 457442 357992 457498 358048
rect 504730 378392 504786 378448
rect 504730 360440 504786 360496
rect 503718 340856 503774 340912
rect 504730 343576 504786 343632
rect 503902 340856 503958 340912
rect 503902 321680 503958 321736
rect 503902 321408 503958 321464
rect 504270 260888 504326 260944
rect 504546 260888 504602 260944
rect 579894 498616 579950 498672
rect 580170 486784 580226 486840
rect 580170 463392 580226 463448
rect 579894 451696 579950 451752
rect 579802 416472 579858 416528
rect 579986 346024 580042 346080
rect 580170 322632 580226 322688
rect 580170 310800 580226 310856
rect 579986 275712 580042 275768
rect 580170 263880 580226 263936
rect 580170 252184 580226 252240
rect 580078 228792 580134 228848
rect 579802 216960 579858 217016
rect 580078 205264 580134 205320
rect 504362 183504 504418 183560
rect 504638 183504 504694 183560
rect 579986 181872 580042 181928
rect 504178 154536 504234 154592
rect 504454 154536 504510 154592
rect 437386 140256 437442 140312
rect 437386 137808 437442 137864
rect 437018 136040 437074 136096
rect 437386 133592 437442 133648
rect 436834 131960 436890 132016
rect 580538 510312 580594 510368
rect 580446 439864 580502 439920
rect 580354 170040 580410 170096
rect 580262 134816 580318 134872
rect 437386 129512 437442 129568
rect 436926 124480 436982 124536
rect 436834 122848 436890 122904
rect 436742 120400 436798 120456
rect 580630 404776 580686 404832
rect 580538 392944 580594 393000
rect 580722 369552 580778 369608
rect 580906 357856 580962 357912
rect 580814 299104 580870 299160
rect 580630 158344 580686 158400
rect 580906 123120 580962 123176
rect 579802 111424 579858 111480
rect 580170 87896 580226 87952
rect 580170 76200 580226 76256
rect 579802 64504 579858 64560
rect 580170 40976 580226 41032
rect 580170 29280 580226 29336
rect 579802 17584 579858 17640
<< metal3 >>
rect 580165 698050 580231 698053
rect 583520 698050 584960 698140
rect 580165 698048 584960 698050
rect 580165 697992 580170 698048
rect 580226 697992 584960 698048
rect 580165 697990 584960 697992
rect 580165 697987 580231 697990
rect 583520 697900 584960 697990
rect -960 696540 480 696780
rect 580165 686354 580231 686357
rect 583520 686354 584960 686444
rect 580165 686352 584960 686354
rect 580165 686296 580170 686352
rect 580226 686296 584960 686352
rect 580165 686294 584960 686296
rect 580165 686291 580231 686294
rect 583520 686204 584960 686294
rect -960 682274 480 682364
rect 3785 682274 3851 682277
rect -960 682272 3851 682274
rect -960 682216 3790 682272
rect 3846 682216 3851 682272
rect -960 682214 3851 682216
rect -960 682124 480 682214
rect 3785 682211 3851 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 3509 653578 3575 653581
rect -960 653576 3575 653578
rect -960 653520 3514 653576
rect 3570 653520 3575 653576
rect -960 653518 3575 653520
rect -960 653428 480 653518
rect 3509 653515 3575 653518
rect 580165 651130 580231 651133
rect 583520 651130 584960 651220
rect 580165 651128 584960 651130
rect 580165 651072 580170 651128
rect 580226 651072 584960 651128
rect 580165 651070 584960 651072
rect 580165 651067 580231 651070
rect 583520 650980 584960 651070
rect 580165 639434 580231 639437
rect 583520 639434 584960 639524
rect 580165 639432 584960 639434
rect 580165 639376 580170 639432
rect 580226 639376 584960 639432
rect 580165 639374 584960 639376
rect 580165 639371 580231 639374
rect 583520 639284 584960 639374
rect -960 639012 480 639252
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3049 624882 3115 624885
rect -960 624880 3115 624882
rect -960 624824 3054 624880
rect 3110 624824 3115 624880
rect -960 624822 3115 624824
rect -960 624732 480 624822
rect 3049 624819 3115 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3601 610466 3667 610469
rect -960 610464 3667 610466
rect -960 610408 3606 610464
rect 3662 610408 3667 610464
rect -960 610406 3667 610408
rect -960 610316 480 610406
rect 3601 610403 3667 610406
rect 580165 604210 580231 604213
rect 583520 604210 584960 604300
rect 580165 604208 584960 604210
rect 580165 604152 580170 604208
rect 580226 604152 584960 604208
rect 580165 604150 584960 604152
rect 580165 604147 580231 604150
rect 583520 604060 584960 604150
rect -960 596050 480 596140
rect 3693 596050 3759 596053
rect -960 596048 3759 596050
rect -960 595992 3698 596048
rect 3754 595992 3759 596048
rect -960 595990 3759 595992
rect -960 595900 480 595990
rect 3693 595987 3759 595990
rect 580165 592514 580231 592517
rect 583520 592514 584960 592604
rect 580165 592512 584960 592514
rect 580165 592456 580170 592512
rect 580226 592456 584960 592512
rect 580165 592454 584960 592456
rect 580165 592451 580231 592454
rect 583520 592364 584960 592454
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 305177 579322 305243 579325
rect 315849 579322 315915 579325
rect 305177 579320 315915 579322
rect 305177 579264 305182 579320
rect 305238 579264 315854 579320
rect 315910 579264 315915 579320
rect 305177 579262 315915 579264
rect 305177 579259 305243 579262
rect 315849 579259 315915 579262
rect 289813 578914 289879 578917
rect 299381 578914 299447 578917
rect 289813 578912 299447 578914
rect 289813 578856 289818 578912
rect 289874 578856 299386 578912
rect 299442 578856 299447 578912
rect 289813 578854 299447 578856
rect 289813 578851 289879 578854
rect 299381 578851 299447 578854
rect 116025 578370 116091 578373
rect 125501 578370 125567 578373
rect 116025 578368 125567 578370
rect 116025 578312 116030 578368
rect 116086 578312 125506 578368
rect 125562 578312 125567 578368
rect 116025 578310 125567 578312
rect 116025 578307 116091 578310
rect 125501 578307 125567 578310
rect 296713 575786 296779 575789
rect 299982 575786 300042 576232
rect 296713 575784 300042 575786
rect 296713 575728 296718 575784
rect 296774 575728 300042 575784
rect 296713 575726 300042 575728
rect 296713 575723 296779 575726
rect 377814 575514 377874 575960
rect 380525 575514 380591 575517
rect 377814 575512 380591 575514
rect 377814 575456 380530 575512
rect 380586 575456 380591 575512
rect 377814 575454 380591 575456
rect 380525 575451 380591 575454
rect 297357 572930 297423 572933
rect 299982 572930 300042 572968
rect 297357 572928 300042 572930
rect 297357 572872 297362 572928
rect 297418 572872 300042 572928
rect 297357 572870 300042 572872
rect 297357 572867 297423 572870
rect 377446 572117 377506 572696
rect 377397 572112 377506 572117
rect 377397 572056 377402 572112
rect 377458 572056 377506 572112
rect 377397 572054 377506 572056
rect 377397 572051 377463 572054
rect 296713 570074 296779 570077
rect 296713 570072 300042 570074
rect 296713 570016 296718 570072
rect 296774 570016 300042 570072
rect 296713 570014 300042 570016
rect 296713 570011 296779 570014
rect 299982 569976 300042 570014
rect 378133 569734 378199 569737
rect 377844 569732 378199 569734
rect 377844 569676 378138 569732
rect 378194 569676 378199 569732
rect 377844 569674 378199 569676
rect 378133 569671 378199 569674
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3877 567354 3943 567357
rect -960 567352 3943 567354
rect -960 567296 3882 567352
rect 3938 567296 3943 567352
rect -960 567294 3943 567296
rect -960 567204 480 567294
rect 3877 567291 3943 567294
rect 296437 566130 296503 566133
rect 299982 566130 300042 566712
rect 378225 566470 378291 566473
rect 377844 566468 378291 566470
rect 377844 566412 378230 566468
rect 378286 566412 378291 566468
rect 377844 566410 378291 566412
rect 378225 566407 378291 566410
rect 296437 566128 300042 566130
rect 296437 566072 296442 566128
rect 296498 566072 300042 566128
rect 296437 566070 300042 566072
rect 296437 566067 296503 566070
rect 296713 563274 296779 563277
rect 299982 563274 300042 563720
rect 378317 563478 378383 563481
rect 377844 563476 378383 563478
rect 377844 563420 378322 563476
rect 378378 563420 378383 563476
rect 377844 563418 378383 563420
rect 378317 563415 378383 563418
rect 296713 563272 300042 563274
rect 296713 563216 296718 563272
rect 296774 563216 300042 563272
rect 296713 563214 300042 563216
rect 296713 563211 296779 563214
rect 271781 563138 271847 563141
rect 271646 563136 271847 563138
rect 271646 563080 271786 563136
rect 271842 563080 271847 563136
rect 271646 563078 271847 563080
rect 271646 563005 271706 563078
rect 271781 563075 271847 563078
rect 271646 563000 271755 563005
rect 271646 562944 271694 563000
rect 271750 562944 271755 563000
rect 271646 562942 271755 562944
rect 271689 562939 271755 562942
rect 297909 560418 297975 560421
rect 299982 560418 300042 560456
rect 297909 560416 300042 560418
rect 297909 560360 297914 560416
rect 297970 560360 300042 560416
rect 297909 560358 300042 560360
rect 297909 560355 297975 560358
rect 271505 560282 271571 560285
rect 271689 560282 271755 560285
rect 271505 560280 271755 560282
rect 271505 560224 271510 560280
rect 271566 560224 271694 560280
rect 271750 560224 271755 560280
rect 271505 560222 271755 560224
rect 271505 560219 271571 560222
rect 271689 560219 271755 560222
rect 377814 559602 377874 560184
rect 378409 559602 378475 559605
rect 377814 559600 378475 559602
rect 377814 559544 378414 559600
rect 378470 559544 378475 559600
rect 377814 559542 378475 559544
rect 378409 559539 378475 559542
rect 198641 556746 198707 556749
rect 200070 556746 200130 557328
rect 297817 556882 297883 556885
rect 299982 556882 300042 557464
rect 580441 557290 580507 557293
rect 583520 557290 584960 557380
rect 580441 557288 584960 557290
rect 580441 557232 580446 557288
rect 580502 557232 584960 557288
rect 580441 557230 584960 557232
rect 580441 557227 580507 557230
rect 297817 556880 300042 556882
rect 297817 556824 297822 556880
rect 297878 556824 300042 556880
rect 297817 556822 300042 556824
rect 297817 556819 297883 556822
rect 198641 556744 200130 556746
rect 198641 556688 198646 556744
rect 198702 556688 200130 556744
rect 198641 556686 200130 556688
rect 198641 556683 198707 556686
rect 219942 556202 220002 556784
rect 377814 556610 377874 557192
rect 583520 557140 584960 557230
rect 378593 556610 378659 556613
rect 377814 556608 378659 556610
rect 377814 556552 378598 556608
rect 378654 556552 378659 556608
rect 377814 556550 378659 556552
rect 378593 556547 378659 556550
rect 222193 556202 222259 556205
rect 219942 556200 222259 556202
rect 219942 556144 222198 556200
rect 222254 556144 222259 556200
rect 219942 556142 222259 556144
rect 222193 556139 222259 556142
rect 297817 553618 297883 553621
rect 299982 553618 300042 554200
rect 297817 553616 300042 553618
rect 297817 553560 297822 553616
rect 297878 553560 300042 553616
rect 297817 553558 300042 553560
rect 297817 553555 297883 553558
rect 377814 553482 377874 553928
rect 379513 553482 379579 553485
rect 377814 553480 379579 553482
rect 377814 553424 379518 553480
rect 379574 553424 379579 553480
rect 377814 553422 379579 553424
rect 379513 553419 379579 553422
rect -960 553074 480 553164
rect 3785 553074 3851 553077
rect -960 553072 3851 553074
rect -960 553016 3790 553072
rect 3846 553016 3851 553072
rect -960 553014 3851 553016
rect -960 552924 480 553014
rect 3785 553011 3851 553014
rect 198549 552122 198615 552125
rect 200070 552122 200130 552704
rect 198549 552120 200130 552122
rect 198549 552064 198554 552120
rect 198610 552064 200130 552120
rect 198549 552062 200130 552064
rect 219942 552122 220002 552160
rect 222285 552122 222351 552125
rect 219942 552120 222351 552122
rect 219942 552064 222290 552120
rect 222346 552064 222351 552120
rect 219942 552062 222351 552064
rect 198549 552059 198615 552062
rect 222285 552059 222351 552062
rect 297725 550762 297791 550765
rect 299982 550762 300042 550936
rect 378685 550762 378751 550765
rect 297725 550760 300042 550762
rect 297725 550704 297730 550760
rect 297786 550704 300042 550760
rect 297725 550702 300042 550704
rect 377814 550760 378751 550762
rect 377814 550704 378690 550760
rect 378746 550704 378751 550760
rect 377814 550702 378751 550704
rect 297725 550699 297791 550702
rect 377814 550664 377874 550702
rect 378685 550699 378751 550702
rect 86358 549949 86418 550528
rect 86358 549944 86467 549949
rect 86358 549888 86406 549944
rect 86462 549888 86467 549944
rect 86358 549886 86467 549888
rect 86401 549883 86467 549886
rect 198917 547906 198983 547909
rect 200070 547906 200130 548080
rect 198917 547904 200130 547906
rect 198917 547848 198922 547904
rect 198978 547848 200130 547904
rect 198917 547846 200130 547848
rect 299105 547906 299171 547909
rect 299982 547906 300042 547944
rect 299105 547904 300042 547906
rect 299105 547848 299110 547904
rect 299166 547848 300042 547904
rect 299105 547846 300042 547848
rect 198917 547843 198983 547846
rect 299105 547843 299171 547846
rect 219942 546954 220002 547536
rect 377814 547090 377874 547672
rect 378869 547090 378935 547093
rect 377814 547088 378935 547090
rect 377814 547032 378874 547088
rect 378930 547032 378935 547088
rect 377814 547030 378935 547032
rect 378869 547027 378935 547030
rect 222377 546954 222443 546957
rect 219942 546952 222443 546954
rect 219942 546896 222382 546952
rect 222438 546896 222443 546952
rect 219942 546894 222443 546896
rect 222377 546891 222443 546894
rect 115614 546546 115674 546720
rect 118049 546546 118115 546549
rect 115614 546544 118115 546546
rect 115614 546488 118054 546544
rect 118110 546488 118115 546544
rect 115614 546486 118115 546488
rect 118049 546483 118115 546486
rect 84101 545866 84167 545869
rect 85990 545866 86050 546448
rect 84101 545864 86050 545866
rect 84101 545808 84106 545864
rect 84162 545808 86050 545864
rect 84101 545806 86050 545808
rect 84101 545803 84167 545806
rect 580349 545594 580415 545597
rect 583520 545594 584960 545684
rect 580349 545592 584960 545594
rect 580349 545536 580354 545592
rect 580410 545536 584960 545592
rect 580349 545534 584960 545536
rect 580349 545531 580415 545534
rect 583520 545444 584960 545534
rect 299013 544098 299079 544101
rect 299982 544098 300042 544680
rect 299013 544096 300042 544098
rect 299013 544040 299018 544096
rect 299074 544040 300042 544096
rect 299013 544038 300042 544040
rect 299013 544035 299079 544038
rect 198457 543826 198523 543829
rect 377814 543826 377874 544408
rect 379605 543826 379671 543829
rect 198457 543824 200130 543826
rect 198457 543768 198462 543824
rect 198518 543768 200130 543824
rect 198457 543766 200130 543768
rect 377814 543824 379671 543826
rect 377814 543768 379610 543824
rect 379666 543768 379671 543824
rect 377814 543766 379671 543768
rect 198457 543763 198523 543766
rect 200070 543728 200130 543766
rect 379605 543763 379671 543766
rect 219942 542602 220002 543184
rect 222469 542602 222535 542605
rect 219942 542600 222535 542602
rect 219942 542544 222474 542600
rect 222530 542544 222535 542600
rect 219942 542542 222535 542544
rect 222469 542539 222535 542542
rect 118601 542466 118667 542469
rect 115614 542464 118667 542466
rect 115614 542408 118606 542464
rect 118662 542408 118667 542464
rect 115614 542406 118667 542408
rect 115614 542368 115674 542406
rect 118601 542403 118667 542406
rect 84009 541514 84075 541517
rect 85990 541514 86050 542096
rect 84009 541512 86050 541514
rect 84009 541456 84014 541512
rect 84070 541456 86050 541512
rect 84009 541454 86050 541456
rect 84009 541451 84075 541454
rect 297265 541106 297331 541109
rect 299982 541106 300042 541688
rect 297265 541104 300042 541106
rect 297265 541048 297270 541104
rect 297326 541048 300042 541104
rect 297265 541046 300042 541048
rect 377814 541106 377874 541416
rect 380341 541106 380407 541109
rect 377814 541104 380407 541106
rect 377814 541048 380346 541104
rect 380402 541048 380407 541104
rect 377814 541046 380407 541048
rect 297265 541043 297331 541046
rect 380341 541043 380407 541046
rect 271689 540970 271755 540973
rect 271965 540970 272031 540973
rect 271689 540968 272031 540970
rect 271689 540912 271694 540968
rect 271750 540912 271970 540968
rect 272026 540912 272031 540968
rect 271689 540910 272031 540912
rect 271689 540907 271755 540910
rect 271965 540907 272031 540910
rect -960 538658 480 538748
rect 3969 538658 4035 538661
rect -960 538656 4035 538658
rect -960 538600 3974 538656
rect 4030 538600 4035 538656
rect -960 538598 4035 538600
rect -960 538508 480 538598
rect 3969 538595 4035 538598
rect 198365 538522 198431 538525
rect 200070 538522 200130 539104
rect 198365 538520 200130 538522
rect 198365 538464 198370 538520
rect 198426 538464 200130 538520
rect 198365 538462 200130 538464
rect 198365 538459 198431 538462
rect 219942 538386 220002 538560
rect 222561 538386 222627 538389
rect 219942 538384 222627 538386
rect 219942 538328 222566 538384
rect 222622 538328 222627 538384
rect 219942 538326 222627 538328
rect 222561 538323 222627 538326
rect 297633 538386 297699 538389
rect 299982 538386 300042 538424
rect 297633 538384 300042 538386
rect 297633 538328 297638 538384
rect 297694 538328 300042 538384
rect 297633 538326 300042 538328
rect 297633 538323 297699 538326
rect 85573 537774 85639 537777
rect 85573 537772 86020 537774
rect 85573 537716 85578 537772
rect 85634 537744 86020 537772
rect 85634 537716 86050 537744
rect 85573 537714 86050 537716
rect 85573 537711 85639 537714
rect 83917 537162 83983 537165
rect 85990 537162 86050 537714
rect 115614 537434 115674 538016
rect 377814 537570 377874 538152
rect 379697 537570 379763 537573
rect 377814 537568 379763 537570
rect 377814 537512 379702 537568
rect 379758 537512 379763 537568
rect 377814 537510 379763 537512
rect 379697 537507 379763 537510
rect 117773 537434 117839 537437
rect 115614 537432 117839 537434
rect 115614 537376 117778 537432
rect 117834 537376 117839 537432
rect 115614 537374 117839 537376
rect 117773 537371 117839 537374
rect 83917 537160 86050 537162
rect 83917 537104 83922 537160
rect 83978 537104 86050 537160
rect 83917 537102 86050 537104
rect 83917 537099 83983 537102
rect 297633 534850 297699 534853
rect 299982 534850 300042 535432
rect 297633 534848 300042 534850
rect 297633 534792 297638 534848
rect 297694 534792 300042 534848
rect 297633 534790 300042 534792
rect 297633 534787 297699 534790
rect 377814 534578 377874 535160
rect 379789 534578 379855 534581
rect 377814 534576 379855 534578
rect 377814 534520 379794 534576
rect 379850 534520 379855 534576
rect 377814 534518 379855 534520
rect 379789 534515 379855 534518
rect 198733 534170 198799 534173
rect 200070 534170 200130 534480
rect 198733 534168 200130 534170
rect 198733 534112 198738 534168
rect 198794 534112 200130 534168
rect 198733 534110 200130 534112
rect 198733 534107 198799 534110
rect 85297 533082 85363 533085
rect 85990 533082 86050 533664
rect 115614 533354 115674 533936
rect 117773 533354 117839 533357
rect 115614 533352 117839 533354
rect 115614 533296 117778 533352
rect 117834 533296 117839 533352
rect 115614 533294 117839 533296
rect 219942 533354 220002 533936
rect 580257 533898 580323 533901
rect 583520 533898 584960 533988
rect 580257 533896 584960 533898
rect 580257 533840 580262 533896
rect 580318 533840 584960 533896
rect 580257 533838 584960 533840
rect 580257 533835 580323 533838
rect 583520 533748 584960 533838
rect 222653 533354 222719 533357
rect 219942 533352 222719 533354
rect 219942 533296 222658 533352
rect 222714 533296 222719 533352
rect 219942 533294 222719 533296
rect 117773 533291 117839 533294
rect 222653 533291 222719 533294
rect 85297 533080 86050 533082
rect 85297 533024 85302 533080
rect 85358 533024 86050 533080
rect 85297 533022 86050 533024
rect 85297 533019 85363 533022
rect 296529 531586 296595 531589
rect 299982 531586 300042 532168
rect 296529 531584 300042 531586
rect 296529 531528 296534 531584
rect 296590 531528 300042 531584
rect 296529 531526 300042 531528
rect 296529 531523 296595 531526
rect 377814 531450 377874 531896
rect 379881 531450 379947 531453
rect 377814 531448 379947 531450
rect 377814 531392 379886 531448
rect 379942 531392 379947 531448
rect 377814 531390 379947 531392
rect 379881 531387 379947 531390
rect 8109 531314 8175 531317
rect 8385 531314 8451 531317
rect 8109 531312 8451 531314
rect 8109 531256 8114 531312
rect 8170 531256 8390 531312
rect 8446 531256 8451 531312
rect 8109 531254 8451 531256
rect 8109 531251 8175 531254
rect 8385 531251 8451 531254
rect 117957 529682 118023 529685
rect 115614 529680 118023 529682
rect 115614 529624 117962 529680
rect 118018 529624 118023 529680
rect 115614 529622 118023 529624
rect 115614 529584 115674 529622
rect 117957 529619 118023 529622
rect 83825 528730 83891 528733
rect 85990 528730 86050 529312
rect 198825 529274 198891 529277
rect 200070 529274 200130 529856
rect 198825 529272 200130 529274
rect 198825 529216 198830 529272
rect 198886 529216 200130 529272
rect 198825 529214 200130 529216
rect 198825 529211 198891 529214
rect 219390 529005 219450 529312
rect 219390 529000 219499 529005
rect 219390 528944 219438 529000
rect 219494 528944 219499 529000
rect 219390 528942 219499 528944
rect 219433 528939 219499 528942
rect 83825 528728 86050 528730
rect 83825 528672 83830 528728
rect 83886 528672 86050 528728
rect 83825 528670 86050 528672
rect 83825 528667 83891 528670
rect 297357 528594 297423 528597
rect 299982 528594 300042 529176
rect 377814 528730 377874 528904
rect 380433 528730 380499 528733
rect 377814 528728 380499 528730
rect 377814 528672 380438 528728
rect 380494 528672 380499 528728
rect 377814 528670 380499 528672
rect 380433 528667 380499 528670
rect 297357 528592 300042 528594
rect 297357 528536 297362 528592
rect 297418 528536 300042 528592
rect 297357 528534 300042 528536
rect 297357 528531 297423 528534
rect 297449 525874 297515 525877
rect 299982 525874 300042 525912
rect 297449 525872 300042 525874
rect 297449 525816 297454 525872
rect 297510 525816 300042 525872
rect 297449 525814 300042 525816
rect 297449 525811 297515 525814
rect 85389 525602 85455 525605
rect 85389 525600 86050 525602
rect 85389 525544 85394 525600
rect 85450 525544 86050 525600
rect 85389 525542 86050 525544
rect 85389 525539 85455 525542
rect 82813 524922 82879 524925
rect 85990 524922 86050 525542
rect 115614 525194 115674 525232
rect 118601 525194 118667 525197
rect 115614 525192 118667 525194
rect 115614 525136 118606 525192
rect 118662 525136 118667 525192
rect 115614 525134 118667 525136
rect 118601 525131 118667 525134
rect 82813 524920 86050 524922
rect 82813 524864 82818 524920
rect 82874 524864 86050 524920
rect 82813 524862 86050 524864
rect 82813 524859 82879 524862
rect 198273 524650 198339 524653
rect 200070 524650 200130 525232
rect 377814 525058 377874 525640
rect 379973 525058 380039 525061
rect 377814 525056 380039 525058
rect 377814 525000 379978 525056
rect 380034 525000 380039 525056
rect 377814 524998 380039 525000
rect 379973 524995 380039 524998
rect 198273 524648 200130 524650
rect 198273 524592 198278 524648
rect 198334 524592 200130 524648
rect 198273 524590 200130 524592
rect 198273 524587 198339 524590
rect 219574 524517 219634 524688
rect 219525 524512 219634 524517
rect 219525 524456 219530 524512
rect 219586 524456 219634 524512
rect 219525 524454 219634 524456
rect 219525 524451 219591 524454
rect -960 524092 480 524332
rect 297541 522066 297607 522069
rect 299982 522066 300042 522648
rect 297541 522064 300042 522066
rect 297541 522008 297546 522064
rect 297602 522008 300042 522064
rect 297541 522006 300042 522008
rect 297541 522003 297607 522006
rect 281257 521930 281323 521933
rect 281214 521928 281323 521930
rect 281214 521872 281262 521928
rect 281318 521872 281323 521928
rect 281214 521867 281323 521872
rect 281214 521692 281274 521867
rect 377814 521794 377874 522376
rect 583520 521916 584960 522156
rect 378501 521794 378567 521797
rect 377814 521792 378567 521794
rect 377814 521736 378506 521792
rect 378562 521736 378567 521792
rect 377814 521734 378567 521736
rect 378501 521731 378567 521734
rect 281349 521692 281415 521695
rect 281214 521690 281415 521692
rect 281214 521634 281354 521690
rect 281410 521634 281415 521690
rect 281214 521632 281415 521634
rect 281349 521629 281415 521632
rect 115614 521114 115674 521152
rect 117313 521114 117379 521117
rect 115614 521112 117379 521114
rect 115614 521056 117318 521112
rect 117374 521056 117379 521112
rect 115614 521054 117379 521056
rect 117313 521051 117379 521054
rect 297449 519074 297515 519077
rect 299982 519074 300042 519656
rect 377630 519213 377690 519384
rect 377630 519208 377739 519213
rect 377630 519152 377678 519208
rect 377734 519152 377739 519208
rect 377630 519150 377739 519152
rect 377673 519147 377739 519150
rect 297449 519072 300042 519074
rect 297449 519016 297454 519072
rect 297510 519016 300042 519072
rect 297449 519014 300042 519016
rect 297449 519011 297515 519014
rect 297449 516218 297515 516221
rect 299982 516218 300042 516392
rect 297449 516216 300042 516218
rect 297449 516160 297454 516216
rect 297510 516160 300042 516216
rect 297449 516158 300042 516160
rect 297449 516155 297515 516158
rect 377814 515538 377874 516120
rect 380065 515538 380131 515541
rect 377814 515536 380131 515538
rect 377814 515480 380070 515536
rect 380126 515480 380131 515536
rect 377814 515478 380131 515480
rect 380065 515475 380131 515478
rect 297449 513498 297515 513501
rect 297449 513496 300042 513498
rect 297449 513440 297454 513496
rect 297510 513440 300042 513496
rect 297449 513438 300042 513440
rect 297449 513435 297515 513438
rect 299982 513400 300042 513438
rect 377814 512546 377874 513128
rect 380157 512546 380223 512549
rect 377814 512544 380223 512546
rect 377814 512488 380162 512544
rect 380218 512488 380223 512544
rect 377814 512486 380223 512488
rect 380157 512483 380223 512486
rect 8109 512002 8175 512005
rect 8385 512002 8451 512005
rect 8109 512000 8451 512002
rect 8109 511944 8114 512000
rect 8170 511944 8390 512000
rect 8446 511944 8451 512000
rect 8109 511942 8451 511944
rect 8109 511939 8175 511942
rect 8385 511939 8451 511942
rect 580533 510370 580599 510373
rect 583520 510370 584960 510460
rect 580533 510368 584960 510370
rect 580533 510312 580538 510368
rect 580594 510312 584960 510368
rect 580533 510310 584960 510312
rect 580533 510307 580599 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 4061 509962 4127 509965
rect -960 509960 4127 509962
rect -960 509904 4066 509960
rect 4122 509904 4127 509960
rect -960 509902 4127 509904
rect -960 509812 480 509902
rect 4061 509899 4127 509902
rect 296713 509554 296779 509557
rect 299982 509554 300042 510136
rect 296713 509552 300042 509554
rect 296713 509496 296718 509552
rect 296774 509496 300042 509552
rect 296713 509494 300042 509496
rect 377814 509554 377874 509864
rect 380249 509554 380315 509557
rect 377814 509552 380315 509554
rect 377814 509496 380254 509552
rect 380310 509496 380315 509552
rect 377814 509494 380315 509496
rect 296713 509491 296779 509494
rect 380249 509491 380315 509494
rect 296713 506562 296779 506565
rect 299982 506562 300042 507144
rect 296713 506560 300042 506562
rect 296713 506504 296718 506560
rect 296774 506504 300042 506560
rect 296713 506502 300042 506504
rect 377814 506562 377874 506872
rect 380341 506562 380407 506565
rect 377814 506560 380407 506562
rect 377814 506504 380346 506560
rect 380402 506504 380407 506560
rect 377814 506502 380407 506504
rect 296713 506499 296779 506502
rect 380341 506499 380407 506502
rect 297357 503842 297423 503845
rect 299982 503842 300042 503880
rect 297357 503840 300042 503842
rect 297357 503784 297362 503840
rect 297418 503784 300042 503840
rect 297357 503782 300042 503784
rect 297357 503779 297423 503782
rect 377814 503026 377874 503608
rect 380709 503026 380775 503029
rect 377814 503024 380775 503026
rect 377814 502968 380714 503024
rect 380770 502968 380775 503024
rect 377814 502966 380775 502968
rect 380709 502963 380775 502966
rect 271597 502348 271663 502349
rect 271597 502344 271644 502348
rect 271708 502346 271714 502348
rect 271597 502288 271602 502344
rect 271597 502284 271644 502288
rect 271708 502286 271754 502346
rect 271708 502284 271714 502286
rect 271597 502283 271663 502284
rect 579889 498674 579955 498677
rect 583520 498674 584960 498764
rect 579889 498672 584960 498674
rect 579889 498616 579894 498672
rect 579950 498616 584960 498672
rect 579889 498614 584960 498616
rect 579889 498611 579955 498614
rect 583520 498524 584960 498614
rect -960 495546 480 495636
rect 3969 495546 4035 495549
rect -960 495544 4035 495546
rect -960 495488 3974 495544
rect 4030 495488 4035 495544
rect -960 495486 4035 495488
rect -960 495396 480 495486
rect 3969 495483 4035 495486
rect 271638 492628 271644 492692
rect 271708 492690 271714 492692
rect 271781 492690 271847 492693
rect 271708 492688 271847 492690
rect 271708 492632 271786 492688
rect 271842 492632 271847 492688
rect 271708 492630 271847 492632
rect 271708 492628 271714 492630
rect 271781 492627 271847 492630
rect 281073 492690 281139 492693
rect 281257 492690 281323 492693
rect 281073 492688 281323 492690
rect 281073 492632 281078 492688
rect 281134 492632 281262 492688
rect 281318 492632 281323 492688
rect 281073 492630 281323 492632
rect 281073 492627 281139 492630
rect 281257 492627 281323 492630
rect 580165 486842 580231 486845
rect 583520 486842 584960 486932
rect 580165 486840 584960 486842
rect 580165 486784 580170 486840
rect 580226 486784 584960 486840
rect 580165 486782 584960 486784
rect 580165 486779 580231 486782
rect 583520 486692 584960 486782
rect 307017 483170 307083 483173
rect 307017 483168 307218 483170
rect 307017 483112 307022 483168
rect 307078 483112 307218 483168
rect 307017 483110 307218 483112
rect 307017 483107 307083 483110
rect 307017 483034 307083 483037
rect 307158 483034 307218 483110
rect 307017 483032 307218 483034
rect 307017 482976 307022 483032
rect 307078 482976 307218 483032
rect 307017 482974 307218 482976
rect 307017 482971 307083 482974
rect -960 481130 480 481220
rect 3141 481130 3207 481133
rect -960 481128 3207 481130
rect -960 481072 3146 481128
rect 3202 481072 3207 481128
rect -960 481070 3207 481072
rect -960 480980 480 481070
rect 3141 481067 3207 481070
rect 583520 474996 584960 475236
rect 7925 473378 7991 473381
rect 8109 473378 8175 473381
rect 7925 473376 8175 473378
rect 7925 473320 7930 473376
rect 7986 473320 8114 473376
rect 8170 473320 8175 473376
rect 7925 473318 8175 473320
rect 7925 473315 7991 473318
rect 8109 473315 8175 473318
rect 301865 473378 301931 473381
rect 302049 473378 302115 473381
rect 301865 473376 302115 473378
rect 301865 473320 301870 473376
rect 301926 473320 302054 473376
rect 302110 473320 302115 473376
rect 301865 473318 302115 473320
rect 301865 473315 301931 473318
rect 302049 473315 302115 473318
rect -960 466700 480 466940
rect 307017 463858 307083 463861
rect 307017 463856 307218 463858
rect 307017 463800 307022 463856
rect 307078 463800 307218 463856
rect 307017 463798 307218 463800
rect 307017 463795 307083 463798
rect 307017 463722 307083 463725
rect 307158 463722 307218 463798
rect 307017 463720 307218 463722
rect 307017 463664 307022 463720
rect 307078 463664 307218 463720
rect 307017 463662 307218 463664
rect 307017 463659 307083 463662
rect 580165 463450 580231 463453
rect 583520 463450 584960 463540
rect 580165 463448 584960 463450
rect 580165 463392 580170 463448
rect 580226 463392 584960 463448
rect 580165 463390 584960 463392
rect 580165 463387 580231 463390
rect 583520 463300 584960 463390
rect 281073 454066 281139 454069
rect 281257 454066 281323 454069
rect 281073 454064 281323 454066
rect 281073 454008 281078 454064
rect 281134 454008 281262 454064
rect 281318 454008 281323 454064
rect 281073 454006 281323 454008
rect 281073 454003 281139 454006
rect 281257 454003 281323 454006
rect 306833 454066 306899 454069
rect 307017 454066 307083 454069
rect 306833 454064 307083 454066
rect 306833 454008 306838 454064
rect 306894 454008 307022 454064
rect 307078 454008 307083 454064
rect 306833 454006 307083 454008
rect 306833 454003 306899 454006
rect 307017 454003 307083 454006
rect -960 452434 480 452524
rect 3233 452434 3299 452437
rect -960 452432 3299 452434
rect -960 452376 3238 452432
rect 3294 452376 3299 452432
rect -960 452374 3299 452376
rect -960 452284 480 452374
rect 3233 452371 3299 452374
rect 579889 451754 579955 451757
rect 583520 451754 584960 451844
rect 579889 451752 584960 451754
rect 579889 451696 579894 451752
rect 579950 451696 584960 451752
rect 579889 451694 584960 451696
rect 579889 451691 579955 451694
rect 583520 451604 584960 451694
rect 580441 439922 580507 439925
rect 583520 439922 584960 440012
rect 580441 439920 584960 439922
rect 580441 439864 580446 439920
rect 580502 439864 584960 439920
rect 580441 439862 584960 439864
rect 580441 439859 580507 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3325 438018 3391 438021
rect -960 438016 3391 438018
rect -960 437960 3330 438016
rect 3386 437960 3391 438016
rect -960 437958 3391 437960
rect -960 437868 480 437958
rect 3325 437955 3391 437958
rect 281073 434754 281139 434757
rect 281257 434754 281323 434757
rect 281073 434752 281323 434754
rect 281073 434696 281078 434752
rect 281134 434696 281262 434752
rect 281318 434696 281323 434752
rect 281073 434694 281323 434696
rect 281073 434691 281139 434694
rect 281257 434691 281323 434694
rect 583520 428076 584960 428316
rect -960 423738 480 423828
rect 3233 423738 3299 423741
rect -960 423736 3299 423738
rect -960 423680 3238 423736
rect 3294 423680 3299 423736
rect -960 423678 3299 423680
rect -960 423588 480 423678
rect 3233 423675 3299 423678
rect 271781 419522 271847 419525
rect 271965 419522 272031 419525
rect 271781 419520 272031 419522
rect 271781 419464 271786 419520
rect 271842 419464 271970 419520
rect 272026 419464 272031 419520
rect 271781 419462 272031 419464
rect 271781 419459 271847 419462
rect 271965 419459 272031 419462
rect 579797 416530 579863 416533
rect 583520 416530 584960 416620
rect 579797 416528 584960 416530
rect 579797 416472 579802 416528
rect 579858 416472 584960 416528
rect 579797 416470 584960 416472
rect 579797 416467 579863 416470
rect 583520 416380 584960 416470
rect 265985 415442 266051 415445
rect 266169 415442 266235 415445
rect 265985 415440 266235 415442
rect 265985 415384 265990 415440
rect 266046 415384 266174 415440
rect 266230 415384 266235 415440
rect 265985 415382 266235 415384
rect 265985 415379 266051 415382
rect 266169 415379 266235 415382
rect -960 409172 480 409412
rect 580625 404834 580691 404837
rect 583520 404834 584960 404924
rect 580625 404832 584960 404834
rect 580625 404776 580630 404832
rect 580686 404776 584960 404832
rect 580625 404774 584960 404776
rect 580625 404771 580691 404774
rect 583520 404684 584960 404774
rect 199009 403746 199075 403749
rect 267733 403746 267799 403749
rect 199009 403744 200100 403746
rect 199009 403688 199014 403744
rect 199070 403688 200100 403744
rect 199009 403686 200100 403688
rect 266524 403744 267799 403746
rect 266524 403688 267738 403744
rect 267794 403688 267799 403744
rect 266524 403686 267799 403688
rect 199009 403683 199075 403686
rect 267733 403683 267799 403686
rect 198181 399666 198247 399669
rect 266813 399666 266879 399669
rect 198181 399664 200100 399666
rect 198181 399608 198186 399664
rect 198242 399608 200100 399664
rect 198181 399606 200100 399608
rect 266524 399664 266879 399666
rect 266524 399608 266818 399664
rect 266874 399608 266879 399664
rect 266524 399606 266879 399608
rect 198181 399603 198247 399606
rect 266813 399603 266879 399606
rect 281625 396130 281691 396133
rect 281398 396128 281691 396130
rect 281398 396072 281630 396128
rect 281686 396072 281691 396128
rect 281398 396070 281691 396072
rect 281398 395994 281458 396070
rect 281625 396067 281691 396070
rect 281625 395994 281691 395997
rect 281398 395992 281691 395994
rect 281398 395936 281630 395992
rect 281686 395936 281691 395992
rect 281398 395934 281691 395936
rect 281625 395931 281691 395934
rect 96613 395858 96679 395861
rect 99281 395858 99347 395861
rect 96613 395856 99347 395858
rect 96613 395800 96618 395856
rect 96674 395800 99286 395856
rect 99342 395800 99347 395856
rect 96613 395798 99347 395800
rect 96613 395795 96679 395798
rect 99281 395795 99347 395798
rect 199101 395314 199167 395317
rect 267825 395314 267891 395317
rect 199101 395312 200100 395314
rect 199101 395256 199106 395312
rect 199162 395256 200100 395312
rect 199101 395254 200100 395256
rect 266524 395312 267891 395314
rect 266524 395256 267830 395312
rect 267886 395256 267891 395312
rect 266524 395254 267891 395256
rect 199101 395251 199167 395254
rect 267825 395251 267891 395254
rect -960 395042 480 395132
rect 3049 395042 3115 395045
rect -960 395040 3115 395042
rect -960 394984 3054 395040
rect 3110 394984 3115 395040
rect -960 394982 3115 394984
rect -960 394892 480 394982
rect 3049 394979 3115 394982
rect 72325 393002 72391 393005
rect 580533 393002 580599 393005
rect 583520 393002 584960 393092
rect 72325 393000 72434 393002
rect 72325 392944 72330 393000
rect 72386 392944 72434 393000
rect 72325 392939 72434 392944
rect 580533 393000 584960 393002
rect 580533 392944 580538 393000
rect 580594 392944 584960 393000
rect 580533 392942 584960 392944
rect 580533 392939 580599 392942
rect 72374 392564 72434 392939
rect 583520 392852 584960 392942
rect 198089 391234 198155 391237
rect 267917 391234 267983 391237
rect 198089 391232 200100 391234
rect 198089 391176 198094 391232
rect 198150 391176 200100 391232
rect 198089 391174 200100 391176
rect 266524 391232 267983 391234
rect 266524 391176 267922 391232
rect 267978 391176 267983 391232
rect 266524 391174 267983 391176
rect 198089 391171 198155 391174
rect 267917 391171 267983 391174
rect 271597 389194 271663 389197
rect 271781 389194 271847 389197
rect 271597 389192 271847 389194
rect 271597 389136 271602 389192
rect 271658 389136 271786 389192
rect 271842 389136 271847 389192
rect 271597 389134 271847 389136
rect 271597 389131 271663 389134
rect 271781 389131 271847 389134
rect 128537 387970 128603 387973
rect 129089 387970 129155 387973
rect 126132 387968 129155 387970
rect 126132 387912 128542 387968
rect 128598 387912 129094 387968
rect 129150 387912 129155 387968
rect 126132 387910 129155 387912
rect 128537 387907 128603 387910
rect 129089 387907 129155 387910
rect 197997 387154 198063 387157
rect 197997 387152 200100 387154
rect 197997 387096 198002 387152
rect 198058 387096 200100 387152
rect 197997 387094 200100 387096
rect 197997 387091 198063 387094
rect 268009 386882 268075 386885
rect 266524 386880 268075 386882
rect 266524 386824 268014 386880
rect 268070 386824 268075 386880
rect 266524 386822 268075 386824
rect 268009 386819 268075 386822
rect 71497 385250 71563 385253
rect 71497 385248 72036 385250
rect 71497 385192 71502 385248
rect 71558 385192 72036 385248
rect 71497 385190 72036 385192
rect 71497 385187 71563 385190
rect 199193 382802 199259 382805
rect 266905 382802 266971 382805
rect 199193 382800 200100 382802
rect 199193 382744 199198 382800
rect 199254 382744 200100 382800
rect 199193 382742 200100 382744
rect 266524 382800 266971 382802
rect 266524 382744 266910 382800
rect 266966 382744 266971 382800
rect 266524 382742 266971 382744
rect 199193 382739 199259 382742
rect 266905 382739 266971 382742
rect 380893 381442 380959 381445
rect 380893 381440 384130 381442
rect 380893 381384 380898 381440
rect 380954 381384 384130 381440
rect 380893 381382 384130 381384
rect 380893 381379 380959 381382
rect 384070 381344 384130 381382
rect 583520 381156 584960 381396
rect 416865 380898 416931 380901
rect 415166 380896 416931 380898
rect 415166 380840 416870 380896
rect 416926 380840 416931 380896
rect 415166 380838 416931 380840
rect 415166 380800 415226 380838
rect 416865 380835 416931 380838
rect -960 380626 480 380716
rect 3141 380626 3207 380629
rect 129181 380626 129247 380629
rect -960 380624 3207 380626
rect -960 380568 3146 380624
rect 3202 380568 3207 380624
rect -960 380566 3207 380568
rect 126132 380624 129247 380626
rect 126132 380568 129186 380624
rect 129242 380568 129247 380624
rect 126132 380566 129247 380568
rect -960 380476 480 380566
rect 3141 380563 3207 380566
rect 129181 380563 129247 380566
rect 197905 378722 197971 378725
rect 197905 378720 200100 378722
rect 197905 378664 197910 378720
rect 197966 378664 200100 378720
rect 197905 378662 200100 378664
rect 197905 378659 197971 378662
rect 268101 378450 268167 378453
rect 266524 378448 268167 378450
rect 266524 378392 268106 378448
rect 268162 378392 268167 378448
rect 266524 378390 268167 378392
rect 268101 378387 268167 378390
rect 504725 378450 504791 378453
rect 504725 378448 504834 378450
rect 504725 378392 504730 378448
rect 504786 378392 504834 378448
rect 504725 378387 504834 378392
rect 504774 378148 504834 378387
rect 70301 377906 70367 377909
rect 71037 377906 71103 377909
rect 70301 377904 72036 377906
rect 70301 377848 70306 377904
rect 70362 377848 71042 377904
rect 71098 377848 72036 377904
rect 70301 377846 72036 377848
rect 70301 377843 70367 377846
rect 71037 377843 71103 377846
rect 380893 377226 380959 377229
rect 384070 377226 384130 377808
rect 380893 377224 384130 377226
rect 380893 377168 380898 377224
rect 380954 377168 384130 377224
rect 380893 377166 384130 377168
rect 380893 377163 380959 377166
rect 415166 376954 415226 377536
rect 417417 376954 417483 376957
rect 415166 376952 417483 376954
rect 415166 376896 417422 376952
rect 417478 376896 417483 376952
rect 415166 376894 417483 376896
rect 417417 376891 417483 376894
rect 456793 375186 456859 375189
rect 456793 375184 460092 375186
rect 456793 375128 456798 375184
rect 456854 375128 460092 375184
rect 456793 375126 460092 375128
rect 456793 375123 456859 375126
rect 416773 374642 416839 374645
rect 415166 374640 416839 374642
rect 415166 374584 416778 374640
rect 416834 374584 416839 374640
rect 415166 374582 416839 374584
rect 199285 374370 199351 374373
rect 268193 374370 268259 374373
rect 199285 374368 200100 374370
rect 199285 374312 199290 374368
rect 199346 374312 200100 374368
rect 199285 374310 200100 374312
rect 266524 374368 268259 374370
rect 266524 374312 268198 374368
rect 268254 374312 268259 374368
rect 266524 374310 268259 374312
rect 199285 374307 199351 374310
rect 268193 374307 268259 374310
rect 380893 374098 380959 374101
rect 384070 374098 384130 374544
rect 380893 374096 384130 374098
rect 380893 374040 380898 374096
rect 380954 374040 384130 374096
rect 380893 374038 384130 374040
rect 380893 374035 380959 374038
rect 415166 374000 415226 374582
rect 416773 374579 416839 374582
rect 128445 373282 128511 373285
rect 126132 373280 128511 373282
rect 126132 373224 128450 373280
rect 128506 373224 128511 373280
rect 126132 373222 128511 373224
rect 128445 373219 128511 373222
rect 128445 372738 128511 372741
rect 129273 372738 129339 372741
rect 128445 372736 129339 372738
rect 128445 372680 128450 372736
rect 128506 372680 129278 372736
rect 129334 372680 129339 372736
rect 128445 372678 129339 372680
rect 128445 372675 128511 372678
rect 129273 372675 129339 372678
rect 380893 370426 380959 370429
rect 384070 370426 384130 371008
rect 380893 370424 384130 370426
rect 380893 370368 380898 370424
rect 380954 370368 384130 370424
rect 380893 370366 384130 370368
rect 380893 370363 380959 370366
rect 70117 370290 70183 370293
rect 70301 370290 70367 370293
rect 197813 370290 197879 370293
rect 70117 370288 72036 370290
rect 70117 370232 70122 370288
rect 70178 370232 70306 370288
rect 70362 370232 72036 370288
rect 70117 370230 72036 370232
rect 197813 370288 200100 370290
rect 197813 370232 197818 370288
rect 197874 370232 200100 370288
rect 197813 370230 200100 370232
rect 70117 370227 70183 370230
rect 70301 370227 70367 370230
rect 197813 370227 197879 370230
rect 415166 370154 415226 370736
rect 416865 370154 416931 370157
rect 415166 370152 416931 370154
rect 415166 370096 416870 370152
rect 416926 370096 416931 370152
rect 415166 370094 416931 370096
rect 416865 370091 416931 370094
rect 268285 370018 268351 370021
rect 266524 370016 268351 370018
rect 266524 369960 268290 370016
rect 268346 369960 268351 370016
rect 266524 369958 268351 369960
rect 268285 369955 268351 369958
rect 580717 369610 580783 369613
rect 583520 369610 584960 369700
rect 580717 369608 584960 369610
rect 580717 369552 580722 369608
rect 580778 369552 584960 369608
rect 580717 369550 584960 369552
rect 580717 369547 580783 369550
rect 583520 369460 584960 369550
rect 381537 367434 381603 367437
rect 384070 367434 384130 367744
rect 381537 367432 384130 367434
rect 381537 367376 381542 367432
rect 381598 367376 384130 367432
rect 381537 367374 384130 367376
rect 381537 367371 381603 367374
rect 415166 367162 415226 367200
rect 416957 367162 417023 367165
rect 415166 367160 417023 367162
rect 415166 367104 416962 367160
rect 417018 367104 417023 367160
rect 415166 367102 417023 367104
rect 416957 367099 417023 367102
rect -960 366210 480 366300
rect 2957 366210 3023 366213
rect -960 366208 3023 366210
rect -960 366152 2962 366208
rect 3018 366152 3023 366208
rect -960 366150 3023 366152
rect -960 366060 480 366150
rect 2957 366147 3023 366150
rect 128905 365938 128971 365941
rect 126132 365936 128971 365938
rect 126132 365880 128910 365936
rect 128966 365880 128971 365936
rect 126132 365878 128971 365880
rect 128905 365875 128971 365878
rect 199377 365938 199443 365941
rect 268377 365938 268443 365941
rect 199377 365936 200100 365938
rect 199377 365880 199382 365936
rect 199438 365880 200100 365936
rect 199377 365878 200100 365880
rect 266524 365936 268443 365938
rect 266524 365880 268382 365936
rect 268438 365880 268443 365936
rect 266524 365878 268443 365880
rect 199377 365875 199443 365878
rect 268377 365875 268443 365878
rect 380893 363626 380959 363629
rect 384070 363626 384130 364208
rect 380893 363624 384130 363626
rect 380893 363568 380898 363624
rect 380954 363568 384130 363624
rect 380893 363566 384130 363568
rect 380893 363563 380959 363566
rect 415166 363354 415226 363936
rect 417049 363354 417115 363357
rect 415166 363352 417115 363354
rect 415166 363296 417054 363352
rect 417110 363296 417115 363352
rect 415166 363294 417115 363296
rect 417049 363291 417115 363294
rect 71589 362946 71655 362949
rect 71589 362944 72036 362946
rect 71589 362888 71594 362944
rect 71650 362888 72036 362944
rect 71589 362886 72036 362888
rect 71589 362883 71655 362886
rect 197721 361858 197787 361861
rect 197721 361856 200100 361858
rect 197721 361800 197726 361856
rect 197782 361800 200100 361856
rect 197721 361798 200100 361800
rect 197721 361795 197787 361798
rect 268469 361586 268535 361589
rect 266524 361584 268535 361586
rect 266524 361528 268474 361584
rect 268530 361528 268535 361584
rect 266524 361526 268535 361528
rect 268469 361523 268535 361526
rect 381629 360362 381695 360365
rect 384070 360362 384130 360944
rect 504774 360501 504834 361012
rect 504725 360496 504834 360501
rect 504725 360440 504730 360496
rect 504786 360440 504834 360496
rect 504725 360438 504834 360440
rect 504725 360435 504791 360438
rect 381629 360360 384130 360362
rect 381629 360304 381634 360360
rect 381690 360304 384130 360360
rect 381629 360302 384130 360304
rect 381629 360299 381695 360302
rect 415166 360226 415226 360400
rect 417141 360226 417207 360229
rect 415166 360224 417207 360226
rect 415166 360168 417146 360224
rect 417202 360168 417207 360224
rect 415166 360166 417207 360168
rect 417141 360163 417207 360166
rect 128629 358730 128695 358733
rect 126102 358728 128695 358730
rect 126102 358672 128634 358728
rect 128690 358672 128695 358728
rect 126102 358670 128695 358672
rect 126102 358292 126162 358670
rect 128629 358667 128695 358670
rect 457437 358050 457503 358053
rect 457437 358048 460092 358050
rect 457437 357992 457442 358048
rect 457498 357992 460092 358048
rect 457437 357990 460092 357992
rect 457437 357987 457503 357990
rect 580901 357914 580967 357917
rect 583520 357914 584960 358004
rect 580901 357912 584960 357914
rect 580901 357856 580906 357912
rect 580962 357856 584960 357912
rect 580901 357854 584960 357856
rect 580901 357851 580967 357854
rect 583520 357764 584960 357854
rect 197629 357506 197695 357509
rect 267089 357506 267155 357509
rect 197629 357504 200100 357506
rect 197629 357448 197634 357504
rect 197690 357448 200100 357504
rect 197629 357446 200100 357448
rect 266524 357504 267155 357506
rect 266524 357448 267094 357504
rect 267150 357448 267155 357504
rect 266524 357446 267155 357448
rect 197629 357443 197695 357446
rect 267089 357443 267155 357446
rect 381721 356826 381787 356829
rect 384070 356826 384130 357408
rect 381721 356824 384130 356826
rect 381721 356768 381726 356824
rect 381782 356768 384130 356824
rect 381721 356766 384130 356768
rect 381721 356763 381787 356766
rect 415166 356554 415226 357136
rect 417233 356554 417299 356557
rect 415166 356552 417299 356554
rect 415166 356496 417238 356552
rect 417294 356496 417299 356552
rect 415166 356494 417299 356496
rect 417233 356491 417299 356494
rect 70117 355602 70183 355605
rect 70117 355600 72036 355602
rect 70117 355544 70122 355600
rect 70178 355544 72036 355600
rect 70117 355542 72036 355544
rect 70117 355539 70183 355542
rect 380893 353562 380959 353565
rect 384070 353562 384130 354144
rect 380893 353560 384130 353562
rect 380893 353504 380898 353560
rect 380954 353504 384130 353560
rect 380893 353502 384130 353504
rect 380893 353499 380959 353502
rect 197537 353426 197603 353429
rect 268561 353426 268627 353429
rect 197537 353424 200100 353426
rect 197537 353368 197542 353424
rect 197598 353368 200100 353424
rect 197537 353366 200100 353368
rect 266524 353424 268627 353426
rect 266524 353368 268566 353424
rect 268622 353368 268627 353424
rect 266524 353366 268627 353368
rect 415166 353426 415226 353600
rect 417325 353426 417391 353429
rect 415166 353424 417391 353426
rect 415166 353368 417330 353424
rect 417386 353368 417391 353424
rect 415166 353366 417391 353368
rect 197537 353363 197603 353366
rect 268561 353363 268627 353366
rect 417325 353363 417391 353366
rect -960 351780 480 352020
rect 129733 350978 129799 350981
rect 126132 350976 129799 350978
rect 126132 350920 129738 350976
rect 129794 350920 129799 350976
rect 126132 350918 129799 350920
rect 129733 350915 129799 350918
rect 197445 349074 197511 349077
rect 267181 349074 267247 349077
rect 197445 349072 200100 349074
rect 197445 349016 197450 349072
rect 197506 349016 200100 349072
rect 197445 349014 200100 349016
rect 266524 349072 267247 349074
rect 266524 349016 267186 349072
rect 267242 349016 267247 349072
rect 266524 349014 267247 349016
rect 197445 349011 197511 349014
rect 267181 349011 267247 349014
rect 70209 348258 70275 348261
rect 71589 348258 71655 348261
rect 70209 348256 72036 348258
rect 70209 348200 70214 348256
rect 70270 348200 71594 348256
rect 71650 348200 72036 348256
rect 70209 348198 72036 348200
rect 70209 348195 70275 348198
rect 71589 348195 71655 348198
rect 579981 346082 580047 346085
rect 583520 346082 584960 346172
rect 579981 346080 584960 346082
rect 579981 346024 579986 346080
rect 580042 346024 584960 346080
rect 579981 346022 584960 346024
rect 579981 346019 580047 346022
rect 583520 345932 584960 346022
rect 199469 344994 199535 344997
rect 268653 344994 268719 344997
rect 199469 344992 200100 344994
rect 199469 344936 199474 344992
rect 199530 344936 200100 344992
rect 199469 344934 200100 344936
rect 266524 344992 268719 344994
rect 266524 344936 268658 344992
rect 268714 344936 268719 344992
rect 266524 344934 268719 344936
rect 199469 344931 199535 344934
rect 268653 344931 268719 344934
rect 504774 343637 504834 343876
rect 128813 343634 128879 343637
rect 126132 343632 128879 343634
rect 126132 343576 128818 343632
rect 128874 343576 128879 343632
rect 126132 343574 128879 343576
rect 128813 343571 128879 343574
rect 504725 343632 504834 343637
rect 504725 343576 504730 343632
rect 504786 343576 504834 343632
rect 504725 343574 504834 343576
rect 504725 343571 504791 343574
rect 70117 341458 70183 341461
rect 134333 341458 134399 341461
rect 185577 341458 185643 341461
rect 70117 341456 185643 341458
rect 70117 341400 70122 341456
rect 70178 341400 134338 341456
rect 134394 341400 185582 341456
rect 185638 341400 185643 341456
rect 70117 341398 185643 341400
rect 70117 341395 70183 341398
rect 134333 341395 134399 341398
rect 185577 341395 185643 341398
rect 503713 340914 503779 340917
rect 503897 340914 503963 340917
rect 503713 340912 503963 340914
rect 503713 340856 503718 340912
rect 503774 340856 503902 340912
rect 503958 340856 503963 340912
rect 503713 340854 503963 340856
rect 503713 340851 503779 340854
rect 503897 340851 503963 340854
rect 154573 340506 154639 340509
rect 157333 340506 157399 340509
rect 154573 340504 157399 340506
rect 154573 340448 154578 340504
rect 154634 340448 157338 340504
rect 157394 340448 157399 340504
rect 154573 340446 157399 340448
rect 154573 340443 154639 340446
rect 157333 340443 157399 340446
rect 240133 340506 240199 340509
rect 249701 340506 249767 340509
rect 240133 340504 249767 340506
rect 240133 340448 240138 340504
rect 240194 340448 249706 340504
rect 249762 340448 249767 340504
rect 240133 340446 249767 340448
rect 240133 340443 240199 340446
rect 249701 340443 249767 340446
rect 259453 340506 259519 340509
rect 268929 340506 268995 340509
rect 259453 340504 268995 340506
rect 259453 340448 259458 340504
rect 259514 340448 268934 340504
rect 268990 340448 268995 340504
rect 259453 340446 268995 340448
rect 259453 340443 259519 340446
rect 268929 340443 268995 340446
rect 269113 340506 269179 340509
rect 273253 340506 273319 340509
rect 269113 340504 273319 340506
rect 269113 340448 269118 340504
rect 269174 340448 273258 340504
rect 273314 340448 273319 340504
rect 269113 340446 273319 340448
rect 269113 340443 269179 340446
rect 273253 340443 273319 340446
rect 193213 340370 193279 340373
rect 202781 340370 202847 340373
rect 193213 340368 202847 340370
rect 193213 340312 193218 340368
rect 193274 340312 202786 340368
rect 202842 340312 202847 340368
rect 193213 340310 202847 340312
rect 193213 340307 193279 340310
rect 202781 340307 202847 340310
rect 230473 340370 230539 340373
rect 240041 340370 240107 340373
rect 230473 340368 240107 340370
rect 230473 340312 230478 340368
rect 230534 340312 240046 340368
rect 240102 340312 240107 340368
rect 230473 340310 240107 340312
rect 230473 340307 230539 340310
rect 240041 340307 240107 340310
rect -960 337514 480 337604
rect 2957 337514 3023 337517
rect -960 337512 3023 337514
rect -960 337456 2962 337512
rect 3018 337456 3023 337512
rect -960 337454 3023 337456
rect -960 337364 480 337454
rect 2957 337451 3023 337454
rect 128353 335338 128419 335341
rect 128537 335338 128603 335341
rect 128353 335336 128603 335338
rect 128353 335280 128358 335336
rect 128414 335280 128542 335336
rect 128598 335280 128603 335336
rect 128353 335278 128603 335280
rect 128353 335275 128419 335278
rect 128537 335275 128603 335278
rect 583520 334236 584960 334476
rect 258165 327042 258231 327045
rect 258349 327042 258415 327045
rect 258165 327040 258415 327042
rect 258165 326984 258170 327040
rect 258226 326984 258354 327040
rect 258410 326984 258415 327040
rect 258165 326982 258415 326984
rect 258165 326979 258231 326982
rect 258349 326979 258415 326982
rect -960 323098 480 323188
rect 2957 323098 3023 323101
rect -960 323096 3023 323098
rect -960 323040 2962 323096
rect 3018 323040 3023 323096
rect -960 323038 3023 323040
rect -960 322948 480 323038
rect 2957 323035 3023 323038
rect 580165 322690 580231 322693
rect 583520 322690 584960 322780
rect 580165 322688 584960 322690
rect 580165 322632 580170 322688
rect 580226 322632 584960 322688
rect 580165 322630 584960 322632
rect 580165 322627 580231 322630
rect 583520 322540 584960 322630
rect 503897 321738 503963 321741
rect 503854 321736 503963 321738
rect 503854 321680 503902 321736
rect 503958 321680 503963 321736
rect 503854 321675 503963 321680
rect 503854 321469 503914 321675
rect 503854 321464 503963 321469
rect 503854 321408 503902 321464
rect 503958 321408 503963 321464
rect 503854 321406 503963 321408
rect 503897 321403 503963 321406
rect 580165 310858 580231 310861
rect 583520 310858 584960 310948
rect 580165 310856 584960 310858
rect 580165 310800 580170 310856
rect 580226 310800 584960 310856
rect 580165 310798 584960 310800
rect 580165 310795 580231 310798
rect 583520 310708 584960 310798
rect 255589 309226 255655 309229
rect 255865 309226 255931 309229
rect 255589 309224 255931 309226
rect 255589 309168 255594 309224
rect 255650 309168 255870 309224
rect 255926 309168 255931 309224
rect 255589 309166 255931 309168
rect 255589 309163 255655 309166
rect 255865 309163 255931 309166
rect 258349 309226 258415 309229
rect 258625 309226 258691 309229
rect 258349 309224 258691 309226
rect 258349 309168 258354 309224
rect 258410 309168 258630 309224
rect 258686 309168 258691 309224
rect 258349 309166 258691 309168
rect 258349 309163 258415 309166
rect 258625 309163 258691 309166
rect -960 308818 480 308908
rect 2957 308818 3023 308821
rect -960 308816 3023 308818
rect -960 308760 2962 308816
rect 3018 308760 3023 308816
rect -960 308758 3023 308760
rect -960 308668 480 308758
rect 2957 308755 3023 308758
rect 580809 299162 580875 299165
rect 583520 299162 584960 299252
rect 580809 299160 584960 299162
rect 580809 299104 580814 299160
rect 580870 299104 584960 299160
rect 580809 299102 584960 299104
rect 580809 299099 580875 299102
rect 583520 299012 584960 299102
rect -960 294402 480 294492
rect 2957 294402 3023 294405
rect -960 294400 3023 294402
rect -960 294344 2962 294400
rect 3018 294344 3023 294400
rect -960 294342 3023 294344
rect -960 294252 480 294342
rect 2957 294339 3023 294342
rect 271965 294130 272031 294133
rect 271830 294128 272031 294130
rect 271830 294072 271970 294128
rect 272026 294072 272031 294128
rect 271830 294070 272031 294072
rect 271830 293997 271890 294070
rect 271965 294067 272031 294070
rect 271781 293992 271890 293997
rect 271781 293936 271786 293992
rect 271842 293936 271890 293992
rect 271781 293934 271890 293936
rect 271781 293931 271847 293934
rect 583520 287316 584960 287556
rect -960 280122 480 280212
rect 2957 280122 3023 280125
rect -960 280120 3023 280122
rect -960 280064 2962 280120
rect 3018 280064 3023 280120
rect -960 280062 3023 280064
rect -960 279972 480 280062
rect 2957 280059 3023 280062
rect 579981 275770 580047 275773
rect 583520 275770 584960 275860
rect 579981 275768 584960 275770
rect 579981 275712 579986 275768
rect 580042 275712 584960 275768
rect 579981 275710 584960 275712
rect 579981 275707 580047 275710
rect 583520 275620 584960 275710
rect 271965 274818 272031 274821
rect 271830 274816 272031 274818
rect 271830 274760 271970 274816
rect 272026 274760 272031 274816
rect 271830 274758 272031 274760
rect 271830 274685 271890 274758
rect 271965 274755 272031 274758
rect 271781 274680 271890 274685
rect 271781 274624 271786 274680
rect 271842 274624 271890 274680
rect 271781 274622 271890 274624
rect 271781 274619 271847 274622
rect -960 265706 480 265796
rect 2865 265706 2931 265709
rect -960 265704 2931 265706
rect -960 265648 2870 265704
rect 2926 265648 2931 265704
rect -960 265646 2931 265648
rect -960 265556 480 265646
rect 2865 265643 2931 265646
rect 580165 263938 580231 263941
rect 583520 263938 584960 264028
rect 580165 263936 584960 263938
rect 580165 263880 580170 263936
rect 580226 263880 584960 263936
rect 580165 263878 584960 263880
rect 580165 263875 580231 263878
rect 583520 263788 584960 263878
rect 504265 260946 504331 260949
rect 504541 260946 504607 260949
rect 504265 260944 504607 260946
rect 504265 260888 504270 260944
rect 504326 260888 504546 260944
rect 504602 260888 504607 260944
rect 504265 260886 504607 260888
rect 504265 260883 504331 260886
rect 504541 260883 504607 260886
rect 281165 260812 281231 260813
rect 281165 260810 281212 260812
rect 281120 260808 281212 260810
rect 281120 260752 281170 260808
rect 281120 260750 281212 260752
rect 281165 260748 281212 260750
rect 281276 260748 281282 260812
rect 281165 260747 281231 260748
rect 271597 255370 271663 255373
rect 271781 255370 271847 255373
rect 271597 255368 271847 255370
rect 271597 255312 271602 255368
rect 271658 255312 271786 255368
rect 271842 255312 271847 255368
rect 271597 255310 271847 255312
rect 271597 255307 271663 255310
rect 271781 255307 271847 255310
rect 580165 252242 580231 252245
rect 583520 252242 584960 252332
rect 580165 252240 584960 252242
rect 580165 252184 580170 252240
rect 580226 252184 584960 252240
rect 580165 252182 584960 252184
rect 580165 252179 580231 252182
rect 583520 252092 584960 252182
rect 308857 251426 308923 251429
rect 308857 251424 309058 251426
rect -960 251290 480 251380
rect 308857 251368 308862 251424
rect 308918 251368 309058 251424
rect 308857 251366 309058 251368
rect 308857 251363 308923 251366
rect 2865 251290 2931 251293
rect -960 251288 2931 251290
rect -960 251232 2870 251288
rect 2926 251232 2931 251288
rect -960 251230 2931 251232
rect -960 251140 480 251230
rect 2865 251227 2931 251230
rect 128077 251290 128143 251293
rect 128445 251290 128511 251293
rect 128077 251288 128511 251290
rect 128077 251232 128082 251288
rect 128138 251232 128450 251288
rect 128506 251232 128511 251288
rect 128077 251230 128511 251232
rect 128077 251227 128143 251230
rect 128445 251227 128511 251230
rect 281206 251228 281212 251292
rect 281276 251228 281282 251292
rect 308857 251290 308923 251293
rect 308998 251290 309058 251366
rect 308857 251288 309058 251290
rect 308857 251232 308862 251288
rect 308918 251232 309058 251288
rect 308857 251230 309058 251232
rect 281073 251154 281139 251157
rect 281214 251154 281274 251228
rect 308857 251227 308923 251230
rect 281073 251152 281274 251154
rect 281073 251096 281078 251152
rect 281134 251096 281274 251152
rect 281073 251094 281274 251096
rect 281073 251091 281139 251094
rect 132861 241498 132927 241501
rect 133505 241498 133571 241501
rect 132861 241496 133571 241498
rect 132861 241440 132866 241496
rect 132922 241440 133510 241496
rect 133566 241440 133571 241496
rect 132861 241438 133571 241440
rect 132861 241435 132927 241438
rect 133505 241435 133571 241438
rect 257981 241498 258047 241501
rect 258165 241498 258231 241501
rect 257981 241496 258231 241498
rect 257981 241440 257986 241496
rect 258042 241440 258170 241496
rect 258226 241440 258231 241496
rect 257981 241438 258231 241440
rect 257981 241435 258047 241438
rect 258165 241435 258231 241438
rect 583520 240396 584960 240636
rect -960 237010 480 237100
rect 2865 237010 2931 237013
rect -960 237008 2931 237010
rect -960 236952 2870 237008
rect 2926 236952 2931 237008
rect -960 236950 2931 236952
rect -960 236860 480 236950
rect 2865 236947 2931 236950
rect 580073 228850 580139 228853
rect 583520 228850 584960 228940
rect 580073 228848 584960 228850
rect 580073 228792 580078 228848
rect 580134 228792 584960 228848
rect 580073 228790 584960 228792
rect 580073 228787 580139 228790
rect 583520 228700 584960 228790
rect -960 222594 480 222684
rect 2773 222594 2839 222597
rect -960 222592 2839 222594
rect -960 222536 2778 222592
rect 2834 222536 2839 222592
rect -960 222534 2839 222536
rect -960 222444 480 222534
rect 2773 222531 2839 222534
rect 579797 217018 579863 217021
rect 583520 217018 584960 217108
rect 579797 217016 584960 217018
rect 579797 216960 579802 217016
rect 579858 216960 584960 217016
rect 579797 216958 584960 216960
rect 579797 216955 579863 216958
rect 583520 216868 584960 216958
rect 122649 212530 122715 212533
rect 122833 212530 122899 212533
rect 122649 212528 122899 212530
rect 122649 212472 122654 212528
rect 122710 212472 122838 212528
rect 122894 212472 122899 212528
rect 122649 212470 122899 212472
rect 122649 212467 122715 212470
rect 122833 212467 122899 212470
rect 128445 212530 128511 212533
rect 128629 212530 128695 212533
rect 128445 212528 128695 212530
rect 128445 212472 128450 212528
rect 128506 212472 128634 212528
rect 128690 212472 128695 212528
rect 128445 212470 128695 212472
rect 128445 212467 128511 212470
rect 128629 212467 128695 212470
rect -960 208178 480 208268
rect 3049 208178 3115 208181
rect -960 208176 3115 208178
rect -960 208120 3054 208176
rect 3110 208120 3115 208176
rect -960 208118 3115 208120
rect -960 208028 480 208118
rect 3049 208115 3115 208118
rect 580073 205322 580139 205325
rect 583520 205322 584960 205412
rect 580073 205320 584960 205322
rect 580073 205264 580078 205320
rect 580134 205264 584960 205320
rect 580073 205262 584960 205264
rect 580073 205259 580139 205262
rect 583520 205172 584960 205262
rect 122649 202874 122715 202877
rect 122925 202874 122991 202877
rect 122649 202872 122991 202874
rect 122649 202816 122654 202872
rect 122710 202816 122930 202872
rect 122986 202816 122991 202872
rect 122649 202814 122991 202816
rect 122649 202811 122715 202814
rect 122925 202811 122991 202814
rect 197261 202874 197327 202877
rect 220353 202874 220419 202877
rect 197261 202872 220419 202874
rect 197261 202816 197266 202872
rect 197322 202816 220358 202872
rect 220414 202816 220419 202872
rect 197261 202814 220419 202816
rect 197261 202811 197327 202814
rect 220353 202811 220419 202814
rect 195697 202738 195763 202741
rect 223849 202738 223915 202741
rect 195697 202736 223915 202738
rect 195697 202680 195702 202736
rect 195758 202680 223854 202736
rect 223910 202680 223915 202736
rect 195697 202678 223915 202680
rect 195697 202675 195763 202678
rect 223849 202675 223915 202678
rect 195789 202602 195855 202605
rect 226333 202602 226399 202605
rect 195789 202600 226399 202602
rect 195789 202544 195794 202600
rect 195850 202544 226338 202600
rect 226394 202544 226399 202600
rect 195789 202542 226399 202544
rect 195789 202539 195855 202542
rect 226333 202539 226399 202542
rect 302233 202602 302299 202605
rect 307201 202602 307267 202605
rect 302233 202600 307267 202602
rect 302233 202544 302238 202600
rect 302294 202544 307206 202600
rect 307262 202544 307267 202600
rect 302233 202542 307267 202544
rect 302233 202539 302299 202542
rect 307201 202539 307267 202542
rect 197169 202466 197235 202469
rect 228633 202466 228699 202469
rect 197169 202464 228699 202466
rect 197169 202408 197174 202464
rect 197230 202408 228638 202464
rect 228694 202408 228699 202464
rect 197169 202406 228699 202408
rect 197169 202403 197235 202406
rect 228633 202403 228699 202406
rect 252645 202466 252711 202469
rect 254117 202466 254183 202469
rect 252645 202464 254183 202466
rect 252645 202408 252650 202464
rect 252706 202408 254122 202464
rect 254178 202408 254183 202464
rect 252645 202406 254183 202408
rect 252645 202403 252711 202406
rect 254117 202403 254183 202406
rect 197077 202330 197143 202333
rect 233417 202330 233483 202333
rect 197077 202328 233483 202330
rect 197077 202272 197082 202328
rect 197138 202272 233422 202328
rect 233478 202272 233483 202328
rect 197077 202270 233483 202272
rect 197077 202267 197143 202270
rect 233417 202267 233483 202270
rect 253473 202330 253539 202333
rect 253933 202330 253999 202333
rect 253473 202328 253999 202330
rect 253473 202272 253478 202328
rect 253534 202272 253938 202328
rect 253994 202272 253999 202328
rect 253473 202270 253999 202272
rect 253473 202267 253539 202270
rect 253933 202267 253999 202270
rect 258533 202330 258599 202333
rect 259453 202330 259519 202333
rect 258533 202328 259519 202330
rect 258533 202272 258538 202328
rect 258594 202272 259458 202328
rect 259514 202272 259519 202328
rect 258533 202270 259519 202272
rect 258533 202267 258599 202270
rect 259453 202267 259519 202270
rect 199009 202194 199075 202197
rect 261937 202194 262003 202197
rect 199009 202192 262003 202194
rect 199009 202136 199014 202192
rect 199070 202136 261942 202192
rect 261998 202136 262003 202192
rect 199009 202134 262003 202136
rect 199009 202131 199075 202134
rect 261937 202131 262003 202134
rect 277301 202194 277367 202197
rect 378409 202194 378475 202197
rect 277301 202192 378475 202194
rect 277301 202136 277306 202192
rect 277362 202136 378414 202192
rect 378470 202136 378475 202192
rect 277301 202134 378475 202136
rect 277301 202131 277367 202134
rect 378409 202131 378475 202134
rect 198641 202058 198707 202061
rect 213453 202058 213519 202061
rect 198641 202056 213519 202058
rect 198641 202000 198646 202056
rect 198702 202000 213458 202056
rect 213514 202000 213519 202056
rect 198641 201998 213519 202000
rect 198641 201995 198707 201998
rect 213453 201995 213519 201998
rect 304257 202058 304323 202061
rect 307293 202058 307359 202061
rect 304257 202056 307359 202058
rect 304257 202000 304262 202056
rect 304318 202000 307298 202056
rect 307354 202000 307359 202056
rect 304257 201998 307359 202000
rect 304257 201995 304323 201998
rect 307293 201995 307359 201998
rect 133086 200092 133092 200156
rect 133156 200154 133162 200156
rect 134333 200154 134399 200157
rect 133156 200152 134399 200154
rect 133156 200096 134338 200152
rect 134394 200096 134399 200152
rect 133156 200094 134399 200096
rect 133156 200092 133162 200094
rect 134333 200091 134399 200094
rect 131205 199338 131271 199341
rect 131205 199336 134044 199338
rect 131205 199280 131210 199336
rect 131266 199280 134044 199336
rect 131205 199278 134044 199280
rect 131205 199275 131271 199278
rect 436829 198930 436895 198933
rect 433934 198928 436895 198930
rect 433934 198872 436834 198928
rect 436890 198872 436895 198928
rect 433934 198870 436895 198872
rect 433934 198764 433994 198870
rect 436829 198867 436895 198870
rect 131205 198250 131271 198253
rect 131205 198248 134044 198250
rect 131205 198192 131210 198248
rect 131266 198192 134044 198248
rect 131205 198190 134044 198192
rect 131205 198187 131271 198190
rect 131297 197162 131363 197165
rect 131297 197160 134044 197162
rect 131297 197104 131302 197160
rect 131358 197104 134044 197160
rect 131297 197102 134044 197104
rect 131297 197099 131363 197102
rect 433934 196210 433994 196724
rect 436369 196210 436435 196213
rect 131254 196150 134044 196210
rect 433934 196208 436435 196210
rect 433934 196152 436374 196208
rect 436430 196152 436435 196208
rect 433934 196150 436435 196152
rect 131254 196077 131314 196150
rect 436369 196147 436435 196150
rect 131205 196072 131314 196077
rect 132861 196076 132927 196077
rect 132861 196074 132908 196076
rect 131205 196016 131210 196072
rect 131266 196016 131314 196072
rect 131205 196014 131314 196016
rect 132816 196072 132908 196074
rect 132816 196016 132866 196072
rect 132816 196014 132908 196016
rect 131205 196011 131271 196014
rect 132861 196012 132908 196014
rect 132972 196012 132978 196076
rect 132861 196011 132927 196012
rect 132861 195940 132927 195941
rect 132861 195938 132908 195940
rect 132816 195936 132908 195938
rect 132816 195880 132866 195936
rect 132816 195878 132908 195880
rect 132861 195876 132908 195878
rect 132972 195876 132978 195940
rect 132861 195875 132927 195876
rect 131205 195122 131271 195125
rect 131205 195120 134044 195122
rect 131205 195064 131210 195120
rect 131266 195064 134044 195120
rect 131205 195062 134044 195064
rect 131205 195059 131271 195062
rect 131205 194034 131271 194037
rect 433934 194034 433994 194548
rect 436461 194034 436527 194037
rect 131205 194032 134044 194034
rect -960 193898 480 193988
rect 131205 193976 131210 194032
rect 131266 193976 134044 194032
rect 131205 193974 134044 193976
rect 433934 194032 436527 194034
rect 433934 193976 436466 194032
rect 436522 193976 436527 194032
rect 433934 193974 436527 193976
rect 131205 193971 131271 193974
rect 436461 193971 436527 193974
rect 3049 193898 3115 193901
rect -960 193896 3115 193898
rect -960 193840 3054 193896
rect 3110 193840 3115 193896
rect -960 193838 3115 193840
rect -960 193748 480 193838
rect 3049 193835 3115 193838
rect 583520 193476 584960 193716
rect 8017 193218 8083 193221
rect 8293 193218 8359 193221
rect 8017 193216 8359 193218
rect 8017 193160 8022 193216
rect 8078 193160 8298 193216
rect 8354 193160 8359 193216
rect 8017 193158 8359 193160
rect 8017 193155 8083 193158
rect 8293 193155 8359 193158
rect 128353 193218 128419 193221
rect 128537 193218 128603 193221
rect 128353 193216 128603 193218
rect 128353 193160 128358 193216
rect 128414 193160 128542 193216
rect 128598 193160 128603 193216
rect 128353 193158 128603 193160
rect 128353 193155 128419 193158
rect 128537 193155 128603 193158
rect 436277 193082 436343 193085
rect 433934 193080 436343 193082
rect 433934 193024 436282 193080
rect 436338 193024 436343 193080
rect 433934 193022 436343 193024
rect 131205 192946 131271 192949
rect 131205 192944 134044 192946
rect 131205 192888 131210 192944
rect 131266 192888 134044 192944
rect 131205 192886 134044 192888
rect 131205 192883 131271 192886
rect 433934 192508 433994 193022
rect 436277 193019 436343 193022
rect 131205 191994 131271 191997
rect 131205 191992 134044 191994
rect 131205 191936 131210 191992
rect 131266 191936 134044 191992
rect 131205 191934 134044 191936
rect 131205 191931 131271 191934
rect 131205 190906 131271 190909
rect 131205 190904 134044 190906
rect 131205 190848 131210 190904
rect 131266 190848 134044 190904
rect 131205 190846 134044 190848
rect 131205 190843 131271 190846
rect 433934 190226 433994 190332
rect 434989 190226 435055 190229
rect 433934 190224 435055 190226
rect 433934 190168 434994 190224
rect 435050 190168 435055 190224
rect 433934 190166 435055 190168
rect 434989 190163 435055 190166
rect 131205 189818 131271 189821
rect 131205 189816 134044 189818
rect 131205 189760 131210 189816
rect 131266 189760 134044 189816
rect 131205 189758 134044 189760
rect 131205 189755 131271 189758
rect 9673 189002 9739 189005
rect 19241 189002 19307 189005
rect 9673 189000 19307 189002
rect 9673 188944 9678 189000
rect 9734 188944 19246 189000
rect 19302 188944 19307 189000
rect 9673 188942 19307 188944
rect 9673 188939 9739 188942
rect 19241 188939 19307 188942
rect 67633 188866 67699 188869
rect 77201 188866 77267 188869
rect 67633 188864 77267 188866
rect 67633 188808 67638 188864
rect 67694 188808 77206 188864
rect 77262 188808 77267 188864
rect 67633 188806 77267 188808
rect 67633 188803 67699 188806
rect 77201 188803 77267 188806
rect 86953 188866 87019 188869
rect 96337 188866 96403 188869
rect 86953 188864 96403 188866
rect 86953 188808 86958 188864
rect 87014 188808 96342 188864
rect 96398 188808 96403 188864
rect 86953 188806 96403 188808
rect 86953 188803 87019 188806
rect 96337 188803 96403 188806
rect 115933 188866 115999 188869
rect 125501 188866 125567 188869
rect 434897 188866 434963 188869
rect 115933 188864 125567 188866
rect 115933 188808 115938 188864
rect 115994 188808 125506 188864
rect 125562 188808 125567 188864
rect 115933 188806 125567 188808
rect 115933 188803 115999 188806
rect 125501 188803 125567 188806
rect 433934 188864 434963 188866
rect 433934 188808 434902 188864
rect 434958 188808 434963 188864
rect 433934 188806 434963 188808
rect 131205 188730 131271 188733
rect 131205 188728 134044 188730
rect 131205 188672 131210 188728
rect 131266 188672 134044 188728
rect 131205 188670 134044 188672
rect 131205 188667 131271 188670
rect 433934 188292 433994 188806
rect 434897 188803 434963 188806
rect 131205 187778 131271 187781
rect 131205 187776 134044 187778
rect 131205 187720 131210 187776
rect 131266 187720 134044 187776
rect 131205 187718 134044 187720
rect 131205 187715 131271 187718
rect 131205 186690 131271 186693
rect 131205 186688 134044 186690
rect 131205 186632 131210 186688
rect 131266 186632 134044 186688
rect 131205 186630 134044 186632
rect 131205 186627 131271 186630
rect 434805 186282 434871 186285
rect 433934 186280 434871 186282
rect 433934 186224 434810 186280
rect 434866 186224 434871 186280
rect 433934 186222 434871 186224
rect 433934 186116 433994 186222
rect 434805 186219 434871 186222
rect 131205 185602 131271 185605
rect 131205 185600 134044 185602
rect 131205 185544 131210 185600
rect 131266 185544 134044 185600
rect 131205 185542 134044 185544
rect 131205 185539 131271 185542
rect 132902 185404 132908 185468
rect 132972 185466 132978 185468
rect 133229 185466 133295 185469
rect 132972 185464 133295 185466
rect 132972 185408 133234 185464
rect 133290 185408 133295 185464
rect 132972 185406 133295 185408
rect 132972 185404 132978 185406
rect 133229 185403 133295 185406
rect 133045 184924 133111 184925
rect 133045 184922 133092 184924
rect 133000 184920 133092 184922
rect 133000 184864 133050 184920
rect 133000 184862 133092 184864
rect 133045 184860 133092 184862
rect 133156 184860 133162 184924
rect 133045 184859 133111 184860
rect 434713 184650 434779 184653
rect 433934 184648 434779 184650
rect 433934 184592 434718 184648
rect 434774 184592 434779 184648
rect 433934 184590 434779 184592
rect 131205 184514 131271 184517
rect 131205 184512 134044 184514
rect 131205 184456 131210 184512
rect 131266 184456 134044 184512
rect 131205 184454 134044 184456
rect 131205 184451 131271 184454
rect 433934 184076 433994 184590
rect 434713 184587 434779 184590
rect 131205 183562 131271 183565
rect 504357 183562 504423 183565
rect 504633 183562 504699 183565
rect 131205 183560 134044 183562
rect 131205 183504 131210 183560
rect 131266 183504 134044 183560
rect 131205 183502 134044 183504
rect 504357 183560 504699 183562
rect 504357 183504 504362 183560
rect 504418 183504 504638 183560
rect 504694 183504 504699 183560
rect 504357 183502 504699 183504
rect 131205 183499 131271 183502
rect 504357 183499 504423 183502
rect 504633 183499 504699 183502
rect 132861 182474 132927 182477
rect 132861 182472 134044 182474
rect 132861 182416 132866 182472
rect 132922 182416 134044 182472
rect 132861 182414 134044 182416
rect 132861 182411 132927 182414
rect 132861 182340 132927 182341
rect 132861 182336 132908 182340
rect 132972 182338 132978 182340
rect 132861 182280 132866 182336
rect 132861 182276 132908 182280
rect 132972 182278 133018 182338
rect 132972 182276 132978 182278
rect 132861 182275 132927 182276
rect 436737 182066 436803 182069
rect 433934 182064 436803 182066
rect 433934 182008 436742 182064
rect 436798 182008 436803 182064
rect 433934 182006 436803 182008
rect 433934 181900 433994 182006
rect 436737 182003 436803 182006
rect 579981 181930 580047 181933
rect 583520 181930 584960 182020
rect 579981 181928 584960 181930
rect 579981 181872 579986 181928
rect 580042 181872 584960 181928
rect 579981 181870 584960 181872
rect 579981 181867 580047 181870
rect 583520 181780 584960 181870
rect 133229 181386 133295 181389
rect 133229 181384 134044 181386
rect 133229 181328 133234 181384
rect 133290 181328 134044 181384
rect 133229 181326 134044 181328
rect 133229 181323 133295 181326
rect 132033 180434 132099 180437
rect 132033 180432 134044 180434
rect 132033 180376 132038 180432
rect 132094 180376 134044 180432
rect 132033 180374 134044 180376
rect 132033 180371 132099 180374
rect 436185 180298 436251 180301
rect 433934 180296 436251 180298
rect 433934 180240 436190 180296
rect 436246 180240 436251 180296
rect 433934 180238 436251 180240
rect 433934 179860 433994 180238
rect 436185 180235 436251 180238
rect -960 179482 480 179572
rect 3693 179482 3759 179485
rect -960 179480 3759 179482
rect -960 179424 3698 179480
rect 3754 179424 3759 179480
rect -960 179422 3759 179424
rect -960 179332 480 179422
rect 3693 179419 3759 179422
rect 133321 179346 133387 179349
rect 133321 179344 134044 179346
rect 133321 179288 133326 179344
rect 133382 179288 134044 179344
rect 133321 179286 134044 179288
rect 133321 179283 133387 179286
rect 132861 178258 132927 178261
rect 132861 178256 134044 178258
rect 132861 178200 132866 178256
rect 132922 178200 134044 178256
rect 132861 178198 134044 178200
rect 132861 178195 132927 178198
rect 436645 177986 436711 177989
rect 433934 177984 436711 177986
rect 433934 177928 436650 177984
rect 436706 177928 436711 177984
rect 433934 177926 436711 177928
rect 433934 177684 433994 177926
rect 436645 177923 436711 177926
rect 133413 177170 133479 177173
rect 133413 177168 134044 177170
rect 133413 177112 133418 177168
rect 133474 177112 134044 177168
rect 133413 177110 134044 177112
rect 133413 177107 133479 177110
rect 133229 176218 133295 176221
rect 436553 176218 436619 176221
rect 133229 176216 134044 176218
rect 133229 176160 133234 176216
rect 133290 176160 134044 176216
rect 133229 176158 134044 176160
rect 433934 176216 436619 176218
rect 433934 176160 436558 176216
rect 436614 176160 436619 176216
rect 433934 176158 436619 176160
rect 133229 176155 133295 176158
rect 433934 175644 433994 176158
rect 436553 176155 436619 176158
rect 131205 175130 131271 175133
rect 131205 175128 134044 175130
rect 131205 175072 131210 175128
rect 131266 175072 134044 175128
rect 131205 175070 134044 175072
rect 131205 175067 131271 175070
rect 132033 174042 132099 174045
rect 132033 174040 134044 174042
rect 132033 173984 132038 174040
rect 132094 173984 134044 174040
rect 132033 173982 134044 173984
rect 132033 173979 132099 173982
rect 434253 173906 434319 173909
rect 433934 173904 434319 173906
rect 433934 173848 434258 173904
rect 434314 173848 434319 173904
rect 433934 173846 434319 173848
rect 433934 173468 433994 173846
rect 434253 173843 434319 173846
rect 130929 172954 130995 172957
rect 130929 172952 134044 172954
rect 130929 172896 130934 172952
rect 130990 172896 134044 172952
rect 130929 172894 134044 172896
rect 130929 172891 130995 172894
rect 130653 172002 130719 172005
rect 434529 172002 434595 172005
rect 130653 172000 134044 172002
rect 130653 171944 130658 172000
rect 130714 171944 134044 172000
rect 130653 171942 134044 171944
rect 433934 172000 434595 172002
rect 433934 171944 434534 172000
rect 434590 171944 434595 172000
rect 433934 171942 434595 171944
rect 130653 171939 130719 171942
rect 433934 171428 433994 171942
rect 434529 171939 434595 171942
rect 130745 170914 130811 170917
rect 130745 170912 134044 170914
rect 130745 170856 130750 170912
rect 130806 170856 134044 170912
rect 130745 170854 134044 170856
rect 130745 170851 130811 170854
rect 580349 170098 580415 170101
rect 583520 170098 584960 170188
rect 580349 170096 584960 170098
rect 580349 170040 580354 170096
rect 580410 170040 584960 170096
rect 580349 170038 584960 170040
rect 580349 170035 580415 170038
rect 583520 169948 584960 170038
rect 130561 169826 130627 169829
rect 130561 169824 134044 169826
rect 130561 169768 130566 169824
rect 130622 169768 134044 169824
rect 130561 169766 134044 169768
rect 130561 169763 130627 169766
rect 434437 169690 434503 169693
rect 433934 169688 434503 169690
rect 433934 169632 434442 169688
rect 434498 169632 434503 169688
rect 433934 169630 434503 169632
rect 433934 169252 433994 169630
rect 434437 169627 434503 169630
rect 132953 168738 133019 168741
rect 132953 168736 134044 168738
rect 132953 168680 132958 168736
rect 133014 168680 134044 168736
rect 132953 168678 134044 168680
rect 132953 168675 133019 168678
rect 132401 167786 132467 167789
rect 434345 167786 434411 167789
rect 132401 167784 134044 167786
rect 132401 167728 132406 167784
rect 132462 167728 134044 167784
rect 132401 167726 134044 167728
rect 433934 167784 434411 167786
rect 433934 167728 434350 167784
rect 434406 167728 434411 167784
rect 433934 167726 434411 167728
rect 132401 167723 132467 167726
rect 433934 167212 433994 167726
rect 434345 167723 434411 167726
rect 132033 166698 132099 166701
rect 132033 166696 134044 166698
rect 132033 166640 132038 166696
rect 132094 166640 134044 166696
rect 132033 166638 134044 166640
rect 132033 166635 132099 166638
rect 131573 165610 131639 165613
rect 434161 165610 434227 165613
rect 131573 165608 134044 165610
rect 131573 165552 131578 165608
rect 131634 165552 134044 165608
rect 131573 165550 134044 165552
rect 433934 165608 434227 165610
rect 433934 165552 434166 165608
rect 434222 165552 434227 165608
rect 433934 165550 434227 165552
rect 131573 165547 131639 165550
rect -960 165066 480 165156
rect 2773 165066 2839 165069
rect -960 165064 2839 165066
rect -960 165008 2778 165064
rect 2834 165008 2839 165064
rect 433934 165036 433994 165550
rect 434161 165547 434227 165550
rect -960 165006 2839 165008
rect -960 164916 480 165006
rect 2773 165003 2839 165006
rect 132677 164522 132743 164525
rect 132677 164520 134044 164522
rect 132677 164464 132682 164520
rect 132738 164464 134044 164520
rect 132677 164462 134044 164464
rect 132677 164459 132743 164462
rect 128353 164250 128419 164253
rect 128537 164250 128603 164253
rect 128353 164248 128603 164250
rect 128353 164192 128358 164248
rect 128414 164192 128542 164248
rect 128598 164192 128603 164248
rect 128353 164190 128603 164192
rect 128353 164187 128419 164190
rect 128537 164187 128603 164190
rect 132953 164250 133019 164253
rect 133137 164250 133203 164253
rect 132953 164248 133203 164250
rect 132953 164192 132958 164248
rect 133014 164192 133142 164248
rect 133198 164192 133203 164248
rect 132953 164190 133203 164192
rect 132953 164187 133019 164190
rect 133137 164187 133203 164190
rect 133505 163570 133571 163573
rect 434069 163570 434135 163573
rect 133505 163568 134044 163570
rect 133505 163512 133510 163568
rect 133566 163512 134044 163568
rect 133505 163510 134044 163512
rect 433934 163568 434135 163570
rect 433934 163512 434074 163568
rect 434130 163512 434135 163568
rect 433934 163510 434135 163512
rect 133505 163507 133571 163510
rect 433934 162996 433994 163510
rect 434069 163507 434135 163510
rect 132401 162482 132467 162485
rect 132401 162480 134044 162482
rect 132401 162424 132406 162480
rect 132462 162424 134044 162480
rect 132401 162422 134044 162424
rect 132401 162419 132467 162422
rect 133505 161394 133571 161397
rect 133505 161392 134044 161394
rect 133505 161336 133510 161392
rect 133566 161336 134044 161392
rect 133505 161334 134044 161336
rect 133505 161331 133571 161334
rect 436093 161258 436159 161261
rect 433934 161256 436159 161258
rect 433934 161200 436098 161256
rect 436154 161200 436159 161256
rect 433934 161198 436159 161200
rect 433934 160956 433994 161198
rect 436093 161195 436159 161198
rect 132033 160442 132099 160445
rect 132033 160440 134044 160442
rect 132033 160384 132038 160440
rect 132094 160384 134044 160440
rect 132033 160382 134044 160384
rect 132033 160379 132099 160382
rect 131205 159354 131271 159357
rect 433977 159354 434043 159357
rect 131205 159352 134044 159354
rect 131205 159296 131210 159352
rect 131266 159296 134044 159352
rect 131205 159294 134044 159296
rect 433934 159352 434043 159354
rect 433934 159296 433982 159352
rect 434038 159296 434043 159352
rect 131205 159291 131271 159294
rect 433934 159291 434043 159296
rect 433934 158780 433994 159291
rect 580625 158402 580691 158405
rect 583520 158402 584960 158492
rect 580625 158400 584960 158402
rect 580625 158344 580630 158400
rect 580686 158344 584960 158400
rect 580625 158342 584960 158344
rect 580625 158339 580691 158342
rect 131573 158266 131639 158269
rect 131573 158264 134044 158266
rect 131573 158208 131578 158264
rect 131634 158208 134044 158264
rect 583520 158252 584960 158342
rect 131573 158206 134044 158208
rect 131573 158203 131639 158206
rect 433885 157314 433951 157317
rect 433885 157312 433994 157314
rect 433885 157256 433890 157312
rect 433946 157256 433994 157312
rect 433885 157251 433994 157256
rect 130929 156634 130995 156637
rect 134014 156634 134074 157148
rect 433934 156740 433994 157251
rect 130929 156632 134074 156634
rect 130929 156576 130934 156632
rect 130990 156576 134074 156632
rect 130929 156574 134074 156576
rect 130929 156571 130995 156574
rect 131205 156226 131271 156229
rect 131205 156224 134044 156226
rect 131205 156168 131210 156224
rect 131266 156168 134044 156224
rect 131205 156166 134044 156168
rect 131205 156163 131271 156166
rect 131205 155138 131271 155141
rect 436093 155138 436159 155141
rect 131205 155136 134044 155138
rect 131205 155080 131210 155136
rect 131266 155080 134044 155136
rect 131205 155078 134044 155080
rect 433934 155136 436159 155138
rect 433934 155080 436098 155136
rect 436154 155080 436159 155136
rect 433934 155078 436159 155080
rect 131205 155075 131271 155078
rect 128537 154868 128603 154869
rect 128486 154866 128492 154868
rect 128446 154806 128492 154866
rect 128556 154864 128603 154868
rect 128598 154808 128603 154864
rect 128486 154804 128492 154806
rect 128556 154804 128603 154808
rect 128537 154803 128603 154804
rect 132953 154730 133019 154733
rect 132953 154728 133154 154730
rect 132953 154672 132958 154728
rect 133014 154672 133154 154728
rect 132953 154670 133154 154672
rect 132953 154667 133019 154670
rect 128537 154596 128603 154597
rect 128486 154532 128492 154596
rect 128556 154594 128603 154596
rect 132953 154594 133019 154597
rect 133094 154594 133154 154670
rect 128556 154592 128648 154594
rect 128598 154536 128648 154592
rect 128556 154534 128648 154536
rect 132953 154592 133154 154594
rect 132953 154536 132958 154592
rect 133014 154536 133154 154592
rect 433934 154564 433994 155078
rect 436093 155075 436159 155078
rect 504173 154594 504239 154597
rect 504449 154594 504515 154597
rect 504173 154592 504515 154594
rect 132953 154534 133154 154536
rect 504173 154536 504178 154592
rect 504234 154536 504454 154592
rect 504510 154536 504515 154592
rect 504173 154534 504515 154536
rect 128556 154532 128603 154534
rect 128537 154531 128603 154532
rect 132953 154531 133019 154534
rect 504173 154531 504239 154534
rect 504449 154531 504515 154534
rect 131205 154050 131271 154053
rect 131205 154048 134044 154050
rect 131205 153992 131210 154048
rect 131266 153992 134044 154048
rect 131205 153990 134044 153992
rect 131205 153987 131271 153990
rect 6913 153098 6979 153101
rect 16481 153098 16547 153101
rect 6913 153096 16547 153098
rect 6913 153040 6918 153096
rect 6974 153040 16486 153096
rect 16542 153040 16547 153096
rect 6913 153038 16547 153040
rect 6913 153035 6979 153038
rect 16481 153035 16547 153038
rect 131205 152962 131271 152965
rect 131205 152960 134044 152962
rect 131205 152904 131210 152960
rect 131266 152904 134044 152960
rect 131205 152902 134044 152904
rect 131205 152899 131271 152902
rect 433934 152282 433994 152524
rect 437381 152282 437447 152285
rect 433934 152280 437447 152282
rect 433934 152224 437386 152280
rect 437442 152224 437447 152280
rect 433934 152222 437447 152224
rect 437381 152219 437447 152222
rect 131205 152010 131271 152013
rect 131205 152008 134044 152010
rect 131205 151952 131210 152008
rect 131266 151952 134044 152008
rect 131205 151950 134044 151952
rect 131205 151947 131271 151950
rect 131205 150922 131271 150925
rect 131205 150920 134044 150922
rect -960 150786 480 150876
rect 131205 150864 131210 150920
rect 131266 150864 134044 150920
rect 131205 150862 134044 150864
rect 131205 150859 131271 150862
rect 4153 150786 4219 150789
rect -960 150784 4219 150786
rect -960 150728 4158 150784
rect 4214 150728 4219 150784
rect -960 150726 4219 150728
rect -960 150636 480 150726
rect 4153 150723 4219 150726
rect 433934 150242 433994 150348
rect 437013 150242 437079 150245
rect 433934 150240 437079 150242
rect 433934 150184 437018 150240
rect 437074 150184 437079 150240
rect 433934 150182 437079 150184
rect 437013 150179 437079 150182
rect 131205 149834 131271 149837
rect 131205 149832 134044 149834
rect 131205 149776 131210 149832
rect 131266 149776 134044 149832
rect 131205 149774 134044 149776
rect 131205 149771 131271 149774
rect 84193 148882 84259 148885
rect 93577 148882 93643 148885
rect 436185 148882 436251 148885
rect 84193 148880 93643 148882
rect 84193 148824 84198 148880
rect 84254 148824 93582 148880
rect 93638 148824 93643 148880
rect 84193 148822 93643 148824
rect 84193 148819 84259 148822
rect 93577 148819 93643 148822
rect 433934 148880 436251 148882
rect 433934 148824 436190 148880
rect 436246 148824 436251 148880
rect 433934 148822 436251 148824
rect 64873 148746 64939 148749
rect 70393 148746 70459 148749
rect 64873 148744 70459 148746
rect 64873 148688 64878 148744
rect 64934 148688 70398 148744
rect 70454 148688 70459 148744
rect 64873 148686 70459 148688
rect 64873 148683 64939 148686
rect 70393 148683 70459 148686
rect 131205 148746 131271 148749
rect 131205 148744 134044 148746
rect 131205 148688 131210 148744
rect 131266 148688 134044 148744
rect 131205 148686 134044 148688
rect 131205 148683 131271 148686
rect 131205 148338 131271 148341
rect 131205 148336 134074 148338
rect 131205 148280 131210 148336
rect 131266 148280 134074 148336
rect 433934 148308 433994 148822
rect 436185 148819 436251 148822
rect 131205 148278 134074 148280
rect 131205 148275 131271 148278
rect 132217 147796 132283 147797
rect 132166 147794 132172 147796
rect 132126 147734 132172 147794
rect 132236 147792 132283 147796
rect 132278 147736 132283 147792
rect 134014 147764 134074 148278
rect 132166 147732 132172 147734
rect 132236 147732 132283 147736
rect 132217 147731 132283 147732
rect 132166 147460 132172 147524
rect 132236 147522 132242 147524
rect 132309 147522 132375 147525
rect 132236 147520 132375 147522
rect 132236 147464 132314 147520
rect 132370 147464 132375 147520
rect 132236 147462 132375 147464
rect 132236 147460 132242 147462
rect 132309 147459 132375 147462
rect 132217 146706 132283 146709
rect 132217 146704 134044 146706
rect 132217 146648 132222 146704
rect 132278 146648 134044 146704
rect 132217 146646 134044 146648
rect 132217 146643 132283 146646
rect 583520 146556 584960 146796
rect 436093 146298 436159 146301
rect 433934 146296 436159 146298
rect 433934 146240 436098 146296
rect 436154 146240 436159 146296
rect 433934 146238 436159 146240
rect 433934 146132 433994 146238
rect 436093 146235 436159 146238
rect 131113 145618 131179 145621
rect 131113 145616 134044 145618
rect 131113 145560 131118 145616
rect 131174 145560 134044 145616
rect 131113 145558 134044 145560
rect 131113 145555 131179 145558
rect 131113 144530 131179 144533
rect 437381 144530 437447 144533
rect 131113 144528 134044 144530
rect 131113 144472 131118 144528
rect 131174 144472 134044 144528
rect 131113 144470 134044 144472
rect 433934 144528 437447 144530
rect 433934 144472 437386 144528
rect 437442 144472 437447 144528
rect 433934 144470 437447 144472
rect 131113 144467 131179 144470
rect 433934 144092 433994 144470
rect 437381 144467 437447 144470
rect 128997 143578 129063 143581
rect 128997 143576 134044 143578
rect 128997 143520 129002 143576
rect 129058 143520 134044 143576
rect 128997 143518 134044 143520
rect 128997 143515 129063 143518
rect 132309 142490 132375 142493
rect 132309 142488 134044 142490
rect 132309 142432 132314 142488
rect 132370 142432 134044 142488
rect 132309 142430 134044 142432
rect 132309 142427 132375 142430
rect 436093 142082 436159 142085
rect 433934 142080 436159 142082
rect 433934 142024 436098 142080
rect 436154 142024 436159 142080
rect 433934 142022 436159 142024
rect 433934 141916 433994 142022
rect 436093 142019 436159 142022
rect 133873 141402 133939 141405
rect 133873 141400 134044 141402
rect 133873 141344 133878 141400
rect 133934 141344 134044 141400
rect 133873 141342 134044 141344
rect 133873 141339 133939 141342
rect 132217 140450 132283 140453
rect 132217 140448 134044 140450
rect 132217 140392 132222 140448
rect 132278 140392 134044 140448
rect 132217 140390 134044 140392
rect 132217 140387 132283 140390
rect 437381 140314 437447 140317
rect 433934 140312 437447 140314
rect 433934 140256 437386 140312
rect 437442 140256 437447 140312
rect 433934 140254 437447 140256
rect 433934 139876 433994 140254
rect 437381 140251 437447 140254
rect 133597 139362 133663 139365
rect 133597 139360 134044 139362
rect 133597 139304 133602 139360
rect 133658 139304 134044 139360
rect 133597 139302 134044 139304
rect 133597 139299 133663 139302
rect 131113 138274 131179 138277
rect 131113 138272 134044 138274
rect 131113 138216 131118 138272
rect 131174 138216 134044 138272
rect 131113 138214 134044 138216
rect 131113 138211 131179 138214
rect 437381 137866 437447 137869
rect 433934 137864 437447 137866
rect 433934 137808 437386 137864
rect 437442 137808 437447 137864
rect 433934 137806 437447 137808
rect 433934 137700 433994 137806
rect 437381 137803 437447 137806
rect 133689 137186 133755 137189
rect 133689 137184 134044 137186
rect 133689 137128 133694 137184
rect 133750 137128 134044 137184
rect 133689 137126 134044 137128
rect 133689 137123 133755 137126
rect -960 136370 480 136460
rect 2773 136370 2839 136373
rect -960 136368 2839 136370
rect -960 136312 2778 136368
rect 2834 136312 2839 136368
rect -960 136310 2839 136312
rect -960 136220 480 136310
rect 2773 136307 2839 136310
rect 132493 136234 132559 136237
rect 132493 136232 134044 136234
rect 132493 136176 132498 136232
rect 132554 136176 134044 136232
rect 132493 136174 134044 136176
rect 132493 136171 132559 136174
rect 437013 136098 437079 136101
rect 433934 136096 437079 136098
rect 433934 136040 437018 136096
rect 437074 136040 437079 136096
rect 433934 136038 437079 136040
rect 433934 135660 433994 136038
rect 437013 136035 437079 136038
rect 132125 135146 132191 135149
rect 132125 135144 134044 135146
rect 132125 135088 132130 135144
rect 132186 135088 134044 135144
rect 132125 135086 134044 135088
rect 132125 135083 132191 135086
rect 580257 134874 580323 134877
rect 583520 134874 584960 134964
rect 580257 134872 584960 134874
rect 580257 134816 580262 134872
rect 580318 134816 584960 134872
rect 580257 134814 584960 134816
rect 580257 134811 580323 134814
rect 583520 134724 584960 134814
rect 131941 134058 132007 134061
rect 131941 134056 134044 134058
rect 131941 134000 131946 134056
rect 132002 134000 134044 134056
rect 131941 133998 134044 134000
rect 131941 133995 132007 133998
rect 437381 133650 437447 133653
rect 433934 133648 437447 133650
rect 433934 133592 437386 133648
rect 437442 133592 437447 133648
rect 433934 133590 437447 133592
rect 133965 133514 134031 133517
rect 133965 133512 134074 133514
rect 133965 133456 133970 133512
rect 134026 133456 134074 133512
rect 433934 133484 433994 133590
rect 437381 133587 437447 133590
rect 133965 133451 134074 133456
rect 134014 132940 134074 133451
rect 131297 132018 131363 132021
rect 436829 132018 436895 132021
rect 131297 132016 134044 132018
rect 131297 131960 131302 132016
rect 131358 131960 134044 132016
rect 131297 131958 134044 131960
rect 433934 132016 436895 132018
rect 433934 131960 436834 132016
rect 436890 131960 436895 132016
rect 433934 131958 436895 131960
rect 131297 131955 131363 131958
rect 433934 131444 433994 131958
rect 436829 131955 436895 131958
rect 131849 130930 131915 130933
rect 131849 130928 134044 130930
rect 131849 130872 131854 130928
rect 131910 130872 134044 130928
rect 131849 130870 134044 130872
rect 131849 130867 131915 130870
rect 134057 130386 134123 130389
rect 134014 130384 134123 130386
rect 134014 130328 134062 130384
rect 134118 130328 134123 130384
rect 134014 130323 134123 130328
rect 134014 129812 134074 130323
rect 437381 129570 437447 129573
rect 433934 129568 437447 129570
rect 433934 129512 437386 129568
rect 437442 129512 437447 129568
rect 433934 129510 437447 129512
rect 433934 129268 433994 129510
rect 437381 129507 437447 129510
rect 131389 128754 131455 128757
rect 131389 128752 134044 128754
rect 131389 128696 131394 128752
rect 131450 128696 134044 128752
rect 131389 128694 134044 128696
rect 131389 128691 131455 128694
rect 131481 127802 131547 127805
rect 436093 127802 436159 127805
rect 131481 127800 134044 127802
rect 131481 127744 131486 127800
rect 131542 127744 134044 127800
rect 131481 127742 134044 127744
rect 433934 127800 436159 127802
rect 433934 127744 436098 127800
rect 436154 127744 436159 127800
rect 433934 127742 436159 127744
rect 131481 127739 131547 127742
rect 433934 127228 433994 127742
rect 436093 127739 436159 127742
rect 131757 126714 131823 126717
rect 131757 126712 134044 126714
rect 131757 126656 131762 126712
rect 131818 126656 134044 126712
rect 131757 126654 134044 126656
rect 131757 126651 131823 126654
rect 128813 125626 128879 125629
rect 129089 125626 129155 125629
rect 128813 125624 129155 125626
rect 128813 125568 128818 125624
rect 128874 125568 129094 125624
rect 129150 125568 129155 125624
rect 128813 125566 129155 125568
rect 128813 125563 128879 125566
rect 129089 125563 129155 125566
rect 131665 125626 131731 125629
rect 131665 125624 134044 125626
rect 131665 125568 131670 125624
rect 131726 125568 134044 125624
rect 131665 125566 134044 125568
rect 131665 125563 131731 125566
rect 132769 124538 132835 124541
rect 433934 124538 433994 125052
rect 436921 124538 436987 124541
rect 132769 124536 134044 124538
rect 132769 124480 132774 124536
rect 132830 124480 134044 124536
rect 132769 124478 134044 124480
rect 433934 124536 436987 124538
rect 433934 124480 436926 124536
rect 436982 124480 436987 124536
rect 433934 124478 436987 124480
rect 132769 124475 132835 124478
rect 436921 124475 436987 124478
rect 134014 123045 134074 123556
rect 580901 123178 580967 123181
rect 583520 123178 584960 123268
rect 580901 123176 584960 123178
rect 580901 123120 580906 123176
rect 580962 123120 584960 123176
rect 580901 123118 584960 123120
rect 580901 123115 580967 123118
rect 133965 123040 134074 123045
rect 133965 122984 133970 123040
rect 134026 122984 134074 123040
rect 583520 123028 584960 123118
rect 133965 122982 134074 122984
rect 133965 122979 134031 122982
rect 433934 122906 433994 123012
rect 436829 122906 436895 122909
rect 433934 122904 436895 122906
rect 433934 122848 436834 122904
rect 436890 122848 436895 122904
rect 433934 122846 436895 122848
rect 436829 122843 436895 122846
rect -960 122090 480 122180
rect 3233 122090 3299 122093
rect -960 122088 3299 122090
rect -960 122032 3238 122088
rect 3294 122032 3299 122088
rect -960 122030 3299 122032
rect -960 121940 480 122030
rect 3233 122027 3299 122030
rect 134014 121957 134074 122468
rect 134014 121952 134123 121957
rect 134014 121896 134062 121952
rect 134118 121896 134123 121952
rect 134014 121894 134123 121896
rect 134057 121891 134123 121894
rect 132309 121410 132375 121413
rect 132309 121408 134044 121410
rect 132309 121352 132314 121408
rect 132370 121352 134044 121408
rect 132309 121350 134044 121352
rect 132309 121347 132375 121350
rect 132125 120458 132191 120461
rect 433934 120458 433994 120972
rect 436737 120458 436803 120461
rect 132125 120456 134044 120458
rect 132125 120400 132130 120456
rect 132186 120400 134044 120456
rect 132125 120398 134044 120400
rect 433934 120456 436803 120458
rect 433934 120400 436742 120456
rect 436798 120400 436803 120456
rect 433934 120398 436803 120400
rect 132125 120395 132191 120398
rect 436737 120395 436803 120398
rect 126973 118690 127039 118693
rect 151813 118690 151879 118693
rect 126973 118688 151879 118690
rect 126973 118632 126978 118688
rect 127034 118632 151818 118688
rect 151874 118632 151879 118688
rect 126973 118630 151879 118632
rect 126973 118627 127039 118630
rect 151813 118627 151879 118630
rect 132953 118554 133019 118557
rect 140773 118554 140839 118557
rect 132953 118552 140839 118554
rect 132953 118496 132958 118552
rect 133014 118496 140778 118552
rect 140834 118496 140839 118552
rect 132953 118494 140839 118496
rect 132953 118491 133019 118494
rect 140773 118491 140839 118494
rect 125777 118418 125843 118421
rect 197629 118418 197695 118421
rect 125777 118416 197695 118418
rect 125777 118360 125782 118416
rect 125838 118360 197634 118416
rect 197690 118360 197695 118416
rect 125777 118358 197695 118360
rect 125777 118355 125843 118358
rect 197629 118355 197695 118358
rect 126237 118282 126303 118285
rect 195973 118282 196039 118285
rect 126237 118280 196039 118282
rect 126237 118224 126242 118280
rect 126298 118224 195978 118280
rect 196034 118224 196039 118280
rect 126237 118222 196039 118224
rect 126237 118219 126303 118222
rect 195973 118219 196039 118222
rect 129181 118146 129247 118149
rect 133229 118146 133295 118149
rect 129181 118144 133295 118146
rect 129181 118088 129186 118144
rect 129242 118088 133234 118144
rect 133290 118088 133295 118144
rect 129181 118086 133295 118088
rect 129181 118083 129247 118086
rect 133229 118083 133295 118086
rect 133822 118084 133828 118148
rect 133892 118146 133898 118148
rect 182173 118146 182239 118149
rect 133892 118086 154498 118146
rect 133892 118084 133898 118086
rect 130377 118010 130443 118013
rect 146477 118010 146543 118013
rect 146845 118010 146911 118013
rect 130377 118008 146911 118010
rect 130377 117952 130382 118008
rect 130438 117952 146482 118008
rect 146538 117952 146850 118008
rect 146906 117952 146911 118008
rect 130377 117950 146911 117952
rect 154438 118010 154498 118086
rect 168974 118144 182239 118146
rect 168974 118088 182178 118144
rect 182234 118088 182239 118144
rect 168974 118086 182239 118088
rect 168974 118010 169034 118086
rect 182173 118083 182239 118086
rect 154438 117950 169034 118010
rect 130377 117947 130443 117950
rect 146477 117947 146543 117950
rect 146845 117947 146911 117950
rect 97993 117874 98059 117877
rect 99281 117874 99347 117877
rect 184933 117874 184999 117877
rect 97993 117872 184999 117874
rect 97993 117816 97998 117872
rect 98054 117816 99286 117872
rect 99342 117816 184938 117872
rect 184994 117816 184999 117872
rect 97993 117814 184999 117816
rect 97993 117811 98059 117814
rect 99281 117811 99347 117814
rect 184933 117811 184999 117814
rect 117221 117738 117287 117741
rect 193949 117738 194015 117741
rect 117221 117736 194015 117738
rect 117221 117680 117226 117736
rect 117282 117680 193954 117736
rect 194010 117680 194015 117736
rect 117221 117678 194015 117680
rect 117221 117675 117287 117678
rect 193949 117675 194015 117678
rect 133045 117602 133111 117605
rect 133822 117602 133828 117604
rect 133045 117600 133828 117602
rect 133045 117544 133050 117600
rect 133106 117544 133828 117600
rect 133045 117542 133828 117544
rect 133045 117539 133111 117542
rect 133822 117540 133828 117542
rect 133892 117540 133898 117604
rect 393221 117602 393287 117605
rect 383702 117600 393287 117602
rect 383702 117544 393226 117600
rect 393282 117544 393287 117600
rect 383702 117542 393287 117544
rect 383702 117469 383762 117542
rect 393221 117539 393287 117542
rect 383653 117464 383762 117469
rect 383653 117408 383658 117464
rect 383714 117408 383762 117464
rect 383653 117406 383762 117408
rect 383653 117403 383719 117406
rect 115933 117330 115999 117333
rect 117221 117330 117287 117333
rect 115933 117328 117287 117330
rect 115933 117272 115938 117328
rect 115994 117272 117226 117328
rect 117282 117272 117287 117328
rect 115933 117270 117287 117272
rect 115933 117267 115999 117270
rect 117221 117267 117287 117270
rect 171133 117194 171199 117197
rect 180701 117194 180767 117197
rect 171133 117192 180767 117194
rect 171133 117136 171138 117192
rect 171194 117136 180706 117192
rect 180762 117136 180767 117192
rect 171133 117134 180767 117136
rect 171133 117131 171199 117134
rect 180701 117131 180767 117134
rect 128813 115970 128879 115973
rect 128997 115970 129063 115973
rect 128813 115968 129063 115970
rect 128813 115912 128818 115968
rect 128874 115912 129002 115968
rect 129058 115912 129063 115968
rect 128813 115910 129063 115912
rect 128813 115907 128879 115910
rect 128997 115907 129063 115910
rect 152181 115970 152247 115973
rect 152457 115970 152523 115973
rect 152181 115968 152523 115970
rect 152181 115912 152186 115968
rect 152242 115912 152462 115968
rect 152518 115912 152523 115968
rect 152181 115910 152523 115912
rect 152181 115907 152247 115910
rect 152457 115907 152523 115910
rect 203057 115970 203123 115973
rect 203701 115970 203767 115973
rect 203057 115968 203767 115970
rect 203057 115912 203062 115968
rect 203118 115912 203706 115968
rect 203762 115912 203767 115968
rect 203057 115910 203767 115912
rect 203057 115907 203123 115910
rect 203701 115907 203767 115910
rect 204529 115970 204595 115973
rect 204897 115970 204963 115973
rect 204529 115968 204963 115970
rect 204529 115912 204534 115968
rect 204590 115912 204902 115968
rect 204958 115912 204963 115968
rect 204529 115910 204963 115912
rect 204529 115907 204595 115910
rect 204897 115907 204963 115910
rect 215937 115970 216003 115973
rect 216121 115970 216187 115973
rect 215937 115968 216187 115970
rect 215937 115912 215942 115968
rect 215998 115912 216126 115968
rect 216182 115912 216187 115968
rect 215937 115910 216187 115912
rect 215937 115907 216003 115910
rect 216121 115907 216187 115910
rect 217041 115970 217107 115973
rect 217409 115970 217475 115973
rect 217041 115968 217475 115970
rect 217041 115912 217046 115968
rect 217102 115912 217414 115968
rect 217470 115912 217475 115968
rect 217041 115910 217475 115912
rect 217041 115907 217107 115910
rect 217409 115907 217475 115910
rect 220169 115970 220235 115973
rect 220353 115970 220419 115973
rect 220169 115968 220419 115970
rect 220169 115912 220174 115968
rect 220230 115912 220358 115968
rect 220414 115912 220419 115968
rect 220169 115910 220419 115912
rect 220169 115907 220235 115910
rect 220353 115907 220419 115910
rect 221457 115970 221523 115973
rect 221641 115970 221707 115973
rect 221457 115968 221707 115970
rect 221457 115912 221462 115968
rect 221518 115912 221646 115968
rect 221702 115912 221707 115968
rect 221457 115910 221707 115912
rect 221457 115907 221523 115910
rect 221641 115907 221707 115910
rect 227989 115970 228055 115973
rect 228265 115970 228331 115973
rect 227989 115968 228331 115970
rect 227989 115912 227994 115968
rect 228050 115912 228270 115968
rect 228326 115912 228331 115968
rect 227989 115910 228331 115912
rect 227989 115907 228055 115910
rect 228265 115907 228331 115910
rect 338665 115970 338731 115973
rect 339033 115970 339099 115973
rect 338665 115968 339099 115970
rect 338665 115912 338670 115968
rect 338726 115912 339038 115968
rect 339094 115912 339099 115968
rect 338665 115910 339099 115912
rect 338665 115907 338731 115910
rect 339033 115907 339099 115910
rect 431309 114746 431375 114749
rect 431309 114744 431786 114746
rect 431309 114688 431314 114744
rect 431370 114688 431786 114744
rect 431309 114686 431786 114688
rect 431309 114683 431375 114686
rect 431585 114610 431651 114613
rect 431726 114610 431786 114686
rect 431585 114608 431786 114610
rect 431585 114552 431590 114608
rect 431646 114552 431786 114608
rect 431585 114550 431786 114552
rect 431585 114547 431651 114550
rect 579797 111482 579863 111485
rect 583520 111482 584960 111572
rect 579797 111480 584960 111482
rect 579797 111424 579802 111480
rect 579858 111424 584960 111480
rect 579797 111422 584960 111424
rect 579797 111419 579863 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3233 107674 3299 107677
rect -960 107672 3299 107674
rect -960 107616 3238 107672
rect 3294 107616 3299 107672
rect -960 107614 3299 107616
rect -960 107524 480 107614
rect 3233 107611 3299 107614
rect 140865 106450 140931 106453
rect 140822 106448 140931 106450
rect 140822 106392 140870 106448
rect 140926 106392 140931 106448
rect 140822 106387 140931 106392
rect 246941 106450 247007 106453
rect 246941 106448 247050 106450
rect 246941 106392 246946 106448
rect 247002 106392 247050 106448
rect 246941 106387 247050 106392
rect 140822 106317 140882 106387
rect 246990 106317 247050 106387
rect 128721 106314 128787 106317
rect 128905 106314 128971 106317
rect 128721 106312 128971 106314
rect 128721 106256 128726 106312
rect 128782 106256 128910 106312
rect 128966 106256 128971 106312
rect 128721 106254 128971 106256
rect 128721 106251 128787 106254
rect 128905 106251 128971 106254
rect 140773 106312 140882 106317
rect 140773 106256 140778 106312
rect 140834 106256 140882 106312
rect 140773 106254 140882 106256
rect 145097 106314 145163 106317
rect 145281 106314 145347 106317
rect 145097 106312 145347 106314
rect 145097 106256 145102 106312
rect 145158 106256 145286 106312
rect 145342 106256 145347 106312
rect 145097 106254 145347 106256
rect 140773 106251 140839 106254
rect 145097 106251 145163 106254
rect 145281 106251 145347 106254
rect 238937 106314 239003 106317
rect 239121 106314 239187 106317
rect 238937 106312 239187 106314
rect 238937 106256 238942 106312
rect 238998 106256 239126 106312
rect 239182 106256 239187 106312
rect 238937 106254 239187 106256
rect 238937 106251 239003 106254
rect 239121 106251 239187 106254
rect 246941 106312 247050 106317
rect 246941 106256 246946 106312
rect 247002 106256 247050 106312
rect 246941 106254 247050 106256
rect 383101 106314 383167 106317
rect 383285 106314 383351 106317
rect 383101 106312 383351 106314
rect 383101 106256 383106 106312
rect 383162 106256 383290 106312
rect 383346 106256 383351 106312
rect 383101 106254 383351 106256
rect 246941 106251 247007 106254
rect 383101 106251 383167 106254
rect 383285 106251 383351 106254
rect 148041 104954 148107 104957
rect 148225 104954 148291 104957
rect 148041 104952 148291 104954
rect 148041 104896 148046 104952
rect 148102 104896 148230 104952
rect 148286 104896 148291 104952
rect 148041 104894 148291 104896
rect 148041 104891 148107 104894
rect 148225 104891 148291 104894
rect 218237 104818 218303 104821
rect 218102 104816 218303 104818
rect 218102 104760 218242 104816
rect 218298 104760 218303 104816
rect 218102 104758 218303 104760
rect 218102 104682 218162 104758
rect 218237 104755 218303 104758
rect 218421 104682 218487 104685
rect 218102 104680 218487 104682
rect 218102 104624 218426 104680
rect 218482 104624 218487 104680
rect 218102 104622 218487 104624
rect 218421 104619 218487 104622
rect 583520 99636 584960 99876
rect 274909 96794 274975 96797
rect 274774 96792 274975 96794
rect 274774 96736 274914 96792
rect 274970 96736 274975 96792
rect 274774 96734 274975 96736
rect 274774 96661 274834 96734
rect 274909 96731 274975 96734
rect 274725 96656 274834 96661
rect 274725 96600 274730 96656
rect 274786 96600 274834 96656
rect 274725 96598 274834 96600
rect 274725 96595 274791 96598
rect -960 93258 480 93348
rect 3417 93258 3483 93261
rect -960 93256 3483 93258
rect -960 93200 3422 93256
rect 3478 93200 3483 93256
rect -960 93198 3483 93200
rect -960 93108 480 93198
rect 3417 93195 3483 93198
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect 204621 87002 204687 87005
rect 204805 87002 204871 87005
rect 204621 87000 204871 87002
rect 204621 86944 204626 87000
rect 204682 86944 204810 87000
rect 204866 86944 204871 87000
rect 204621 86942 204871 86944
rect 204621 86939 204687 86942
rect 204805 86939 204871 86942
rect 209957 87002 210023 87005
rect 210141 87002 210207 87005
rect 209957 87000 210207 87002
rect 209957 86944 209962 87000
rect 210018 86944 210146 87000
rect 210202 86944 210207 87000
rect 209957 86942 210207 86944
rect 209957 86939 210023 86942
rect 210141 86939 210207 86942
rect 274449 87002 274515 87005
rect 274633 87002 274699 87005
rect 274449 87000 274699 87002
rect 274449 86944 274454 87000
rect 274510 86944 274638 87000
rect 274694 86944 274699 87000
rect 274449 86942 274699 86944
rect 274449 86939 274515 86942
rect 274633 86939 274699 86942
rect 425973 87002 426039 87005
rect 426157 87002 426223 87005
rect 425973 87000 426223 87002
rect 425973 86944 425978 87000
rect 426034 86944 426162 87000
rect 426218 86944 426223 87000
rect 425973 86942 426223 86944
rect 425973 86939 426039 86942
rect 426157 86939 426223 86942
rect 276105 85642 276171 85645
rect 276289 85642 276355 85645
rect 276105 85640 276355 85642
rect 276105 85584 276110 85640
rect 276166 85584 276294 85640
rect 276350 85584 276355 85640
rect 276105 85582 276355 85584
rect 276105 85579 276171 85582
rect 276289 85579 276355 85582
rect 233417 80202 233483 80205
rect 233374 80200 233483 80202
rect 233374 80144 233422 80200
rect 233478 80144 233483 80200
rect 233374 80139 233483 80144
rect 233233 79930 233299 79933
rect 233374 79930 233434 80139
rect 233233 79928 233434 79930
rect 233233 79872 233238 79928
rect 233294 79872 233434 79928
rect 233233 79870 233434 79872
rect 233233 79867 233299 79870
rect -960 78978 480 79068
rect 3141 78978 3207 78981
rect -960 78976 3207 78978
rect -960 78920 3146 78976
rect 3202 78920 3207 78976
rect -960 78918 3207 78920
rect -960 78828 480 78918
rect 3141 78915 3207 78918
rect 383193 77210 383259 77213
rect 383653 77210 383719 77213
rect 383193 77208 383719 77210
rect 383193 77152 383198 77208
rect 383254 77152 383658 77208
rect 383714 77152 383719 77208
rect 383193 77150 383719 77152
rect 383193 77147 383259 77150
rect 383653 77147 383719 77150
rect 420729 77210 420795 77213
rect 421005 77210 421071 77213
rect 420729 77208 421071 77210
rect 420729 77152 420734 77208
rect 420790 77152 421010 77208
rect 421066 77152 421071 77208
rect 420729 77150 421071 77152
rect 420729 77147 420795 77150
rect 421005 77147 421071 77150
rect 580165 76258 580231 76261
rect 583520 76258 584960 76348
rect 580165 76256 584960 76258
rect 580165 76200 580170 76256
rect 580226 76200 584960 76256
rect 580165 76198 584960 76200
rect 580165 76195 580231 76198
rect 583520 76108 584960 76198
rect 144821 75850 144887 75853
rect 145005 75850 145071 75853
rect 144821 75848 145071 75850
rect 144821 75792 144826 75848
rect 144882 75792 145010 75848
rect 145066 75792 145071 75848
rect 144821 75790 145071 75792
rect 144821 75787 144887 75790
rect 145005 75787 145071 75790
rect 244273 75850 244339 75853
rect 244641 75850 244707 75853
rect 244273 75848 244707 75850
rect 244273 75792 244278 75848
rect 244334 75792 244646 75848
rect 244702 75792 244707 75848
rect 244273 75790 244707 75792
rect 244273 75787 244339 75790
rect 244641 75787 244707 75790
rect 128905 67826 128971 67829
rect 128905 67824 129290 67826
rect 128905 67768 128910 67824
rect 128966 67768 129290 67824
rect 128905 67766 129290 67768
rect 128905 67763 128971 67766
rect 129089 67690 129155 67693
rect 129230 67690 129290 67766
rect 129089 67688 129290 67690
rect 129089 67632 129094 67688
rect 129150 67632 129290 67688
rect 129089 67630 129290 67632
rect 129089 67627 129155 67630
rect 221089 66330 221155 66333
rect 221273 66330 221339 66333
rect 221089 66328 221339 66330
rect 221089 66272 221094 66328
rect 221150 66272 221278 66328
rect 221334 66272 221339 66328
rect 221089 66270 221339 66272
rect 221089 66267 221155 66270
rect 221273 66267 221339 66270
rect 431585 66330 431651 66333
rect 431769 66330 431835 66333
rect 431585 66328 431835 66330
rect 431585 66272 431590 66328
rect 431646 66272 431774 66328
rect 431830 66272 431835 66328
rect 431585 66270 431835 66272
rect 431585 66267 431651 66270
rect 431769 66267 431835 66270
rect 145097 66194 145163 66197
rect 145097 66192 145298 66194
rect 145097 66136 145102 66192
rect 145158 66136 145298 66192
rect 145097 66134 145298 66136
rect 145097 66131 145163 66134
rect 145238 66061 145298 66134
rect 145189 66056 145298 66061
rect 145189 66000 145194 66056
rect 145250 66000 145298 66056
rect 145189 65998 145298 66000
rect 145189 65995 145255 65998
rect 426065 64970 426131 64973
rect 426433 64970 426499 64973
rect 426065 64968 426499 64970
rect 426065 64912 426070 64968
rect 426126 64912 426438 64968
rect 426494 64912 426499 64968
rect 426065 64910 426499 64912
rect 426065 64907 426131 64910
rect 426433 64907 426499 64910
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 140773 60892 140839 60893
rect 140773 60888 140820 60892
rect 140884 60890 140890 60892
rect 140773 60832 140778 60888
rect 140773 60828 140820 60832
rect 140884 60830 140930 60890
rect 140884 60828 140890 60830
rect 140773 60827 140839 60828
rect 140773 55316 140839 55317
rect 140773 55312 140820 55316
rect 140884 55314 140890 55316
rect 140773 55256 140778 55312
rect 140773 55252 140820 55256
rect 140884 55254 140930 55314
rect 140884 55252 140890 55254
rect 140773 55251 140839 55252
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 4061 50146 4127 50149
rect -960 50144 4127 50146
rect -960 50088 4066 50144
rect 4122 50088 4127 50144
rect -960 50086 4127 50088
rect -960 49996 480 50086
rect 4061 50083 4127 50086
rect 420453 48378 420519 48381
rect 420637 48378 420703 48381
rect 420453 48376 420703 48378
rect 420453 48320 420458 48376
rect 420514 48320 420642 48376
rect 420698 48320 420703 48376
rect 420453 48318 420703 48320
rect 420453 48315 420519 48318
rect 420637 48315 420703 48318
rect 143717 44162 143783 44165
rect 143993 44162 144059 44165
rect 143717 44160 144059 44162
rect 143717 44104 143722 44160
rect 143778 44104 143998 44160
rect 144054 44104 144059 44160
rect 143717 44102 144059 44104
rect 143717 44099 143783 44102
rect 143993 44099 144059 44102
rect 425789 44162 425855 44165
rect 425973 44162 426039 44165
rect 425789 44160 426039 44162
rect 425789 44104 425794 44160
rect 425850 44104 425978 44160
rect 426034 44104 426039 44160
rect 425789 44102 426039 44104
rect 425789 44099 425855 44102
rect 425973 44099 426039 44102
rect 140865 41442 140931 41445
rect 140822 41440 140931 41442
rect 140822 41384 140870 41440
rect 140926 41384 140931 41440
rect 140822 41379 140931 41384
rect 140822 41309 140882 41379
rect 140773 41304 140882 41309
rect 140773 41248 140778 41304
rect 140834 41248 140882 41304
rect 140773 41246 140882 41248
rect 140773 41243 140839 41246
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect 183369 37226 183435 37229
rect 183645 37226 183711 37229
rect 183369 37224 183711 37226
rect 183369 37168 183374 37224
rect 183430 37168 183650 37224
rect 183706 37168 183711 37224
rect 183369 37166 183711 37168
rect 183369 37163 183435 37166
rect 183645 37163 183711 37166
rect -960 35866 480 35956
rect 3417 35866 3483 35869
rect -960 35864 3483 35866
rect -960 35808 3422 35864
rect 3478 35808 3483 35864
rect -960 35806 3483 35808
rect -960 35716 480 35806
rect 3417 35803 3483 35806
rect 580165 29338 580231 29341
rect 583520 29338 584960 29428
rect 580165 29336 584960 29338
rect 580165 29280 580170 29336
rect 580226 29280 584960 29336
rect 580165 29278 584960 29280
rect 580165 29275 580231 29278
rect 164601 29202 164667 29205
rect 164374 29200 164667 29202
rect 164374 29144 164606 29200
rect 164662 29144 164667 29200
rect 583520 29188 584960 29278
rect 164374 29142 164667 29144
rect 164374 29066 164434 29142
rect 164601 29139 164667 29142
rect 164509 29066 164575 29069
rect 164374 29064 164575 29066
rect 164374 29008 164514 29064
rect 164570 29008 164575 29064
rect 164374 29006 164575 29008
rect 164509 29003 164575 29006
rect 189073 29066 189139 29069
rect 420453 29066 420519 29069
rect 189073 29064 189274 29066
rect 189073 29008 189078 29064
rect 189134 29008 189274 29064
rect 189073 29006 189274 29008
rect 189073 29003 189139 29006
rect 189214 28930 189274 29006
rect 420453 29064 420562 29066
rect 420453 29008 420458 29064
rect 420514 29032 420562 29064
rect 420637 29032 420703 29035
rect 420514 29030 420703 29032
rect 420514 29008 420642 29030
rect 420453 29003 420642 29008
rect 420502 28974 420642 29003
rect 420698 28974 420703 29030
rect 420502 28972 420703 28974
rect 420637 28969 420703 28972
rect 189349 28930 189415 28933
rect 189214 28928 189415 28930
rect 189214 28872 189354 28928
rect 189410 28872 189415 28928
rect 189214 28870 189415 28872
rect 189349 28867 189415 28870
rect 227805 28930 227871 28933
rect 227989 28930 228055 28933
rect 227805 28928 228055 28930
rect 227805 28872 227810 28928
rect 227866 28872 227994 28928
rect 228050 28872 228055 28928
rect 227805 28870 228055 28872
rect 227805 28867 227871 28870
rect 227989 28867 228055 28870
rect 383285 28932 383351 28933
rect 383285 28928 383332 28932
rect 383396 28930 383402 28932
rect 383285 28872 383290 28928
rect 383285 28868 383332 28872
rect 383396 28870 383442 28930
rect 383396 28868 383402 28870
rect 383285 28867 383351 28868
rect 383377 21996 383443 21997
rect 383326 21994 383332 21996
rect 383286 21934 383332 21994
rect 383396 21992 383443 21996
rect 383438 21936 383443 21992
rect 383326 21932 383332 21934
rect 383396 21932 383443 21936
rect 383377 21931 383443 21932
rect -960 21450 480 21540
rect 2773 21450 2839 21453
rect -960 21448 2839 21450
rect -960 21392 2778 21448
rect 2834 21392 2839 21448
rect -960 21390 2839 21392
rect -960 21300 480 21390
rect 2773 21387 2839 21390
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect 183921 9890 183987 9893
rect 246941 9890 247007 9893
rect 183510 9888 183987 9890
rect 183510 9832 183926 9888
rect 183982 9832 183987 9888
rect 183510 9830 183987 9832
rect 183510 9754 183570 9830
rect 183921 9827 183987 9830
rect 246622 9888 247007 9890
rect 246622 9832 246946 9888
rect 247002 9832 247007 9888
rect 246622 9830 247007 9832
rect 183645 9754 183711 9757
rect 183510 9752 183711 9754
rect 183510 9696 183650 9752
rect 183706 9696 183711 9752
rect 183510 9694 183711 9696
rect 246622 9754 246682 9830
rect 246941 9827 247007 9830
rect 246757 9754 246823 9757
rect 246622 9752 246823 9754
rect 246622 9696 246762 9752
rect 246818 9696 246823 9752
rect 246622 9694 246823 9696
rect 183645 9691 183711 9694
rect 246757 9691 246823 9694
rect 174261 9618 174327 9621
rect 181069 9618 181135 9621
rect 174261 9616 181135 9618
rect 174261 9560 174266 9616
rect 174322 9560 181074 9616
rect 181130 9560 181135 9616
rect 174261 9558 181135 9560
rect 174261 9555 174327 9558
rect 181069 9555 181135 9558
rect -960 7170 480 7260
rect 3877 7170 3943 7173
rect -960 7168 3943 7170
rect -960 7112 3882 7168
rect 3938 7112 3943 7168
rect -960 7110 3943 7112
rect -960 7020 480 7110
rect 3877 7107 3943 7110
rect 376753 6898 376819 6901
rect 379605 6898 379671 6901
rect 376753 6896 379671 6898
rect 376753 6840 376758 6896
rect 376814 6840 379610 6896
rect 379666 6840 379671 6896
rect 376753 6838 379671 6840
rect 376753 6835 376819 6838
rect 379605 6835 379671 6838
rect 583520 5796 584960 6036
<< via3 >>
rect 271644 502344 271708 502348
rect 271644 502288 271658 502344
rect 271658 502288 271708 502344
rect 271644 502284 271708 502288
rect 271644 492628 271708 492692
rect 281212 260808 281276 260812
rect 281212 260752 281226 260808
rect 281226 260752 281276 260808
rect 281212 260748 281276 260752
rect 281212 251228 281276 251292
rect 133092 200092 133156 200156
rect 132908 196072 132972 196076
rect 132908 196016 132922 196072
rect 132922 196016 132972 196072
rect 132908 196012 132972 196016
rect 132908 195936 132972 195940
rect 132908 195880 132922 195936
rect 132922 195880 132972 195936
rect 132908 195876 132972 195880
rect 132908 185404 132972 185468
rect 133092 184920 133156 184924
rect 133092 184864 133106 184920
rect 133106 184864 133156 184920
rect 133092 184860 133156 184864
rect 132908 182336 132972 182340
rect 132908 182280 132922 182336
rect 132922 182280 132972 182336
rect 132908 182276 132972 182280
rect 128492 154864 128556 154868
rect 128492 154808 128542 154864
rect 128542 154808 128556 154864
rect 128492 154804 128556 154808
rect 128492 154592 128556 154596
rect 128492 154536 128542 154592
rect 128542 154536 128556 154592
rect 128492 154532 128556 154536
rect 132172 147792 132236 147796
rect 132172 147736 132222 147792
rect 132222 147736 132236 147792
rect 132172 147732 132236 147736
rect 132172 147460 132236 147524
rect 133828 118084 133892 118148
rect 133828 117540 133892 117604
rect 140820 60888 140884 60892
rect 140820 60832 140834 60888
rect 140834 60832 140884 60888
rect 140820 60828 140884 60832
rect 140820 55312 140884 55316
rect 140820 55256 140834 55312
rect 140834 55256 140884 55312
rect 140820 55252 140884 55256
rect 383332 28928 383396 28932
rect 383332 28872 383346 28928
rect 383346 28872 383396 28928
rect 383332 28868 383396 28872
rect 383332 21992 383396 21996
rect 383332 21936 383382 21992
rect 383382 21936 383396 21992
rect 383332 21932 383396 21936
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 679254 -7976 710862
rect -8576 679018 -8394 679254
rect -8158 679018 -7976 679254
rect -8576 678934 -7976 679018
rect -8576 678698 -8394 678934
rect -8158 678698 -7976 678934
rect -8576 643254 -7976 678698
rect -8576 643018 -8394 643254
rect -8158 643018 -7976 643254
rect -8576 642934 -7976 643018
rect -8576 642698 -8394 642934
rect -8158 642698 -7976 642934
rect -8576 607254 -7976 642698
rect -8576 607018 -8394 607254
rect -8158 607018 -7976 607254
rect -8576 606934 -7976 607018
rect -8576 606698 -8394 606934
rect -8158 606698 -7976 606934
rect -8576 571254 -7976 606698
rect -8576 571018 -8394 571254
rect -8158 571018 -7976 571254
rect -8576 570934 -7976 571018
rect -8576 570698 -8394 570934
rect -8158 570698 -7976 570934
rect -8576 535254 -7976 570698
rect -8576 535018 -8394 535254
rect -8158 535018 -7976 535254
rect -8576 534934 -7976 535018
rect -8576 534698 -8394 534934
rect -8158 534698 -7976 534934
rect -8576 499254 -7976 534698
rect -8576 499018 -8394 499254
rect -8158 499018 -7976 499254
rect -8576 498934 -7976 499018
rect -8576 498698 -8394 498934
rect -8158 498698 -7976 498934
rect -8576 463254 -7976 498698
rect -8576 463018 -8394 463254
rect -8158 463018 -7976 463254
rect -8576 462934 -7976 463018
rect -8576 462698 -8394 462934
rect -8158 462698 -7976 462934
rect -8576 427254 -7976 462698
rect -8576 427018 -8394 427254
rect -8158 427018 -7976 427254
rect -8576 426934 -7976 427018
rect -8576 426698 -8394 426934
rect -8158 426698 -7976 426934
rect -8576 391254 -7976 426698
rect -8576 391018 -8394 391254
rect -8158 391018 -7976 391254
rect -8576 390934 -7976 391018
rect -8576 390698 -8394 390934
rect -8158 390698 -7976 390934
rect -8576 355254 -7976 390698
rect -8576 355018 -8394 355254
rect -8158 355018 -7976 355254
rect -8576 354934 -7976 355018
rect -8576 354698 -8394 354934
rect -8158 354698 -7976 354934
rect -8576 319254 -7976 354698
rect -8576 319018 -8394 319254
rect -8158 319018 -7976 319254
rect -8576 318934 -7976 319018
rect -8576 318698 -8394 318934
rect -8158 318698 -7976 318934
rect -8576 283254 -7976 318698
rect -8576 283018 -8394 283254
rect -8158 283018 -7976 283254
rect -8576 282934 -7976 283018
rect -8576 282698 -8394 282934
rect -8158 282698 -7976 282934
rect -8576 247254 -7976 282698
rect -8576 247018 -8394 247254
rect -8158 247018 -7976 247254
rect -8576 246934 -7976 247018
rect -8576 246698 -8394 246934
rect -8158 246698 -7976 246934
rect -8576 211254 -7976 246698
rect -8576 211018 -8394 211254
rect -8158 211018 -7976 211254
rect -8576 210934 -7976 211018
rect -8576 210698 -8394 210934
rect -8158 210698 -7976 210934
rect -8576 175254 -7976 210698
rect -8576 175018 -8394 175254
rect -8158 175018 -7976 175254
rect -8576 174934 -7976 175018
rect -8576 174698 -8394 174934
rect -8158 174698 -7976 174934
rect -8576 139254 -7976 174698
rect -8576 139018 -8394 139254
rect -8158 139018 -7976 139254
rect -8576 138934 -7976 139018
rect -8576 138698 -8394 138934
rect -8158 138698 -7976 138934
rect -8576 103254 -7976 138698
rect -8576 103018 -8394 103254
rect -8158 103018 -7976 103254
rect -8576 102934 -7976 103018
rect -8576 102698 -8394 102934
rect -8158 102698 -7976 102934
rect -8576 67254 -7976 102698
rect -8576 67018 -8394 67254
rect -8158 67018 -7976 67254
rect -8576 66934 -7976 67018
rect -8576 66698 -8394 66934
rect -8158 66698 -7976 66934
rect -8576 31254 -7976 66698
rect -8576 31018 -8394 31254
rect -8158 31018 -7976 31254
rect -8576 30934 -7976 31018
rect -8576 30698 -8394 30934
rect -8158 30698 -7976 30934
rect -8576 -6926 -7976 30698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 697254 -7036 709922
rect 11604 710478 12204 711440
rect 11604 710242 11786 710478
rect 12022 710242 12204 710478
rect 11604 710158 12204 710242
rect 11604 709922 11786 710158
rect 12022 709922 12204 710158
rect -7636 697018 -7454 697254
rect -7218 697018 -7036 697254
rect -7636 696934 -7036 697018
rect -7636 696698 -7454 696934
rect -7218 696698 -7036 696934
rect -7636 661254 -7036 696698
rect -7636 661018 -7454 661254
rect -7218 661018 -7036 661254
rect -7636 660934 -7036 661018
rect -7636 660698 -7454 660934
rect -7218 660698 -7036 660934
rect -7636 625254 -7036 660698
rect -7636 625018 -7454 625254
rect -7218 625018 -7036 625254
rect -7636 624934 -7036 625018
rect -7636 624698 -7454 624934
rect -7218 624698 -7036 624934
rect -7636 589254 -7036 624698
rect -7636 589018 -7454 589254
rect -7218 589018 -7036 589254
rect -7636 588934 -7036 589018
rect -7636 588698 -7454 588934
rect -7218 588698 -7036 588934
rect -7636 553254 -7036 588698
rect -7636 553018 -7454 553254
rect -7218 553018 -7036 553254
rect -7636 552934 -7036 553018
rect -7636 552698 -7454 552934
rect -7218 552698 -7036 552934
rect -7636 517254 -7036 552698
rect -7636 517018 -7454 517254
rect -7218 517018 -7036 517254
rect -7636 516934 -7036 517018
rect -7636 516698 -7454 516934
rect -7218 516698 -7036 516934
rect -7636 481254 -7036 516698
rect -7636 481018 -7454 481254
rect -7218 481018 -7036 481254
rect -7636 480934 -7036 481018
rect -7636 480698 -7454 480934
rect -7218 480698 -7036 480934
rect -7636 445254 -7036 480698
rect -7636 445018 -7454 445254
rect -7218 445018 -7036 445254
rect -7636 444934 -7036 445018
rect -7636 444698 -7454 444934
rect -7218 444698 -7036 444934
rect -7636 409254 -7036 444698
rect -7636 409018 -7454 409254
rect -7218 409018 -7036 409254
rect -7636 408934 -7036 409018
rect -7636 408698 -7454 408934
rect -7218 408698 -7036 408934
rect -7636 373254 -7036 408698
rect -7636 373018 -7454 373254
rect -7218 373018 -7036 373254
rect -7636 372934 -7036 373018
rect -7636 372698 -7454 372934
rect -7218 372698 -7036 372934
rect -7636 337254 -7036 372698
rect -7636 337018 -7454 337254
rect -7218 337018 -7036 337254
rect -7636 336934 -7036 337018
rect -7636 336698 -7454 336934
rect -7218 336698 -7036 336934
rect -7636 301254 -7036 336698
rect -7636 301018 -7454 301254
rect -7218 301018 -7036 301254
rect -7636 300934 -7036 301018
rect -7636 300698 -7454 300934
rect -7218 300698 -7036 300934
rect -7636 265254 -7036 300698
rect -7636 265018 -7454 265254
rect -7218 265018 -7036 265254
rect -7636 264934 -7036 265018
rect -7636 264698 -7454 264934
rect -7218 264698 -7036 264934
rect -7636 229254 -7036 264698
rect -7636 229018 -7454 229254
rect -7218 229018 -7036 229254
rect -7636 228934 -7036 229018
rect -7636 228698 -7454 228934
rect -7218 228698 -7036 228934
rect -7636 193254 -7036 228698
rect -7636 193018 -7454 193254
rect -7218 193018 -7036 193254
rect -7636 192934 -7036 193018
rect -7636 192698 -7454 192934
rect -7218 192698 -7036 192934
rect -7636 157254 -7036 192698
rect -7636 157018 -7454 157254
rect -7218 157018 -7036 157254
rect -7636 156934 -7036 157018
rect -7636 156698 -7454 156934
rect -7218 156698 -7036 156934
rect -7636 121254 -7036 156698
rect -7636 121018 -7454 121254
rect -7218 121018 -7036 121254
rect -7636 120934 -7036 121018
rect -7636 120698 -7454 120934
rect -7218 120698 -7036 120934
rect -7636 85254 -7036 120698
rect -7636 85018 -7454 85254
rect -7218 85018 -7036 85254
rect -7636 84934 -7036 85018
rect -7636 84698 -7454 84934
rect -7218 84698 -7036 84934
rect -7636 49254 -7036 84698
rect -7636 49018 -7454 49254
rect -7218 49018 -7036 49254
rect -7636 48934 -7036 49018
rect -7636 48698 -7454 48934
rect -7218 48698 -7036 48934
rect -7636 13254 -7036 48698
rect -7636 13018 -7454 13254
rect -7218 13018 -7036 13254
rect -7636 12934 -7036 13018
rect -7636 12698 -7454 12934
rect -7218 12698 -7036 12934
rect -7636 -5986 -7036 12698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 675654 -6096 708982
rect -6696 675418 -6514 675654
rect -6278 675418 -6096 675654
rect -6696 675334 -6096 675418
rect -6696 675098 -6514 675334
rect -6278 675098 -6096 675334
rect -6696 639654 -6096 675098
rect -6696 639418 -6514 639654
rect -6278 639418 -6096 639654
rect -6696 639334 -6096 639418
rect -6696 639098 -6514 639334
rect -6278 639098 -6096 639334
rect -6696 603654 -6096 639098
rect -6696 603418 -6514 603654
rect -6278 603418 -6096 603654
rect -6696 603334 -6096 603418
rect -6696 603098 -6514 603334
rect -6278 603098 -6096 603334
rect -6696 567654 -6096 603098
rect -6696 567418 -6514 567654
rect -6278 567418 -6096 567654
rect -6696 567334 -6096 567418
rect -6696 567098 -6514 567334
rect -6278 567098 -6096 567334
rect -6696 531654 -6096 567098
rect -6696 531418 -6514 531654
rect -6278 531418 -6096 531654
rect -6696 531334 -6096 531418
rect -6696 531098 -6514 531334
rect -6278 531098 -6096 531334
rect -6696 495654 -6096 531098
rect -6696 495418 -6514 495654
rect -6278 495418 -6096 495654
rect -6696 495334 -6096 495418
rect -6696 495098 -6514 495334
rect -6278 495098 -6096 495334
rect -6696 459654 -6096 495098
rect -6696 459418 -6514 459654
rect -6278 459418 -6096 459654
rect -6696 459334 -6096 459418
rect -6696 459098 -6514 459334
rect -6278 459098 -6096 459334
rect -6696 423654 -6096 459098
rect -6696 423418 -6514 423654
rect -6278 423418 -6096 423654
rect -6696 423334 -6096 423418
rect -6696 423098 -6514 423334
rect -6278 423098 -6096 423334
rect -6696 387654 -6096 423098
rect -6696 387418 -6514 387654
rect -6278 387418 -6096 387654
rect -6696 387334 -6096 387418
rect -6696 387098 -6514 387334
rect -6278 387098 -6096 387334
rect -6696 351654 -6096 387098
rect -6696 351418 -6514 351654
rect -6278 351418 -6096 351654
rect -6696 351334 -6096 351418
rect -6696 351098 -6514 351334
rect -6278 351098 -6096 351334
rect -6696 315654 -6096 351098
rect -6696 315418 -6514 315654
rect -6278 315418 -6096 315654
rect -6696 315334 -6096 315418
rect -6696 315098 -6514 315334
rect -6278 315098 -6096 315334
rect -6696 279654 -6096 315098
rect -6696 279418 -6514 279654
rect -6278 279418 -6096 279654
rect -6696 279334 -6096 279418
rect -6696 279098 -6514 279334
rect -6278 279098 -6096 279334
rect -6696 243654 -6096 279098
rect -6696 243418 -6514 243654
rect -6278 243418 -6096 243654
rect -6696 243334 -6096 243418
rect -6696 243098 -6514 243334
rect -6278 243098 -6096 243334
rect -6696 207654 -6096 243098
rect -6696 207418 -6514 207654
rect -6278 207418 -6096 207654
rect -6696 207334 -6096 207418
rect -6696 207098 -6514 207334
rect -6278 207098 -6096 207334
rect -6696 171654 -6096 207098
rect -6696 171418 -6514 171654
rect -6278 171418 -6096 171654
rect -6696 171334 -6096 171418
rect -6696 171098 -6514 171334
rect -6278 171098 -6096 171334
rect -6696 135654 -6096 171098
rect -6696 135418 -6514 135654
rect -6278 135418 -6096 135654
rect -6696 135334 -6096 135418
rect -6696 135098 -6514 135334
rect -6278 135098 -6096 135334
rect -6696 99654 -6096 135098
rect -6696 99418 -6514 99654
rect -6278 99418 -6096 99654
rect -6696 99334 -6096 99418
rect -6696 99098 -6514 99334
rect -6278 99098 -6096 99334
rect -6696 63654 -6096 99098
rect -6696 63418 -6514 63654
rect -6278 63418 -6096 63654
rect -6696 63334 -6096 63418
rect -6696 63098 -6514 63334
rect -6278 63098 -6096 63334
rect -6696 27654 -6096 63098
rect -6696 27418 -6514 27654
rect -6278 27418 -6096 27654
rect -6696 27334 -6096 27418
rect -6696 27098 -6514 27334
rect -6278 27098 -6096 27334
rect -6696 -5046 -6096 27098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 693654 -5156 708042
rect 8004 708598 8604 709560
rect 8004 708362 8186 708598
rect 8422 708362 8604 708598
rect 8004 708278 8604 708362
rect 8004 708042 8186 708278
rect 8422 708042 8604 708278
rect -5756 693418 -5574 693654
rect -5338 693418 -5156 693654
rect -5756 693334 -5156 693418
rect -5756 693098 -5574 693334
rect -5338 693098 -5156 693334
rect -5756 657654 -5156 693098
rect -5756 657418 -5574 657654
rect -5338 657418 -5156 657654
rect -5756 657334 -5156 657418
rect -5756 657098 -5574 657334
rect -5338 657098 -5156 657334
rect -5756 621654 -5156 657098
rect -5756 621418 -5574 621654
rect -5338 621418 -5156 621654
rect -5756 621334 -5156 621418
rect -5756 621098 -5574 621334
rect -5338 621098 -5156 621334
rect -5756 585654 -5156 621098
rect -5756 585418 -5574 585654
rect -5338 585418 -5156 585654
rect -5756 585334 -5156 585418
rect -5756 585098 -5574 585334
rect -5338 585098 -5156 585334
rect -5756 549654 -5156 585098
rect -5756 549418 -5574 549654
rect -5338 549418 -5156 549654
rect -5756 549334 -5156 549418
rect -5756 549098 -5574 549334
rect -5338 549098 -5156 549334
rect -5756 513654 -5156 549098
rect -5756 513418 -5574 513654
rect -5338 513418 -5156 513654
rect -5756 513334 -5156 513418
rect -5756 513098 -5574 513334
rect -5338 513098 -5156 513334
rect -5756 477654 -5156 513098
rect -5756 477418 -5574 477654
rect -5338 477418 -5156 477654
rect -5756 477334 -5156 477418
rect -5756 477098 -5574 477334
rect -5338 477098 -5156 477334
rect -5756 441654 -5156 477098
rect -5756 441418 -5574 441654
rect -5338 441418 -5156 441654
rect -5756 441334 -5156 441418
rect -5756 441098 -5574 441334
rect -5338 441098 -5156 441334
rect -5756 405654 -5156 441098
rect -5756 405418 -5574 405654
rect -5338 405418 -5156 405654
rect -5756 405334 -5156 405418
rect -5756 405098 -5574 405334
rect -5338 405098 -5156 405334
rect -5756 369654 -5156 405098
rect -5756 369418 -5574 369654
rect -5338 369418 -5156 369654
rect -5756 369334 -5156 369418
rect -5756 369098 -5574 369334
rect -5338 369098 -5156 369334
rect -5756 333654 -5156 369098
rect -5756 333418 -5574 333654
rect -5338 333418 -5156 333654
rect -5756 333334 -5156 333418
rect -5756 333098 -5574 333334
rect -5338 333098 -5156 333334
rect -5756 297654 -5156 333098
rect -5756 297418 -5574 297654
rect -5338 297418 -5156 297654
rect -5756 297334 -5156 297418
rect -5756 297098 -5574 297334
rect -5338 297098 -5156 297334
rect -5756 261654 -5156 297098
rect -5756 261418 -5574 261654
rect -5338 261418 -5156 261654
rect -5756 261334 -5156 261418
rect -5756 261098 -5574 261334
rect -5338 261098 -5156 261334
rect -5756 225654 -5156 261098
rect -5756 225418 -5574 225654
rect -5338 225418 -5156 225654
rect -5756 225334 -5156 225418
rect -5756 225098 -5574 225334
rect -5338 225098 -5156 225334
rect -5756 189654 -5156 225098
rect -5756 189418 -5574 189654
rect -5338 189418 -5156 189654
rect -5756 189334 -5156 189418
rect -5756 189098 -5574 189334
rect -5338 189098 -5156 189334
rect -5756 153654 -5156 189098
rect -5756 153418 -5574 153654
rect -5338 153418 -5156 153654
rect -5756 153334 -5156 153418
rect -5756 153098 -5574 153334
rect -5338 153098 -5156 153334
rect -5756 117654 -5156 153098
rect -5756 117418 -5574 117654
rect -5338 117418 -5156 117654
rect -5756 117334 -5156 117418
rect -5756 117098 -5574 117334
rect -5338 117098 -5156 117334
rect -5756 81654 -5156 117098
rect -5756 81418 -5574 81654
rect -5338 81418 -5156 81654
rect -5756 81334 -5156 81418
rect -5756 81098 -5574 81334
rect -5338 81098 -5156 81334
rect -5756 45654 -5156 81098
rect -5756 45418 -5574 45654
rect -5338 45418 -5156 45654
rect -5756 45334 -5156 45418
rect -5756 45098 -5574 45334
rect -5338 45098 -5156 45334
rect -5756 9654 -5156 45098
rect -5756 9418 -5574 9654
rect -5338 9418 -5156 9654
rect -5756 9334 -5156 9418
rect -5756 9098 -5574 9334
rect -5338 9098 -5156 9334
rect -5756 -4106 -5156 9098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 672054 -4216 707102
rect -4816 671818 -4634 672054
rect -4398 671818 -4216 672054
rect -4816 671734 -4216 671818
rect -4816 671498 -4634 671734
rect -4398 671498 -4216 671734
rect -4816 636054 -4216 671498
rect -4816 635818 -4634 636054
rect -4398 635818 -4216 636054
rect -4816 635734 -4216 635818
rect -4816 635498 -4634 635734
rect -4398 635498 -4216 635734
rect -4816 600054 -4216 635498
rect -4816 599818 -4634 600054
rect -4398 599818 -4216 600054
rect -4816 599734 -4216 599818
rect -4816 599498 -4634 599734
rect -4398 599498 -4216 599734
rect -4816 564054 -4216 599498
rect -4816 563818 -4634 564054
rect -4398 563818 -4216 564054
rect -4816 563734 -4216 563818
rect -4816 563498 -4634 563734
rect -4398 563498 -4216 563734
rect -4816 528054 -4216 563498
rect -4816 527818 -4634 528054
rect -4398 527818 -4216 528054
rect -4816 527734 -4216 527818
rect -4816 527498 -4634 527734
rect -4398 527498 -4216 527734
rect -4816 492054 -4216 527498
rect -4816 491818 -4634 492054
rect -4398 491818 -4216 492054
rect -4816 491734 -4216 491818
rect -4816 491498 -4634 491734
rect -4398 491498 -4216 491734
rect -4816 456054 -4216 491498
rect -4816 455818 -4634 456054
rect -4398 455818 -4216 456054
rect -4816 455734 -4216 455818
rect -4816 455498 -4634 455734
rect -4398 455498 -4216 455734
rect -4816 420054 -4216 455498
rect -4816 419818 -4634 420054
rect -4398 419818 -4216 420054
rect -4816 419734 -4216 419818
rect -4816 419498 -4634 419734
rect -4398 419498 -4216 419734
rect -4816 384054 -4216 419498
rect -4816 383818 -4634 384054
rect -4398 383818 -4216 384054
rect -4816 383734 -4216 383818
rect -4816 383498 -4634 383734
rect -4398 383498 -4216 383734
rect -4816 348054 -4216 383498
rect -4816 347818 -4634 348054
rect -4398 347818 -4216 348054
rect -4816 347734 -4216 347818
rect -4816 347498 -4634 347734
rect -4398 347498 -4216 347734
rect -4816 312054 -4216 347498
rect -4816 311818 -4634 312054
rect -4398 311818 -4216 312054
rect -4816 311734 -4216 311818
rect -4816 311498 -4634 311734
rect -4398 311498 -4216 311734
rect -4816 276054 -4216 311498
rect -4816 275818 -4634 276054
rect -4398 275818 -4216 276054
rect -4816 275734 -4216 275818
rect -4816 275498 -4634 275734
rect -4398 275498 -4216 275734
rect -4816 240054 -4216 275498
rect -4816 239818 -4634 240054
rect -4398 239818 -4216 240054
rect -4816 239734 -4216 239818
rect -4816 239498 -4634 239734
rect -4398 239498 -4216 239734
rect -4816 204054 -4216 239498
rect -4816 203818 -4634 204054
rect -4398 203818 -4216 204054
rect -4816 203734 -4216 203818
rect -4816 203498 -4634 203734
rect -4398 203498 -4216 203734
rect -4816 168054 -4216 203498
rect -4816 167818 -4634 168054
rect -4398 167818 -4216 168054
rect -4816 167734 -4216 167818
rect -4816 167498 -4634 167734
rect -4398 167498 -4216 167734
rect -4816 132054 -4216 167498
rect -4816 131818 -4634 132054
rect -4398 131818 -4216 132054
rect -4816 131734 -4216 131818
rect -4816 131498 -4634 131734
rect -4398 131498 -4216 131734
rect -4816 96054 -4216 131498
rect -4816 95818 -4634 96054
rect -4398 95818 -4216 96054
rect -4816 95734 -4216 95818
rect -4816 95498 -4634 95734
rect -4398 95498 -4216 95734
rect -4816 60054 -4216 95498
rect -4816 59818 -4634 60054
rect -4398 59818 -4216 60054
rect -4816 59734 -4216 59818
rect -4816 59498 -4634 59734
rect -4398 59498 -4216 59734
rect -4816 24054 -4216 59498
rect -4816 23818 -4634 24054
rect -4398 23818 -4216 24054
rect -4816 23734 -4216 23818
rect -4816 23498 -4634 23734
rect -4398 23498 -4216 23734
rect -4816 -3166 -4216 23498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 690054 -3276 706162
rect 4404 706718 5004 707680
rect 4404 706482 4586 706718
rect 4822 706482 5004 706718
rect 4404 706398 5004 706482
rect 4404 706162 4586 706398
rect 4822 706162 5004 706398
rect -3876 689818 -3694 690054
rect -3458 689818 -3276 690054
rect -3876 689734 -3276 689818
rect -3876 689498 -3694 689734
rect -3458 689498 -3276 689734
rect -3876 654054 -3276 689498
rect -3876 653818 -3694 654054
rect -3458 653818 -3276 654054
rect -3876 653734 -3276 653818
rect -3876 653498 -3694 653734
rect -3458 653498 -3276 653734
rect -3876 618054 -3276 653498
rect -3876 617818 -3694 618054
rect -3458 617818 -3276 618054
rect -3876 617734 -3276 617818
rect -3876 617498 -3694 617734
rect -3458 617498 -3276 617734
rect -3876 582054 -3276 617498
rect -3876 581818 -3694 582054
rect -3458 581818 -3276 582054
rect -3876 581734 -3276 581818
rect -3876 581498 -3694 581734
rect -3458 581498 -3276 581734
rect -3876 546054 -3276 581498
rect -3876 545818 -3694 546054
rect -3458 545818 -3276 546054
rect -3876 545734 -3276 545818
rect -3876 545498 -3694 545734
rect -3458 545498 -3276 545734
rect -3876 510054 -3276 545498
rect -3876 509818 -3694 510054
rect -3458 509818 -3276 510054
rect -3876 509734 -3276 509818
rect -3876 509498 -3694 509734
rect -3458 509498 -3276 509734
rect -3876 474054 -3276 509498
rect -3876 473818 -3694 474054
rect -3458 473818 -3276 474054
rect -3876 473734 -3276 473818
rect -3876 473498 -3694 473734
rect -3458 473498 -3276 473734
rect -3876 438054 -3276 473498
rect -3876 437818 -3694 438054
rect -3458 437818 -3276 438054
rect -3876 437734 -3276 437818
rect -3876 437498 -3694 437734
rect -3458 437498 -3276 437734
rect -3876 402054 -3276 437498
rect -3876 401818 -3694 402054
rect -3458 401818 -3276 402054
rect -3876 401734 -3276 401818
rect -3876 401498 -3694 401734
rect -3458 401498 -3276 401734
rect -3876 366054 -3276 401498
rect -3876 365818 -3694 366054
rect -3458 365818 -3276 366054
rect -3876 365734 -3276 365818
rect -3876 365498 -3694 365734
rect -3458 365498 -3276 365734
rect -3876 330054 -3276 365498
rect -3876 329818 -3694 330054
rect -3458 329818 -3276 330054
rect -3876 329734 -3276 329818
rect -3876 329498 -3694 329734
rect -3458 329498 -3276 329734
rect -3876 294054 -3276 329498
rect -3876 293818 -3694 294054
rect -3458 293818 -3276 294054
rect -3876 293734 -3276 293818
rect -3876 293498 -3694 293734
rect -3458 293498 -3276 293734
rect -3876 258054 -3276 293498
rect -3876 257818 -3694 258054
rect -3458 257818 -3276 258054
rect -3876 257734 -3276 257818
rect -3876 257498 -3694 257734
rect -3458 257498 -3276 257734
rect -3876 222054 -3276 257498
rect -3876 221818 -3694 222054
rect -3458 221818 -3276 222054
rect -3876 221734 -3276 221818
rect -3876 221498 -3694 221734
rect -3458 221498 -3276 221734
rect -3876 186054 -3276 221498
rect -3876 185818 -3694 186054
rect -3458 185818 -3276 186054
rect -3876 185734 -3276 185818
rect -3876 185498 -3694 185734
rect -3458 185498 -3276 185734
rect -3876 150054 -3276 185498
rect -3876 149818 -3694 150054
rect -3458 149818 -3276 150054
rect -3876 149734 -3276 149818
rect -3876 149498 -3694 149734
rect -3458 149498 -3276 149734
rect -3876 114054 -3276 149498
rect -3876 113818 -3694 114054
rect -3458 113818 -3276 114054
rect -3876 113734 -3276 113818
rect -3876 113498 -3694 113734
rect -3458 113498 -3276 113734
rect -3876 78054 -3276 113498
rect -3876 77818 -3694 78054
rect -3458 77818 -3276 78054
rect -3876 77734 -3276 77818
rect -3876 77498 -3694 77734
rect -3458 77498 -3276 77734
rect -3876 42054 -3276 77498
rect -3876 41818 -3694 42054
rect -3458 41818 -3276 42054
rect -3876 41734 -3276 41818
rect -3876 41498 -3694 41734
rect -3458 41498 -3276 41734
rect -3876 6054 -3276 41498
rect -3876 5818 -3694 6054
rect -3458 5818 -3276 6054
rect -3876 5734 -3276 5818
rect -3876 5498 -3694 5734
rect -3458 5498 -3276 5734
rect -3876 -2226 -3276 5498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 4404 690054 5004 706162
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 4404 -2226 5004 5498
rect 4404 -2462 4586 -2226
rect 4822 -2462 5004 -2226
rect 4404 -2546 5004 -2462
rect 4404 -2782 4586 -2546
rect 4822 -2782 5004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 4404 -3744 5004 -2782
rect 8004 693654 8604 708042
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 8004 -4106 8604 9098
rect 8004 -4342 8186 -4106
rect 8422 -4342 8604 -4106
rect 8004 -4426 8604 -4342
rect 8004 -4662 8186 -4426
rect 8422 -4662 8604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 8004 -5624 8604 -4662
rect 11604 697254 12204 709922
rect 29604 711418 30204 711440
rect 29604 711182 29786 711418
rect 30022 711182 30204 711418
rect 29604 711098 30204 711182
rect 29604 710862 29786 711098
rect 30022 710862 30204 711098
rect 26004 709538 26604 709560
rect 26004 709302 26186 709538
rect 26422 709302 26604 709538
rect 26004 709218 26604 709302
rect 26004 708982 26186 709218
rect 26422 708982 26604 709218
rect 22404 707658 23004 707680
rect 22404 707422 22586 707658
rect 22822 707422 23004 707658
rect 22404 707338 23004 707422
rect 22404 707102 22586 707338
rect 22822 707102 23004 707338
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 11604 -5986 12204 12698
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 22404 672054 23004 707102
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3166 23004 23498
rect 22404 -3402 22586 -3166
rect 22822 -3402 23004 -3166
rect 22404 -3486 23004 -3402
rect 22404 -3722 22586 -3486
rect 22822 -3722 23004 -3486
rect 22404 -3744 23004 -3722
rect 26004 675654 26604 708982
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -5046 26604 27098
rect 26004 -5282 26186 -5046
rect 26422 -5282 26604 -5046
rect 26004 -5366 26604 -5282
rect 26004 -5602 26186 -5366
rect 26422 -5602 26604 -5366
rect 26004 -5624 26604 -5602
rect 29604 679254 30204 710862
rect 47604 710478 48204 711440
rect 47604 710242 47786 710478
rect 48022 710242 48204 710478
rect 47604 710158 48204 710242
rect 47604 709922 47786 710158
rect 48022 709922 48204 710158
rect 44004 708598 44604 709560
rect 44004 708362 44186 708598
rect 44422 708362 44604 708598
rect 44004 708278 44604 708362
rect 44004 708042 44186 708278
rect 44422 708042 44604 708278
rect 40404 706718 41004 707680
rect 40404 706482 40586 706718
rect 40822 706482 41004 706718
rect 40404 706398 41004 706482
rect 40404 706162 40586 706398
rect 40822 706162 41004 706398
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6222 11786 -5986
rect 12022 -6222 12204 -5986
rect 11604 -6306 12204 -6222
rect 11604 -6542 11786 -6306
rect 12022 -6542 12204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 11604 -7504 12204 -6542
rect 29604 -6926 30204 30698
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 40404 690054 41004 706162
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2226 41004 5498
rect 40404 -2462 40586 -2226
rect 40822 -2462 41004 -2226
rect 40404 -2546 41004 -2462
rect 40404 -2782 40586 -2546
rect 40822 -2782 41004 -2546
rect 40404 -3744 41004 -2782
rect 44004 693654 44604 708042
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4106 44604 9098
rect 44004 -4342 44186 -4106
rect 44422 -4342 44604 -4106
rect 44004 -4426 44604 -4342
rect 44004 -4662 44186 -4426
rect 44422 -4662 44604 -4426
rect 44004 -5624 44604 -4662
rect 47604 697254 48204 709922
rect 65604 711418 66204 711440
rect 65604 711182 65786 711418
rect 66022 711182 66204 711418
rect 65604 711098 66204 711182
rect 65604 710862 65786 711098
rect 66022 710862 66204 711098
rect 62004 709538 62604 709560
rect 62004 709302 62186 709538
rect 62422 709302 62604 709538
rect 62004 709218 62604 709302
rect 62004 708982 62186 709218
rect 62422 708982 62604 709218
rect 58404 707658 59004 707680
rect 58404 707422 58586 707658
rect 58822 707422 59004 707658
rect 58404 707338 59004 707422
rect 58404 707102 58586 707338
rect 58822 707102 59004 707338
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7162 29786 -6926
rect 30022 -7162 30204 -6926
rect 29604 -7246 30204 -7162
rect 29604 -7482 29786 -7246
rect 30022 -7482 30204 -7246
rect 29604 -7504 30204 -7482
rect 47604 -5986 48204 12698
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 58404 672054 59004 707102
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3166 59004 23498
rect 58404 -3402 58586 -3166
rect 58822 -3402 59004 -3166
rect 58404 -3486 59004 -3402
rect 58404 -3722 58586 -3486
rect 58822 -3722 59004 -3486
rect 58404 -3744 59004 -3722
rect 62004 675654 62604 708982
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -5046 62604 27098
rect 62004 -5282 62186 -5046
rect 62422 -5282 62604 -5046
rect 62004 -5366 62604 -5282
rect 62004 -5602 62186 -5366
rect 62422 -5602 62604 -5366
rect 62004 -5624 62604 -5602
rect 65604 679254 66204 710862
rect 83604 710478 84204 711440
rect 83604 710242 83786 710478
rect 84022 710242 84204 710478
rect 83604 710158 84204 710242
rect 83604 709922 83786 710158
rect 84022 709922 84204 710158
rect 80004 708598 80604 709560
rect 80004 708362 80186 708598
rect 80422 708362 80604 708598
rect 80004 708278 80604 708362
rect 80004 708042 80186 708278
rect 80422 708042 80604 708278
rect 76404 706718 77004 707680
rect 76404 706482 76586 706718
rect 76822 706482 77004 706718
rect 76404 706398 77004 706482
rect 76404 706162 76586 706398
rect 76822 706162 77004 706398
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 396550 73404 397898
rect 76404 690054 77004 706162
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 396550 77004 401498
rect 80004 693654 80604 708042
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 396550 80604 405098
rect 83604 697254 84204 709922
rect 101604 711418 102204 711440
rect 101604 711182 101786 711418
rect 102022 711182 102204 711418
rect 101604 711098 102204 711182
rect 101604 710862 101786 711098
rect 102022 710862 102204 711098
rect 98004 709538 98604 709560
rect 98004 709302 98186 709538
rect 98422 709302 98604 709538
rect 98004 709218 98604 709302
rect 98004 708982 98186 709218
rect 98422 708982 98604 709218
rect 94404 707658 95004 707680
rect 94404 707422 94586 707658
rect 94822 707422 95004 707658
rect 94404 707338 95004 707422
rect 94404 707102 94586 707338
rect 94822 707102 95004 707338
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 552104 91404 559898
rect 94404 672054 95004 707102
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 552104 95004 563498
rect 98004 675654 98604 708982
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 552104 98604 567098
rect 101604 679254 102204 710862
rect 119604 710478 120204 711440
rect 119604 710242 119786 710478
rect 120022 710242 120204 710478
rect 119604 710158 120204 710242
rect 119604 709922 119786 710158
rect 120022 709922 120204 710158
rect 116004 708598 116604 709560
rect 116004 708362 116186 708598
rect 116422 708362 116604 708598
rect 116004 708278 116604 708362
rect 116004 708042 116186 708278
rect 116422 708042 116604 708278
rect 112404 706718 113004 707680
rect 112404 706482 112586 706718
rect 112822 706482 113004 706718
rect 112404 706398 113004 706482
rect 112404 706162 112586 706398
rect 112822 706162 113004 706398
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 552104 102204 570698
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 552104 109404 577898
rect 112404 690054 113004 706162
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 552104 113004 581498
rect 116004 693654 116604 708042
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 91529 542454 91849 542476
rect 91529 542218 91571 542454
rect 91807 542218 91849 542454
rect 91529 542134 91849 542218
rect 91529 541898 91571 542134
rect 91807 541898 91849 542134
rect 91529 541876 91849 541898
rect 96113 524454 96433 524476
rect 96113 524218 96155 524454
rect 96391 524218 96433 524454
rect 96113 524134 96433 524218
rect 96113 523898 96155 524134
rect 96391 523898 96433 524134
rect 96113 523876 96433 523898
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 396550 84204 408698
rect 90804 488454 91404 519800
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 396550 91404 415898
rect 94404 492054 95004 519800
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 396550 95004 419498
rect 98004 495654 98604 519800
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 396550 98604 423098
rect 101604 499254 102204 519800
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 396550 102204 426698
rect 108804 506454 109404 519800
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 396550 109404 397898
rect 112404 510054 113004 519800
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 396550 113004 401498
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 396550 116604 405098
rect 119604 697254 120204 709922
rect 137604 711418 138204 711440
rect 137604 711182 137786 711418
rect 138022 711182 138204 711418
rect 137604 711098 138204 711182
rect 137604 710862 137786 711098
rect 138022 710862 138204 711098
rect 134004 709538 134604 709560
rect 134004 709302 134186 709538
rect 134422 709302 134604 709538
rect 134004 709218 134604 709302
rect 134004 708982 134186 709218
rect 134422 708982 134604 709218
rect 130404 707658 131004 707680
rect 130404 707422 130586 707658
rect 130822 707422 131004 707658
rect 130404 707338 131004 707422
rect 130404 707102 130586 707338
rect 130822 707102 131004 707338
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 553254 120204 588698
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 396550 120204 408698
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 91568 380454 91888 380476
rect 91568 380218 91610 380454
rect 91846 380218 91888 380454
rect 91568 380134 91888 380218
rect 91568 379898 91610 380134
rect 91846 379898 91888 380134
rect 91568 379876 91888 379898
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 76208 362454 76528 362476
rect 76208 362218 76250 362454
rect 76486 362218 76528 362454
rect 76208 362134 76528 362218
rect 76208 361898 76250 362134
rect 76486 361898 76528 362134
rect 76208 361876 76528 361898
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 91568 344454 91888 344476
rect 91568 344218 91610 344454
rect 91846 344218 91888 344454
rect 91568 344134 91888 344218
rect 91568 343898 91610 344134
rect 91846 343898 91888 344134
rect 91568 343876 91888 343898
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6222 47786 -5986
rect 48022 -6222 48204 -5986
rect 47604 -6306 48204 -6222
rect 47604 -6542 47786 -6306
rect 48022 -6542 48204 -6306
rect 47604 -7504 48204 -6542
rect 65604 -6926 66204 30698
rect 72804 326454 73404 339800
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 76404 330054 77004 339800
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2226 77004 5498
rect 76404 -2462 76586 -2226
rect 76822 -2462 77004 -2226
rect 76404 -2546 77004 -2462
rect 76404 -2782 76586 -2546
rect 76822 -2782 77004 -2546
rect 76404 -3744 77004 -2782
rect 80004 333654 80604 339800
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4106 80604 9098
rect 80004 -4342 80186 -4106
rect 80422 -4342 80604 -4106
rect 80004 -4426 80604 -4342
rect 80004 -4662 80186 -4426
rect 80422 -4662 80604 -4426
rect 80004 -5624 80604 -4662
rect 83604 337254 84204 339800
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7162 65786 -6926
rect 66022 -7162 66204 -6926
rect 65604 -7246 66204 -7162
rect 65604 -7482 65786 -7246
rect 66022 -7482 66204 -7246
rect 65604 -7504 66204 -7482
rect 83604 -5986 84204 12698
rect 90804 308454 91404 339800
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 94404 312054 95004 339800
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3166 95004 23498
rect 94404 -3402 94586 -3166
rect 94822 -3402 95004 -3166
rect 94404 -3486 95004 -3402
rect 94404 -3722 94586 -3486
rect 94822 -3722 95004 -3486
rect 94404 -3744 95004 -3722
rect 98004 315654 98604 339800
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -5046 98604 27098
rect 98004 -5282 98186 -5046
rect 98422 -5282 98604 -5046
rect 98004 -5366 98604 -5282
rect 98004 -5602 98186 -5366
rect 98422 -5602 98604 -5366
rect 98004 -5624 98604 -5602
rect 101604 319254 102204 339800
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6222 83786 -5986
rect 84022 -6222 84204 -5986
rect 83604 -6306 84204 -6222
rect 83604 -6542 83786 -6306
rect 84022 -6542 84204 -6306
rect 83604 -7504 84204 -6542
rect 101604 -6926 102204 30698
rect 108804 326454 109404 339800
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 112404 330054 113004 339800
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2226 113004 5498
rect 112404 -2462 112586 -2226
rect 112822 -2462 113004 -2226
rect 112404 -2546 113004 -2462
rect 112404 -2782 112586 -2546
rect 112822 -2782 113004 -2546
rect 112404 -3744 113004 -2782
rect 116004 333654 116604 339800
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4106 116604 9098
rect 116004 -4342 116186 -4106
rect 116422 -4342 116604 -4106
rect 116004 -4426 116604 -4342
rect 116004 -4662 116186 -4426
rect 116422 -4662 116604 -4426
rect 116004 -5624 116604 -4662
rect 119604 337254 120204 339800
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7162 101786 -6926
rect 102022 -7162 102204 -6926
rect 101604 -7246 102204 -7162
rect 101604 -7482 101786 -7246
rect 102022 -7482 102204 -7246
rect 101604 -7504 102204 -7482
rect 119604 -5986 120204 12698
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 130404 672054 131004 707102
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 134004 675654 134604 708982
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 200200 134604 207098
rect 137604 679254 138204 710862
rect 155604 710478 156204 711440
rect 155604 710242 155786 710478
rect 156022 710242 156204 710478
rect 155604 710158 156204 710242
rect 155604 709922 155786 710158
rect 156022 709922 156204 710158
rect 152004 708598 152604 709560
rect 152004 708362 152186 708598
rect 152422 708362 152604 708598
rect 152004 708278 152604 708362
rect 152004 708042 152186 708278
rect 152422 708042 152604 708278
rect 148404 706718 149004 707680
rect 148404 706482 148586 706718
rect 148822 706482 149004 706718
rect 148404 706398 149004 706482
rect 148404 706162 148586 706398
rect 148822 706162 149004 706398
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 535254 138204 570698
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 200200 138204 210698
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 200200 145404 217898
rect 148404 690054 149004 706162
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 200200 149004 221498
rect 152004 693654 152604 708042
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 200200 152604 225098
rect 155604 697254 156204 709922
rect 173604 711418 174204 711440
rect 173604 711182 173786 711418
rect 174022 711182 174204 711418
rect 173604 711098 174204 711182
rect 173604 710862 173786 711098
rect 174022 710862 174204 711098
rect 170004 709538 170604 709560
rect 170004 709302 170186 709538
rect 170422 709302 170604 709538
rect 170004 709218 170604 709302
rect 170004 708982 170186 709218
rect 170422 708982 170604 709218
rect 166404 707658 167004 707680
rect 166404 707422 166586 707658
rect 166822 707422 167004 707658
rect 166404 707338 167004 707422
rect 166404 707102 166586 707338
rect 166822 707102 167004 707338
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 409254 156204 444698
rect 155604 409018 155786 409254
rect 156022 409018 156204 409254
rect 155604 408934 156204 409018
rect 155604 408698 155786 408934
rect 156022 408698 156204 408934
rect 155604 373254 156204 408698
rect 155604 373018 155786 373254
rect 156022 373018 156204 373254
rect 155604 372934 156204 373018
rect 155604 372698 155786 372934
rect 156022 372698 156204 372934
rect 155604 337254 156204 372698
rect 155604 337018 155786 337254
rect 156022 337018 156204 337254
rect 155604 336934 156204 337018
rect 155604 336698 155786 336934
rect 156022 336698 156204 336934
rect 155604 301254 156204 336698
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 200200 156204 228698
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200200 163404 235898
rect 166404 672054 167004 707102
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 384054 167004 419498
rect 166404 383818 166586 384054
rect 166822 383818 167004 384054
rect 166404 383734 167004 383818
rect 166404 383498 166586 383734
rect 166822 383498 167004 383734
rect 166404 348054 167004 383498
rect 166404 347818 166586 348054
rect 166822 347818 167004 348054
rect 166404 347734 167004 347818
rect 166404 347498 166586 347734
rect 166822 347498 167004 347734
rect 166404 312054 167004 347498
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 200200 167004 203498
rect 170004 675654 170604 708982
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 387654 170604 423098
rect 170004 387418 170186 387654
rect 170422 387418 170604 387654
rect 170004 387334 170604 387418
rect 170004 387098 170186 387334
rect 170422 387098 170604 387334
rect 170004 351654 170604 387098
rect 170004 351418 170186 351654
rect 170422 351418 170604 351654
rect 170004 351334 170604 351418
rect 170004 351098 170186 351334
rect 170422 351098 170604 351334
rect 170004 315654 170604 351098
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 200200 170604 207098
rect 173604 679254 174204 710862
rect 191604 710478 192204 711440
rect 191604 710242 191786 710478
rect 192022 710242 192204 710478
rect 191604 710158 192204 710242
rect 191604 709922 191786 710158
rect 192022 709922 192204 710158
rect 188004 708598 188604 709560
rect 188004 708362 188186 708598
rect 188422 708362 188604 708598
rect 188004 708278 188604 708362
rect 188004 708042 188186 708278
rect 188422 708042 188604 708278
rect 184404 706718 185004 707680
rect 184404 706482 184586 706718
rect 184822 706482 185004 706718
rect 184404 706398 185004 706482
rect 184404 706162 184586 706398
rect 184822 706162 185004 706398
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 391254 174204 426698
rect 173604 391018 173786 391254
rect 174022 391018 174204 391254
rect 173604 390934 174204 391018
rect 173604 390698 173786 390934
rect 174022 390698 174204 390934
rect 173604 355254 174204 390698
rect 173604 355018 173786 355254
rect 174022 355018 174204 355254
rect 173604 354934 174204 355018
rect 173604 354698 173786 354934
rect 174022 354698 174204 354934
rect 173604 319254 174204 354698
rect 173604 319018 173786 319254
rect 174022 319018 174204 319254
rect 173604 318934 174204 319018
rect 173604 318698 173786 318934
rect 174022 318698 174204 318934
rect 173604 283254 174204 318698
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 200200 174204 210698
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 200200 181404 217898
rect 184404 690054 185004 706162
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 402054 185004 437498
rect 184404 401818 184586 402054
rect 184822 401818 185004 402054
rect 184404 401734 185004 401818
rect 184404 401498 184586 401734
rect 184822 401498 185004 401734
rect 184404 366054 185004 401498
rect 184404 365818 184586 366054
rect 184822 365818 185004 366054
rect 184404 365734 185004 365818
rect 184404 365498 184586 365734
rect 184822 365498 185004 365734
rect 184404 330054 185004 365498
rect 184404 329818 184586 330054
rect 184822 329818 185004 330054
rect 184404 329734 185004 329818
rect 184404 329498 184586 329734
rect 184822 329498 185004 329734
rect 184404 294054 185004 329498
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 200200 185004 221498
rect 188004 693654 188604 708042
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 405654 188604 441098
rect 188004 405418 188186 405654
rect 188422 405418 188604 405654
rect 188004 405334 188604 405418
rect 188004 405098 188186 405334
rect 188422 405098 188604 405334
rect 188004 369654 188604 405098
rect 188004 369418 188186 369654
rect 188422 369418 188604 369654
rect 188004 369334 188604 369418
rect 188004 369098 188186 369334
rect 188422 369098 188604 369334
rect 188004 333654 188604 369098
rect 188004 333418 188186 333654
rect 188422 333418 188604 333654
rect 188004 333334 188604 333418
rect 188004 333098 188186 333334
rect 188422 333098 188604 333334
rect 188004 297654 188604 333098
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 200200 188604 225098
rect 191604 697254 192204 709922
rect 209604 711418 210204 711440
rect 209604 711182 209786 711418
rect 210022 711182 210204 711418
rect 209604 711098 210204 711182
rect 209604 710862 209786 711098
rect 210022 710862 210204 711098
rect 206004 709538 206604 709560
rect 206004 709302 206186 709538
rect 206422 709302 206604 709538
rect 206004 709218 206604 709302
rect 206004 708982 206186 709218
rect 206422 708982 206604 709218
rect 202404 707658 203004 707680
rect 202404 707422 202586 707658
rect 202822 707422 203004 707658
rect 202404 707338 203004 707422
rect 202404 707102 202586 707338
rect 202822 707102 203004 707338
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 409254 192204 444698
rect 191604 409018 191786 409254
rect 192022 409018 192204 409254
rect 191604 408934 192204 409018
rect 191604 408698 191786 408934
rect 192022 408698 192204 408934
rect 191604 373254 192204 408698
rect 191604 373018 191786 373254
rect 192022 373018 192204 373254
rect 191604 372934 192204 373018
rect 191604 372698 191786 372934
rect 192022 372698 192204 372934
rect 191604 337254 192204 372698
rect 191604 337018 191786 337254
rect 192022 337018 192204 337254
rect 191604 336934 192204 337018
rect 191604 336698 191786 336934
rect 192022 336698 192204 336934
rect 191604 301254 192204 336698
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 200200 192204 228698
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 202404 672054 203004 707102
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 202404 560200 203004 563498
rect 206004 675654 206604 708982
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 560200 206604 567098
rect 209604 679254 210204 710862
rect 227604 710478 228204 711440
rect 227604 710242 227786 710478
rect 228022 710242 228204 710478
rect 227604 710158 228204 710242
rect 227604 709922 227786 710158
rect 228022 709922 228204 710158
rect 224004 708598 224604 709560
rect 224004 708362 224186 708598
rect 224422 708362 224604 708598
rect 224004 708278 224604 708362
rect 224004 708042 224186 708278
rect 224422 708042 224604 708278
rect 220404 706718 221004 707680
rect 220404 706482 220586 706718
rect 220822 706482 221004 706718
rect 220404 706398 221004 706482
rect 220404 706162 220586 706398
rect 220822 706162 221004 706398
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 560200 210204 570698
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 560200 217404 577898
rect 220404 690054 221004 706162
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198804 524454 199404 559898
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 203909 542454 204229 542476
rect 203909 542218 203951 542454
rect 204187 542218 204229 542454
rect 203909 542134 204229 542218
rect 203909 541898 203951 542134
rect 204187 541898 204229 542134
rect 203909 541876 204229 541898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 206875 524454 207195 524476
rect 206875 524218 206917 524454
rect 207153 524218 207195 524454
rect 206875 524134 207195 524218
rect 206875 523898 206917 524134
rect 207153 523898 207195 524134
rect 206875 523876 207195 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 202404 492054 203004 519800
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 409022 203004 419498
rect 206004 495654 206604 519800
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 409022 206604 423098
rect 209604 499254 210204 519800
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 409022 210204 426698
rect 216804 506454 217404 519800
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 409022 217404 433898
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 409022 221004 437498
rect 224004 693654 224604 708042
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 549654 224604 585098
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 409022 224604 441098
rect 227604 697254 228204 709922
rect 245604 711418 246204 711440
rect 245604 711182 245786 711418
rect 246022 711182 246204 711418
rect 245604 711098 246204 711182
rect 245604 710862 245786 711098
rect 246022 710862 246204 711098
rect 242004 709538 242604 709560
rect 242004 709302 242186 709538
rect 242422 709302 242604 709538
rect 242004 709218 242604 709302
rect 242004 708982 242186 709218
rect 242422 708982 242604 709218
rect 238404 707658 239004 707680
rect 238404 707422 238586 707658
rect 238822 707422 239004 707658
rect 238404 707338 239004 707422
rect 238404 707102 238586 707338
rect 238822 707102 239004 707338
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 553254 228204 588698
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 409022 228204 444698
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 234804 409022 235404 415898
rect 238404 672054 239004 707102
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 564054 239004 599498
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 420054 239004 455498
rect 238404 419818 238586 420054
rect 238822 419818 239004 420054
rect 238404 419734 239004 419818
rect 238404 419498 238586 419734
rect 238822 419498 239004 419734
rect 238404 409022 239004 419498
rect 242004 675654 242604 708982
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 567654 242604 603098
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 242004 495654 242604 531098
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 242004 423654 242604 459098
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 242004 409022 242604 423098
rect 245604 679254 246204 710862
rect 263604 710478 264204 711440
rect 263604 710242 263786 710478
rect 264022 710242 264204 710478
rect 263604 710158 264204 710242
rect 263604 709922 263786 710158
rect 264022 709922 264204 710158
rect 260004 708598 260604 709560
rect 260004 708362 260186 708598
rect 260422 708362 260604 708598
rect 260004 708278 260604 708362
rect 260004 708042 260186 708278
rect 260422 708042 260604 708278
rect 256404 706718 257004 707680
rect 256404 706482 256586 706718
rect 256822 706482 257004 706718
rect 256404 706398 257004 706482
rect 256404 706162 256586 706398
rect 256822 706162 257004 706398
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 571254 246204 606698
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 535254 246204 570698
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 245604 499254 246204 534698
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 245604 427254 246204 462698
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 245604 409022 246204 426698
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 252804 409022 253404 433898
rect 256404 690054 257004 706162
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 409022 257004 437498
rect 260004 693654 260604 708042
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 477654 260604 513098
rect 260004 477418 260186 477654
rect 260422 477418 260604 477654
rect 260004 477334 260604 477418
rect 260004 477098 260186 477334
rect 260422 477098 260604 477334
rect 260004 441654 260604 477098
rect 260004 441418 260186 441654
rect 260422 441418 260604 441654
rect 260004 441334 260604 441418
rect 260004 441098 260186 441334
rect 260422 441098 260604 441334
rect 260004 409022 260604 441098
rect 263604 697254 264204 709922
rect 281604 711418 282204 711440
rect 281604 711182 281786 711418
rect 282022 711182 282204 711418
rect 281604 711098 282204 711182
rect 281604 710862 281786 711098
rect 282022 710862 282204 711098
rect 278004 709538 278604 709560
rect 278004 709302 278186 709538
rect 278422 709302 278604 709538
rect 278004 709218 278604 709302
rect 278004 708982 278186 709218
rect 278422 708982 278604 709218
rect 274404 707658 275004 707680
rect 274404 707422 274586 707658
rect 274822 707422 275004 707658
rect 274404 707338 275004 707422
rect 274404 707102 274586 707338
rect 274822 707102 275004 707338
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 517254 264204 552698
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 481254 264204 516698
rect 263604 481018 263786 481254
rect 264022 481018 264204 481254
rect 263604 480934 264204 481018
rect 263604 480698 263786 480934
rect 264022 480698 264204 480934
rect 263604 445254 264204 480698
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 409022 264204 444698
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 274404 672054 275004 707102
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 271643 502348 271709 502349
rect 271643 502284 271644 502348
rect 271708 502284 271709 502348
rect 271643 502283 271709 502284
rect 271646 492693 271706 502283
rect 271643 492692 271709 492693
rect 271643 492628 271644 492692
rect 271708 492628 271709 492692
rect 271643 492627 271709 492628
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 204208 398454 204528 398476
rect 204208 398218 204250 398454
rect 204486 398218 204528 398454
rect 204208 398134 204528 398218
rect 204208 397898 204250 398134
rect 204486 397898 204528 398134
rect 204208 397876 204528 397898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 219568 380454 219888 380476
rect 219568 380218 219610 380454
rect 219846 380218 219888 380454
rect 219568 380134 219888 380218
rect 219568 379898 219610 380134
rect 219846 379898 219888 380134
rect 219568 379876 219888 379898
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 204208 362454 204528 362476
rect 204208 362218 204250 362454
rect 204486 362218 204528 362454
rect 204208 362134 204528 362218
rect 204208 361898 204250 362134
rect 204486 361898 204528 362134
rect 204208 361876 204528 361898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 219568 344454 219888 344476
rect 219568 344218 219610 344454
rect 219846 344218 219888 344454
rect 219568 344134 219888 344218
rect 219568 343898 219610 344134
rect 219846 343898 219888 344134
rect 219568 343876 219888 343898
rect 270804 344454 271404 379898
rect 270804 344218 270986 344454
rect 271222 344218 271404 344454
rect 270804 344134 271404 344218
rect 270804 343898 270986 344134
rect 271222 343898 271404 344134
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198804 200200 199404 235898
rect 202404 312054 203004 339800
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 202404 200200 203004 203498
rect 206004 315654 206604 339800
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 200200 206604 207098
rect 209604 319254 210204 339800
rect 209604 319018 209786 319254
rect 210022 319018 210204 319254
rect 209604 318934 210204 319018
rect 209604 318698 209786 318934
rect 210022 318698 210204 318934
rect 209604 283254 210204 318698
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 200200 210204 210698
rect 216804 326454 217404 339800
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 200200 217404 217898
rect 220404 330054 221004 339800
rect 220404 329818 220586 330054
rect 220822 329818 221004 330054
rect 220404 329734 221004 329818
rect 220404 329498 220586 329734
rect 220822 329498 221004 329734
rect 220404 294054 221004 329498
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 200200 221004 221498
rect 224004 333654 224604 339800
rect 224004 333418 224186 333654
rect 224422 333418 224604 333654
rect 224004 333334 224604 333418
rect 224004 333098 224186 333334
rect 224422 333098 224604 333334
rect 224004 297654 224604 333098
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 200200 224604 225098
rect 227604 337254 228204 339800
rect 227604 337018 227786 337254
rect 228022 337018 228204 337254
rect 227604 336934 228204 337018
rect 227604 336698 227786 336934
rect 228022 336698 228204 336934
rect 227604 301254 228204 336698
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 200200 228204 228698
rect 234804 308454 235404 339800
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200200 235404 235898
rect 238404 312054 239004 339800
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 200200 239004 203498
rect 242004 315654 242604 339800
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 200200 242604 207098
rect 245604 319254 246204 339800
rect 245604 319018 245786 319254
rect 246022 319018 246204 319254
rect 245604 318934 246204 319018
rect 245604 318698 245786 318934
rect 246022 318698 246204 318934
rect 245604 283254 246204 318698
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 200200 246204 210698
rect 252804 326454 253404 339800
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 200200 253404 217898
rect 256404 330054 257004 339800
rect 256404 329818 256586 330054
rect 256822 329818 257004 330054
rect 256404 329734 257004 329818
rect 256404 329498 256586 329734
rect 256822 329498 257004 329734
rect 256404 294054 257004 329498
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 200200 257004 221498
rect 260004 333654 260604 339800
rect 260004 333418 260186 333654
rect 260422 333418 260604 333654
rect 260004 333334 260604 333418
rect 260004 333098 260186 333334
rect 260422 333098 260604 333334
rect 260004 297654 260604 333098
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 200200 260604 225098
rect 263604 337254 264204 339800
rect 263604 337018 263786 337254
rect 264022 337018 264204 337254
rect 263604 336934 264204 337018
rect 263604 336698 263786 336934
rect 264022 336698 264204 336934
rect 263604 301254 264204 336698
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 200200 264204 228698
rect 270804 308454 271404 343898
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 270804 200200 271404 235898
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 420054 275004 455498
rect 274404 419818 274586 420054
rect 274822 419818 275004 420054
rect 274404 419734 275004 419818
rect 274404 419498 274586 419734
rect 274822 419498 275004 419734
rect 274404 384054 275004 419498
rect 274404 383818 274586 384054
rect 274822 383818 275004 384054
rect 274404 383734 275004 383818
rect 274404 383498 274586 383734
rect 274822 383498 275004 383734
rect 274404 348054 275004 383498
rect 274404 347818 274586 348054
rect 274822 347818 275004 348054
rect 274404 347734 275004 347818
rect 274404 347498 274586 347734
rect 274822 347498 275004 347734
rect 274404 312054 275004 347498
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 200200 275004 203498
rect 278004 675654 278604 708982
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 459654 278604 495098
rect 278004 459418 278186 459654
rect 278422 459418 278604 459654
rect 278004 459334 278604 459418
rect 278004 459098 278186 459334
rect 278422 459098 278604 459334
rect 278004 423654 278604 459098
rect 278004 423418 278186 423654
rect 278422 423418 278604 423654
rect 278004 423334 278604 423418
rect 278004 423098 278186 423334
rect 278422 423098 278604 423334
rect 278004 387654 278604 423098
rect 278004 387418 278186 387654
rect 278422 387418 278604 387654
rect 278004 387334 278604 387418
rect 278004 387098 278186 387334
rect 278422 387098 278604 387334
rect 278004 351654 278604 387098
rect 278004 351418 278186 351654
rect 278422 351418 278604 351654
rect 278004 351334 278604 351418
rect 278004 351098 278186 351334
rect 278422 351098 278604 351334
rect 278004 315654 278604 351098
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 281604 679254 282204 710862
rect 299604 710478 300204 711440
rect 299604 710242 299786 710478
rect 300022 710242 300204 710478
rect 299604 710158 300204 710242
rect 299604 709922 299786 710158
rect 300022 709922 300204 710158
rect 296004 708598 296604 709560
rect 296004 708362 296186 708598
rect 296422 708362 296604 708598
rect 296004 708278 296604 708362
rect 296004 708042 296186 708278
rect 296422 708042 296604 708278
rect 292404 706718 293004 707680
rect 292404 706482 292586 706718
rect 292822 706482 293004 706718
rect 292404 706398 293004 706482
rect 292404 706162 292586 706398
rect 292822 706162 293004 706398
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 463254 282204 498698
rect 281604 463018 281786 463254
rect 282022 463018 282204 463254
rect 281604 462934 282204 463018
rect 281604 462698 281786 462934
rect 282022 462698 282204 462934
rect 281604 427254 282204 462698
rect 281604 427018 281786 427254
rect 282022 427018 282204 427254
rect 281604 426934 282204 427018
rect 281604 426698 281786 426934
rect 282022 426698 282204 426934
rect 281604 391254 282204 426698
rect 281604 391018 281786 391254
rect 282022 391018 282204 391254
rect 281604 390934 282204 391018
rect 281604 390698 281786 390934
rect 282022 390698 282204 390934
rect 281604 355254 282204 390698
rect 281604 355018 281786 355254
rect 282022 355018 282204 355254
rect 281604 354934 282204 355018
rect 281604 354698 281786 354934
rect 282022 354698 282204 354934
rect 281604 319254 282204 354698
rect 281604 319018 281786 319254
rect 282022 319018 282204 319254
rect 281604 318934 282204 319018
rect 281604 318698 281786 318934
rect 282022 318698 282204 318934
rect 281604 283254 282204 318698
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281211 260812 281277 260813
rect 281211 260748 281212 260812
rect 281276 260748 281277 260812
rect 281211 260747 281277 260748
rect 281214 251293 281274 260747
rect 281211 251292 281277 251293
rect 281211 251228 281212 251292
rect 281276 251228 281277 251292
rect 281211 251227 281277 251228
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 200200 278604 207098
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 200200 282204 210698
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 200200 289404 217898
rect 292404 690054 293004 706162
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 200200 293004 221498
rect 296004 693654 296604 708042
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 299604 697254 300204 709922
rect 317604 711418 318204 711440
rect 317604 711182 317786 711418
rect 318022 711182 318204 711418
rect 317604 711098 318204 711182
rect 317604 710862 317786 711098
rect 318022 710862 318204 711098
rect 314004 709538 314604 709560
rect 314004 709302 314186 709538
rect 314422 709302 314604 709538
rect 314004 709218 314604 709302
rect 314004 708982 314186 709218
rect 314422 708982 314604 709218
rect 310404 707658 311004 707680
rect 310404 707422 310586 707658
rect 310822 707422 311004 707658
rect 310404 707338 311004 707422
rect 310404 707102 310586 707338
rect 310822 707102 311004 707338
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 580211 300204 588698
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 580211 307404 595898
rect 310404 672054 311004 707102
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 580211 311004 599498
rect 314004 675654 314604 708982
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 580211 314604 603098
rect 317604 679254 318204 710862
rect 335604 710478 336204 711440
rect 335604 710242 335786 710478
rect 336022 710242 336204 710478
rect 335604 710158 336204 710242
rect 335604 709922 335786 710158
rect 336022 709922 336204 710158
rect 332004 708598 332604 709560
rect 332004 708362 332186 708598
rect 332422 708362 332604 708598
rect 332004 708278 332604 708362
rect 332004 708042 332186 708278
rect 332422 708042 332604 708278
rect 328404 706718 329004 707680
rect 328404 706482 328586 706718
rect 328822 706482 329004 706718
rect 328404 706398 329004 706482
rect 328404 706162 328586 706398
rect 328822 706162 329004 706398
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 580211 318204 606698
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 580211 325404 613898
rect 328404 690054 329004 706162
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 580211 329004 581498
rect 332004 693654 332604 708042
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 580211 332604 585098
rect 335604 697254 336204 709922
rect 353604 711418 354204 711440
rect 353604 711182 353786 711418
rect 354022 711182 354204 711418
rect 353604 711098 354204 711182
rect 353604 710862 353786 711098
rect 354022 710862 354204 711098
rect 350004 709538 350604 709560
rect 350004 709302 350186 709538
rect 350422 709302 350604 709538
rect 350004 709218 350604 709302
rect 350004 708982 350186 709218
rect 350422 708982 350604 709218
rect 346404 707658 347004 707680
rect 346404 707422 346586 707658
rect 346822 707422 347004 707658
rect 346404 707338 347004 707422
rect 346404 707102 346586 707338
rect 346822 707102 347004 707338
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 580211 336204 588698
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 580211 343404 595898
rect 346404 672054 347004 707102
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 580211 347004 599498
rect 350004 675654 350604 708982
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 580211 350604 603098
rect 353604 679254 354204 710862
rect 371604 710478 372204 711440
rect 371604 710242 371786 710478
rect 372022 710242 372204 710478
rect 371604 710158 372204 710242
rect 371604 709922 371786 710158
rect 372022 709922 372204 710158
rect 368004 708598 368604 709560
rect 368004 708362 368186 708598
rect 368422 708362 368604 708598
rect 368004 708278 368604 708362
rect 368004 708042 368186 708278
rect 368422 708042 368604 708278
rect 364404 706718 365004 707680
rect 364404 706482 364586 706718
rect 364822 706482 365004 706718
rect 364404 706398 365004 706482
rect 364404 706162 364586 706398
rect 364822 706162 365004 706398
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 580211 354204 606698
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 580211 361404 613898
rect 364404 690054 365004 706162
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 580211 365004 581498
rect 368004 693654 368604 708042
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 580211 368604 585098
rect 371604 697254 372204 709922
rect 389604 711418 390204 711440
rect 389604 711182 389786 711418
rect 390022 711182 390204 711418
rect 389604 711098 390204 711182
rect 389604 710862 389786 711098
rect 390022 710862 390204 711098
rect 386004 709538 386604 709560
rect 386004 709302 386186 709538
rect 386422 709302 386604 709538
rect 386004 709218 386604 709302
rect 386004 708982 386186 709218
rect 386422 708982 386604 709218
rect 382404 707658 383004 707680
rect 382404 707422 382586 707658
rect 382822 707422 383004 707658
rect 382404 707338 383004 707422
rect 382404 707102 382586 707338
rect 382822 707102 383004 707338
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 580211 372204 588698
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 319568 560454 319888 560476
rect 319568 560218 319610 560454
rect 319846 560218 319888 560454
rect 319568 560134 319888 560218
rect 319568 559898 319610 560134
rect 319846 559898 319888 560134
rect 319568 559876 319888 559898
rect 378804 560454 379404 595898
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 304208 542454 304528 542476
rect 304208 542218 304250 542454
rect 304486 542218 304528 542454
rect 304208 542134 304528 542218
rect 304208 541898 304250 542134
rect 304486 541898 304528 542134
rect 304208 541876 304528 541898
rect 319568 524454 319888 524476
rect 319568 524218 319610 524454
rect 319846 524218 319888 524454
rect 319568 524134 319888 524218
rect 319568 523898 319610 524134
rect 319846 523898 319888 524134
rect 319568 523876 319888 523898
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 304208 506454 304528 506476
rect 304208 506218 304250 506454
rect 304486 506218 304528 506454
rect 304208 506134 304528 506218
rect 304208 505898 304250 506134
rect 304486 505898 304528 506134
rect 304208 505876 304528 505898
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 200200 296604 225098
rect 299604 481254 300204 499800
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299604 301254 300204 336698
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 200200 300204 228698
rect 306804 488454 307404 499800
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200200 307404 235898
rect 310404 492054 311004 499800
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 200200 311004 203498
rect 314004 495654 314604 499800
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 200200 314604 207098
rect 317604 499254 318204 499800
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 200200 318204 210698
rect 324804 470454 325404 499800
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 200200 325404 217898
rect 328404 474054 329004 499800
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 294054 329004 329498
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 200200 329004 221498
rect 332004 477654 332604 499800
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 297654 332604 333098
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 200200 332604 225098
rect 335604 481254 336204 499800
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 335604 301254 336204 336698
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 200200 336204 228698
rect 342804 488454 343404 499800
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200200 343404 235898
rect 346404 492054 347004 499800
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 384054 347004 419498
rect 346404 383818 346586 384054
rect 346822 383818 347004 384054
rect 346404 383734 347004 383818
rect 346404 383498 346586 383734
rect 346822 383498 347004 383734
rect 346404 348054 347004 383498
rect 346404 347818 346586 348054
rect 346822 347818 347004 348054
rect 346404 347734 347004 347818
rect 346404 347498 346586 347734
rect 346822 347498 347004 347734
rect 346404 312054 347004 347498
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 200200 347004 203498
rect 350004 495654 350604 499800
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 387654 350604 423098
rect 350004 387418 350186 387654
rect 350422 387418 350604 387654
rect 350004 387334 350604 387418
rect 350004 387098 350186 387334
rect 350422 387098 350604 387334
rect 350004 351654 350604 387098
rect 350004 351418 350186 351654
rect 350422 351418 350604 351654
rect 350004 351334 350604 351418
rect 350004 351098 350186 351334
rect 350422 351098 350604 351334
rect 350004 315654 350604 351098
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 200200 350604 207098
rect 353604 499254 354204 499800
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 391254 354204 426698
rect 353604 391018 353786 391254
rect 354022 391018 354204 391254
rect 353604 390934 354204 391018
rect 353604 390698 353786 390934
rect 354022 390698 354204 390934
rect 353604 355254 354204 390698
rect 353604 355018 353786 355254
rect 354022 355018 354204 355254
rect 353604 354934 354204 355018
rect 353604 354698 353786 354934
rect 354022 354698 354204 354934
rect 353604 319254 354204 354698
rect 353604 319018 353786 319254
rect 354022 319018 354204 319254
rect 353604 318934 354204 319018
rect 353604 318698 353786 318934
rect 354022 318698 354204 318934
rect 353604 283254 354204 318698
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 200200 354204 210698
rect 360804 470454 361404 499800
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 200200 361404 217898
rect 364404 474054 365004 499800
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 402054 365004 437498
rect 364404 401818 364586 402054
rect 364822 401818 365004 402054
rect 364404 401734 365004 401818
rect 364404 401498 364586 401734
rect 364822 401498 365004 401734
rect 364404 366054 365004 401498
rect 364404 365818 364586 366054
rect 364822 365818 365004 366054
rect 364404 365734 365004 365818
rect 364404 365498 364586 365734
rect 364822 365498 365004 365734
rect 364404 330054 365004 365498
rect 364404 329818 364586 330054
rect 364822 329818 365004 330054
rect 364404 329734 365004 329818
rect 364404 329498 364586 329734
rect 364822 329498 365004 329734
rect 364404 294054 365004 329498
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 200200 365004 221498
rect 368004 477654 368604 499800
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 405654 368604 441098
rect 368004 405418 368186 405654
rect 368422 405418 368604 405654
rect 368004 405334 368604 405418
rect 368004 405098 368186 405334
rect 368422 405098 368604 405334
rect 368004 369654 368604 405098
rect 368004 369418 368186 369654
rect 368422 369418 368604 369654
rect 368004 369334 368604 369418
rect 368004 369098 368186 369334
rect 368422 369098 368604 369334
rect 368004 333654 368604 369098
rect 368004 333418 368186 333654
rect 368422 333418 368604 333654
rect 368004 333334 368604 333418
rect 368004 333098 368186 333334
rect 368422 333098 368604 333334
rect 368004 297654 368604 333098
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 200200 368604 225098
rect 371604 481254 372204 499800
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 409254 372204 444698
rect 371604 409018 371786 409254
rect 372022 409018 372204 409254
rect 371604 408934 372204 409018
rect 371604 408698 371786 408934
rect 372022 408698 372204 408934
rect 371604 373254 372204 408698
rect 371604 373018 371786 373254
rect 372022 373018 372204 373254
rect 371604 372934 372204 373018
rect 371604 372698 371786 372934
rect 372022 372698 372204 372934
rect 371604 337254 372204 372698
rect 371604 337018 371786 337254
rect 372022 337018 372204 337254
rect 371604 336934 372204 337018
rect 371604 336698 371786 336934
rect 372022 336698 372204 336934
rect 371604 301254 372204 336698
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 200200 372204 228698
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200200 379404 235898
rect 382404 672054 383004 707102
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 384054 383004 419498
rect 382404 383818 382586 384054
rect 382822 383818 383004 384054
rect 382404 383734 383004 383818
rect 382404 383498 382586 383734
rect 382822 383498 383004 383734
rect 386004 675654 386604 708982
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 387654 386604 423098
rect 386004 387418 386186 387654
rect 386422 387418 386604 387654
rect 386004 387334 386604 387418
rect 386004 387098 386186 387334
rect 386422 387098 386604 387334
rect 386004 383619 386604 387098
rect 389604 679254 390204 710862
rect 407604 710478 408204 711440
rect 407604 710242 407786 710478
rect 408022 710242 408204 710478
rect 407604 710158 408204 710242
rect 407604 709922 407786 710158
rect 408022 709922 408204 710158
rect 404004 708598 404604 709560
rect 404004 708362 404186 708598
rect 404422 708362 404604 708598
rect 404004 708278 404604 708362
rect 404004 708042 404186 708278
rect 404422 708042 404604 708278
rect 400404 706718 401004 707680
rect 400404 706482 400586 706718
rect 400822 706482 401004 706718
rect 400404 706398 401004 706482
rect 400404 706162 400586 706398
rect 400822 706162 401004 706398
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 391254 390204 426698
rect 389604 391018 389786 391254
rect 390022 391018 390204 391254
rect 389604 390934 390204 391018
rect 389604 390698 389786 390934
rect 390022 390698 390204 390934
rect 389604 383619 390204 390698
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 383619 397404 397898
rect 400404 690054 401004 706162
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 383619 401004 401498
rect 404004 693654 404604 708042
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 383619 404604 405098
rect 407604 697254 408204 709922
rect 425604 711418 426204 711440
rect 425604 711182 425786 711418
rect 426022 711182 426204 711418
rect 425604 711098 426204 711182
rect 425604 710862 425786 711098
rect 426022 710862 426204 711098
rect 422004 709538 422604 709560
rect 422004 709302 422186 709538
rect 422422 709302 422604 709538
rect 422004 709218 422604 709302
rect 422004 708982 422186 709218
rect 422422 708982 422604 709218
rect 418404 707658 419004 707680
rect 418404 707422 418586 707658
rect 418822 707422 419004 707658
rect 418404 707338 419004 707422
rect 418404 707102 418586 707338
rect 418822 707102 419004 707338
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 383619 408204 408698
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 383619 415404 415898
rect 418404 672054 419004 707102
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 382404 348054 383004 383498
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 394604 380454 394924 380476
rect 394604 380218 394646 380454
rect 394882 380218 394924 380454
rect 394604 380134 394924 380218
rect 394604 379898 394646 380134
rect 394882 379898 394924 380134
rect 394604 379876 394924 379898
rect 389774 362454 390094 362476
rect 389774 362218 389816 362454
rect 390052 362218 390094 362454
rect 389774 362134 390094 362218
rect 389774 361898 389816 362134
rect 390052 361898 390094 362134
rect 389774 361876 390094 361898
rect 382404 347818 382586 348054
rect 382822 347818 383004 348054
rect 382404 347734 383004 347818
rect 382404 347498 382586 347734
rect 382822 347498 383004 347734
rect 382404 312054 383004 347498
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 200200 383004 203498
rect 386004 315654 386604 349800
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 200200 386604 207098
rect 389604 319254 390204 349800
rect 389604 319018 389786 319254
rect 390022 319018 390204 319254
rect 389604 318934 390204 319018
rect 389604 318698 389786 318934
rect 390022 318698 390204 318934
rect 389604 283254 390204 318698
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 200200 390204 210698
rect 396804 326454 397404 349800
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 200200 397404 217898
rect 400404 330054 401004 349800
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 200200 401004 221498
rect 404004 333654 404604 349800
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 297654 404604 333098
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 200200 404604 225098
rect 407604 337254 408204 349800
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 301254 408204 336698
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 200200 408204 228698
rect 414804 344454 415404 349800
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200200 415404 235898
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 200200 419004 203498
rect 422004 675654 422604 708982
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 200200 422604 207098
rect 425604 679254 426204 710862
rect 443604 710478 444204 711440
rect 443604 710242 443786 710478
rect 444022 710242 444204 710478
rect 443604 710158 444204 710242
rect 443604 709922 443786 710158
rect 444022 709922 444204 710158
rect 440004 708598 440604 709560
rect 440004 708362 440186 708598
rect 440422 708362 440604 708598
rect 440004 708278 440604 708362
rect 440004 708042 440186 708278
rect 440422 708042 440604 708278
rect 436404 706718 437004 707680
rect 436404 706482 436586 706718
rect 436822 706482 437004 706718
rect 436404 706398 437004 706482
rect 436404 706162 436586 706398
rect 436822 706162 437004 706398
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 200200 426204 210698
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 200200 433404 217898
rect 436404 690054 437004 706162
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 133091 200156 133157 200157
rect 133091 200092 133092 200156
rect 133156 200092 133157 200156
rect 133091 200091 133157 200092
rect 132907 196076 132973 196077
rect 132907 196012 132908 196076
rect 132972 196012 132973 196076
rect 132907 196011 132973 196012
rect 132910 195941 132970 196011
rect 132907 195940 132973 195941
rect 132907 195876 132908 195940
rect 132972 195876 132973 195940
rect 132907 195875 132973 195876
rect 132907 185468 132973 185469
rect 132907 185404 132908 185468
rect 132972 185404 132973 185468
rect 132907 185403 132973 185404
rect 132910 182341 132970 185403
rect 133094 184925 133154 200091
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 133091 184924 133157 184925
rect 133091 184860 133092 184924
rect 133156 184860 133157 184924
rect 133091 184859 133157 184860
rect 138208 182454 138528 182476
rect 132907 182340 132973 182341
rect 132907 182276 132908 182340
rect 132972 182276 132973 182340
rect 132907 182275 132973 182276
rect 138208 182218 138250 182454
rect 138486 182218 138528 182454
rect 138208 182134 138528 182218
rect 138208 181898 138250 182134
rect 138486 181898 138528 182134
rect 138208 181876 138528 181898
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 128491 154868 128557 154869
rect 128491 154804 128492 154868
rect 128556 154804 128557 154868
rect 128491 154803 128557 154804
rect 128494 154597 128554 154803
rect 128491 154596 128557 154597
rect 128491 154532 128492 154596
rect 128556 154532 128557 154596
rect 128491 154531 128557 154532
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 130404 132054 131004 167498
rect 153568 164454 153888 164476
rect 153568 164218 153610 164454
rect 153846 164218 153888 164454
rect 153568 164134 153888 164218
rect 153568 163898 153610 164134
rect 153846 163898 153888 164134
rect 153568 163876 153888 163898
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 132171 147796 132237 147797
rect 132171 147732 132172 147796
rect 132236 147732 132237 147796
rect 132171 147731 132237 147732
rect 132174 147525 132234 147731
rect 132171 147524 132237 147525
rect 132171 147460 132172 147524
rect 132236 147460 132237 147524
rect 132171 147459 132237 147460
rect 138208 146454 138528 146476
rect 138208 146218 138250 146454
rect 138486 146218 138528 146454
rect 138208 146134 138528 146218
rect 138208 145898 138250 146134
rect 138486 145898 138528 146134
rect 138208 145876 138528 145898
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 153568 128454 153888 128476
rect 153568 128218 153610 128454
rect 153846 128218 153888 128454
rect 153568 128134 153888 128218
rect 153568 127898 153610 128134
rect 153846 127898 153888 128134
rect 153568 127876 153888 127898
rect 133827 118148 133893 118149
rect 133827 118084 133828 118148
rect 133892 118084 133893 118148
rect 133827 118083 133893 118084
rect 133830 117605 133890 118083
rect 133827 117604 133893 117605
rect 133827 117540 133828 117604
rect 133892 117540 133893 117604
rect 133827 117539 133893 117540
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3166 131004 23498
rect 130404 -3402 130586 -3166
rect 130822 -3402 131004 -3166
rect 130404 -3486 131004 -3402
rect 130404 -3722 130586 -3486
rect 130822 -3722 131004 -3486
rect 130404 -3744 131004 -3722
rect 134004 99654 134604 119800
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -5046 134604 27098
rect 134004 -5282 134186 -5046
rect 134422 -5282 134604 -5046
rect 134004 -5366 134604 -5282
rect 134004 -5602 134186 -5366
rect 134422 -5602 134604 -5366
rect 134004 -5624 134604 -5602
rect 137604 103254 138204 119800
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 144804 110454 145404 119800
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 140819 60892 140885 60893
rect 140819 60828 140820 60892
rect 140884 60828 140885 60892
rect 140819 60827 140885 60828
rect 140822 55317 140882 60827
rect 140819 55316 140885 55317
rect 140819 55252 140820 55316
rect 140884 55252 140885 55316
rect 140819 55251 140885 55252
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6222 119786 -5986
rect 120022 -6222 120204 -5986
rect 119604 -6306 120204 -6222
rect 119604 -6542 119786 -6306
rect 120022 -6542 120204 -6306
rect 119604 -7504 120204 -6542
rect 137604 -6926 138204 30698
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 148404 114054 149004 119800
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2226 149004 5498
rect 148404 -2462 148586 -2226
rect 148822 -2462 149004 -2226
rect 148404 -2546 149004 -2462
rect 148404 -2782 148586 -2546
rect 148822 -2782 149004 -2546
rect 148404 -3744 149004 -2782
rect 152004 117654 152604 119800
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4106 152604 9098
rect 152004 -4342 152186 -4106
rect 152422 -4342 152604 -4106
rect 152004 -4426 152604 -4342
rect 152004 -4662 152186 -4426
rect 152422 -4662 152604 -4426
rect 152004 -5624 152604 -4662
rect 155604 85254 156204 119800
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7162 137786 -6926
rect 138022 -7162 138204 -6926
rect 137604 -7246 138204 -7162
rect 137604 -7482 137786 -7246
rect 138022 -7482 138204 -7246
rect 137604 -7504 138204 -7482
rect 155604 -5986 156204 12698
rect 162804 92454 163404 119800
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 166404 96054 167004 119800
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3166 167004 23498
rect 166404 -3402 166586 -3166
rect 166822 -3402 167004 -3166
rect 166404 -3486 167004 -3402
rect 166404 -3722 166586 -3486
rect 166822 -3722 167004 -3486
rect 166404 -3744 167004 -3722
rect 170004 99654 170604 119800
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -5046 170604 27098
rect 170004 -5282 170186 -5046
rect 170422 -5282 170604 -5046
rect 170004 -5366 170604 -5282
rect 170004 -5602 170186 -5366
rect 170422 -5602 170604 -5366
rect 170004 -5624 170604 -5602
rect 173604 103254 174204 119800
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6222 155786 -5986
rect 156022 -6222 156204 -5986
rect 155604 -6306 156204 -6222
rect 155604 -6542 155786 -6306
rect 156022 -6542 156204 -6306
rect 155604 -7504 156204 -6542
rect 173604 -6926 174204 30698
rect 180804 110454 181404 119800
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 184404 114054 185004 119800
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2226 185004 5498
rect 184404 -2462 184586 -2226
rect 184822 -2462 185004 -2226
rect 184404 -2546 185004 -2462
rect 184404 -2782 184586 -2546
rect 184822 -2782 185004 -2546
rect 184404 -3744 185004 -2782
rect 188004 117654 188604 119800
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4106 188604 9098
rect 188004 -4342 188186 -4106
rect 188422 -4342 188604 -4106
rect 188004 -4426 188604 -4342
rect 188004 -4662 188186 -4426
rect 188422 -4662 188604 -4426
rect 188004 -5624 188604 -4662
rect 191604 85254 192204 119800
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7162 173786 -6926
rect 174022 -7162 174204 -6926
rect 173604 -7246 174204 -7162
rect 173604 -7482 173786 -7246
rect 174022 -7482 174204 -7246
rect 173604 -7504 174204 -7482
rect 191604 -5986 192204 12698
rect 198804 92454 199404 119800
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 202404 96054 203004 119800
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3166 203004 23498
rect 202404 -3402 202586 -3166
rect 202822 -3402 203004 -3166
rect 202404 -3486 203004 -3402
rect 202404 -3722 202586 -3486
rect 202822 -3722 203004 -3486
rect 202404 -3744 203004 -3722
rect 206004 99654 206604 119800
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -5046 206604 27098
rect 206004 -5282 206186 -5046
rect 206422 -5282 206604 -5046
rect 206004 -5366 206604 -5282
rect 206004 -5602 206186 -5366
rect 206422 -5602 206604 -5366
rect 206004 -5624 206604 -5602
rect 209604 103254 210204 119800
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6222 191786 -5986
rect 192022 -6222 192204 -5986
rect 191604 -6306 192204 -6222
rect 191604 -6542 191786 -6306
rect 192022 -6542 192204 -6306
rect 191604 -7504 192204 -6542
rect 209604 -6926 210204 30698
rect 216804 110454 217404 119800
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 220404 114054 221004 119800
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2226 221004 5498
rect 220404 -2462 220586 -2226
rect 220822 -2462 221004 -2226
rect 220404 -2546 221004 -2462
rect 220404 -2782 220586 -2546
rect 220822 -2782 221004 -2546
rect 220404 -3744 221004 -2782
rect 224004 117654 224604 119800
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4106 224604 9098
rect 224004 -4342 224186 -4106
rect 224422 -4342 224604 -4106
rect 224004 -4426 224604 -4342
rect 224004 -4662 224186 -4426
rect 224422 -4662 224604 -4426
rect 224004 -5624 224604 -4662
rect 227604 85254 228204 119800
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7162 209786 -6926
rect 210022 -7162 210204 -6926
rect 209604 -7246 210204 -7162
rect 209604 -7482 209786 -7246
rect 210022 -7482 210204 -7246
rect 209604 -7504 210204 -7482
rect 227604 -5986 228204 12698
rect 234804 92454 235404 119800
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 238404 96054 239004 119800
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3166 239004 23498
rect 238404 -3402 238586 -3166
rect 238822 -3402 239004 -3166
rect 238404 -3486 239004 -3402
rect 238404 -3722 238586 -3486
rect 238822 -3722 239004 -3486
rect 238404 -3744 239004 -3722
rect 242004 99654 242604 119800
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -5046 242604 27098
rect 242004 -5282 242186 -5046
rect 242422 -5282 242604 -5046
rect 242004 -5366 242604 -5282
rect 242004 -5602 242186 -5366
rect 242422 -5602 242604 -5366
rect 242004 -5624 242604 -5602
rect 245604 103254 246204 119800
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6222 227786 -5986
rect 228022 -6222 228204 -5986
rect 227604 -6306 228204 -6222
rect 227604 -6542 227786 -6306
rect 228022 -6542 228204 -6306
rect 227604 -7504 228204 -6542
rect 245604 -6926 246204 30698
rect 252804 110454 253404 119800
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 256404 114054 257004 119800
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2226 257004 5498
rect 256404 -2462 256586 -2226
rect 256822 -2462 257004 -2226
rect 256404 -2546 257004 -2462
rect 256404 -2782 256586 -2546
rect 256822 -2782 257004 -2546
rect 256404 -3744 257004 -2782
rect 260004 117654 260604 119800
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4106 260604 9098
rect 260004 -4342 260186 -4106
rect 260422 -4342 260604 -4106
rect 260004 -4426 260604 -4342
rect 260004 -4662 260186 -4426
rect 260422 -4662 260604 -4426
rect 260004 -5624 260604 -4662
rect 263604 85254 264204 119800
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7162 245786 -6926
rect 246022 -7162 246204 -6926
rect 245604 -7246 246204 -7162
rect 245604 -7482 245786 -7246
rect 246022 -7482 246204 -7246
rect 245604 -7504 246204 -7482
rect 263604 -5986 264204 12698
rect 270804 92454 271404 119800
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 274404 96054 275004 119800
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3166 275004 23498
rect 274404 -3402 274586 -3166
rect 274822 -3402 275004 -3166
rect 274404 -3486 275004 -3402
rect 274404 -3722 274586 -3486
rect 274822 -3722 275004 -3486
rect 274404 -3744 275004 -3722
rect 278004 99654 278604 119800
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -5046 278604 27098
rect 278004 -5282 278186 -5046
rect 278422 -5282 278604 -5046
rect 278004 -5366 278604 -5282
rect 278004 -5602 278186 -5366
rect 278422 -5602 278604 -5366
rect 278004 -5624 278604 -5602
rect 281604 103254 282204 119800
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6222 263786 -5986
rect 264022 -6222 264204 -5986
rect 263604 -6306 264204 -6222
rect 263604 -6542 263786 -6306
rect 264022 -6542 264204 -6306
rect 263604 -7504 264204 -6542
rect 281604 -6926 282204 30698
rect 288804 110454 289404 119800
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 292404 114054 293004 119800
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2226 293004 5498
rect 292404 -2462 292586 -2226
rect 292822 -2462 293004 -2226
rect 292404 -2546 293004 -2462
rect 292404 -2782 292586 -2546
rect 292822 -2782 293004 -2546
rect 292404 -3744 293004 -2782
rect 296004 117654 296604 119800
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4106 296604 9098
rect 296004 -4342 296186 -4106
rect 296422 -4342 296604 -4106
rect 296004 -4426 296604 -4342
rect 296004 -4662 296186 -4426
rect 296422 -4662 296604 -4426
rect 296004 -5624 296604 -4662
rect 299604 85254 300204 119800
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7162 281786 -6926
rect 282022 -7162 282204 -6926
rect 281604 -7246 282204 -7162
rect 281604 -7482 281786 -7246
rect 282022 -7482 282204 -7246
rect 281604 -7504 282204 -7482
rect 299604 -5986 300204 12698
rect 306804 92454 307404 119800
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 310404 96054 311004 119800
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3166 311004 23498
rect 310404 -3402 310586 -3166
rect 310822 -3402 311004 -3166
rect 310404 -3486 311004 -3402
rect 310404 -3722 310586 -3486
rect 310822 -3722 311004 -3486
rect 310404 -3744 311004 -3722
rect 314004 99654 314604 119800
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -5046 314604 27098
rect 314004 -5282 314186 -5046
rect 314422 -5282 314604 -5046
rect 314004 -5366 314604 -5282
rect 314004 -5602 314186 -5366
rect 314422 -5602 314604 -5366
rect 314004 -5624 314604 -5602
rect 317604 103254 318204 119800
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6222 299786 -5986
rect 300022 -6222 300204 -5986
rect 299604 -6306 300204 -6222
rect 299604 -6542 299786 -6306
rect 300022 -6542 300204 -6306
rect 299604 -7504 300204 -6542
rect 317604 -6926 318204 30698
rect 324804 110454 325404 119800
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 328404 114054 329004 119800
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2226 329004 5498
rect 328404 -2462 328586 -2226
rect 328822 -2462 329004 -2226
rect 328404 -2546 329004 -2462
rect 328404 -2782 328586 -2546
rect 328822 -2782 329004 -2546
rect 328404 -3744 329004 -2782
rect 332004 117654 332604 119800
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4106 332604 9098
rect 332004 -4342 332186 -4106
rect 332422 -4342 332604 -4106
rect 332004 -4426 332604 -4342
rect 332004 -4662 332186 -4426
rect 332422 -4662 332604 -4426
rect 332004 -5624 332604 -4662
rect 335604 85254 336204 119800
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7162 317786 -6926
rect 318022 -7162 318204 -6926
rect 317604 -7246 318204 -7162
rect 317604 -7482 317786 -7246
rect 318022 -7482 318204 -7246
rect 317604 -7504 318204 -7482
rect 335604 -5986 336204 12698
rect 342804 92454 343404 119800
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 346404 96054 347004 119800
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3166 347004 23498
rect 346404 -3402 346586 -3166
rect 346822 -3402 347004 -3166
rect 346404 -3486 347004 -3402
rect 346404 -3722 346586 -3486
rect 346822 -3722 347004 -3486
rect 346404 -3744 347004 -3722
rect 350004 99654 350604 119800
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -5046 350604 27098
rect 350004 -5282 350186 -5046
rect 350422 -5282 350604 -5046
rect 350004 -5366 350604 -5282
rect 350004 -5602 350186 -5366
rect 350422 -5602 350604 -5366
rect 350004 -5624 350604 -5602
rect 353604 103254 354204 119800
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6222 335786 -5986
rect 336022 -6222 336204 -5986
rect 335604 -6306 336204 -6222
rect 335604 -6542 335786 -6306
rect 336022 -6542 336204 -6306
rect 335604 -7504 336204 -6542
rect 353604 -6926 354204 30698
rect 360804 110454 361404 119800
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 364404 114054 365004 119800
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2226 365004 5498
rect 364404 -2462 364586 -2226
rect 364822 -2462 365004 -2226
rect 364404 -2546 365004 -2462
rect 364404 -2782 364586 -2546
rect 364822 -2782 365004 -2546
rect 364404 -3744 365004 -2782
rect 368004 117654 368604 119800
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4106 368604 9098
rect 368004 -4342 368186 -4106
rect 368422 -4342 368604 -4106
rect 368004 -4426 368604 -4342
rect 368004 -4662 368186 -4426
rect 368422 -4662 368604 -4426
rect 368004 -5624 368604 -4662
rect 371604 85254 372204 119800
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7162 353786 -6926
rect 354022 -7162 354204 -6926
rect 353604 -7246 354204 -7162
rect 353604 -7482 353786 -7246
rect 354022 -7482 354204 -7246
rect 353604 -7504 354204 -7482
rect 371604 -5986 372204 12698
rect 378804 92454 379404 119800
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 382404 96054 383004 119800
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 386004 99654 386604 119800
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 383331 28932 383397 28933
rect 383331 28868 383332 28932
rect 383396 28868 383397 28932
rect 383331 28867 383397 28868
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3166 383004 23498
rect 383334 21997 383394 28867
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 383331 21996 383397 21997
rect 383331 21932 383332 21996
rect 383396 21932 383397 21996
rect 383331 21931 383397 21932
rect 382404 -3402 382586 -3166
rect 382822 -3402 383004 -3166
rect 382404 -3486 383004 -3402
rect 382404 -3722 382586 -3486
rect 382822 -3722 383004 -3486
rect 382404 -3744 383004 -3722
rect 386004 -5046 386604 27098
rect 386004 -5282 386186 -5046
rect 386422 -5282 386604 -5046
rect 386004 -5366 386604 -5282
rect 386004 -5602 386186 -5366
rect 386422 -5602 386604 -5366
rect 386004 -5624 386604 -5602
rect 389604 103254 390204 119800
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6222 371786 -5986
rect 372022 -6222 372204 -5986
rect 371604 -6306 372204 -6222
rect 371604 -6542 371786 -6306
rect 372022 -6542 372204 -6306
rect 371604 -7504 372204 -6542
rect 389604 -6926 390204 30698
rect 396804 110454 397404 119800
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 400404 114054 401004 119800
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2226 401004 5498
rect 400404 -2462 400586 -2226
rect 400822 -2462 401004 -2226
rect 400404 -2546 401004 -2462
rect 400404 -2782 400586 -2546
rect 400822 -2782 401004 -2546
rect 400404 -3744 401004 -2782
rect 404004 117654 404604 119800
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4106 404604 9098
rect 404004 -4342 404186 -4106
rect 404422 -4342 404604 -4106
rect 404004 -4426 404604 -4342
rect 404004 -4662 404186 -4426
rect 404422 -4662 404604 -4426
rect 404004 -5624 404604 -4662
rect 407604 85254 408204 119800
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7162 389786 -6926
rect 390022 -7162 390204 -6926
rect 389604 -7246 390204 -7162
rect 389604 -7482 389786 -7246
rect 390022 -7482 390204 -7246
rect 389604 -7504 390204 -7482
rect 407604 -5986 408204 12698
rect 414804 92454 415404 119800
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 418404 96054 419004 119800
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3166 419004 23498
rect 418404 -3402 418586 -3166
rect 418822 -3402 419004 -3166
rect 418404 -3486 419004 -3402
rect 418404 -3722 418586 -3486
rect 418822 -3722 419004 -3486
rect 418404 -3744 419004 -3722
rect 422004 99654 422604 119800
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -5046 422604 27098
rect 422004 -5282 422186 -5046
rect 422422 -5282 422604 -5046
rect 422004 -5366 422604 -5282
rect 422004 -5602 422186 -5366
rect 422422 -5602 422604 -5366
rect 422004 -5624 422604 -5602
rect 425604 103254 426204 119800
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6222 407786 -5986
rect 408022 -6222 408204 -5986
rect 407604 -6306 408204 -6222
rect 407604 -6542 407786 -6306
rect 408022 -6542 408204 -6306
rect 407604 -7504 408204 -6542
rect 425604 -6926 426204 30698
rect 432804 110454 433404 119800
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2226 437004 5498
rect 436404 -2462 436586 -2226
rect 436822 -2462 437004 -2226
rect 436404 -2546 437004 -2462
rect 436404 -2782 436586 -2546
rect 436822 -2782 437004 -2546
rect 436404 -3744 437004 -2782
rect 440004 693654 440604 708042
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4106 440604 9098
rect 440004 -4342 440186 -4106
rect 440422 -4342 440604 -4106
rect 440004 -4426 440604 -4342
rect 440004 -4662 440186 -4426
rect 440422 -4662 440604 -4426
rect 440004 -5624 440604 -4662
rect 443604 697254 444204 709922
rect 461604 711418 462204 711440
rect 461604 711182 461786 711418
rect 462022 711182 462204 711418
rect 461604 711098 462204 711182
rect 461604 710862 461786 711098
rect 462022 710862 462204 711098
rect 458004 709538 458604 709560
rect 458004 709302 458186 709538
rect 458422 709302 458604 709538
rect 458004 709218 458604 709302
rect 458004 708982 458186 709218
rect 458422 708982 458604 709218
rect 454404 707658 455004 707680
rect 454404 707422 454586 707658
rect 454822 707422 455004 707658
rect 454404 707338 455004 707422
rect 454404 707102 454586 707338
rect 454822 707102 455004 707338
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7162 425786 -6926
rect 426022 -7162 426204 -6926
rect 425604 -7246 426204 -7162
rect 425604 -7482 425786 -7246
rect 426022 -7482 426204 -7246
rect 425604 -7504 426204 -7482
rect 443604 -5986 444204 12698
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 454404 672054 455004 707102
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3166 455004 23498
rect 454404 -3402 454586 -3166
rect 454822 -3402 455004 -3166
rect 454404 -3486 455004 -3402
rect 454404 -3722 454586 -3486
rect 454822 -3722 455004 -3486
rect 454404 -3744 455004 -3722
rect 458004 675654 458604 708982
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 461604 679254 462204 710862
rect 479604 710478 480204 711440
rect 479604 710242 479786 710478
rect 480022 710242 480204 710478
rect 479604 710158 480204 710242
rect 479604 709922 479786 710158
rect 480022 709922 480204 710158
rect 476004 708598 476604 709560
rect 476004 708362 476186 708598
rect 476422 708362 476604 708598
rect 476004 708278 476604 708362
rect 476004 708042 476186 708278
rect 476422 708042 476604 708278
rect 472404 706718 473004 707680
rect 472404 706482 472586 706718
rect 472822 706482 473004 706718
rect 472404 706398 473004 706482
rect 472404 706162 472586 706398
rect 472822 706162 473004 706398
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 387749 462204 390698
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 387749 469404 397898
rect 472404 690054 473004 706162
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 387749 473004 401498
rect 476004 693654 476604 708042
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 479604 697254 480204 709922
rect 497604 711418 498204 711440
rect 497604 711182 497786 711418
rect 498022 711182 498204 711418
rect 497604 711098 498204 711182
rect 497604 710862 497786 711098
rect 498022 710862 498204 711098
rect 494004 709538 494604 709560
rect 494004 709302 494186 709538
rect 494422 709302 494604 709538
rect 494004 709218 494604 709302
rect 494004 708982 494186 709218
rect 494422 708982 494604 709218
rect 490404 707658 491004 707680
rect 490404 707422 490586 707658
rect 490822 707422 491004 707658
rect 490404 707338 491004 707422
rect 490404 707102 490586 707338
rect 490822 707102 491004 707338
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 554964 480204 588698
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 554964 487404 559898
rect 490404 672054 491004 707102
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 554964 491004 563498
rect 494004 675654 494604 708982
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 554964 494604 567098
rect 497604 679254 498204 710862
rect 515604 710478 516204 711440
rect 515604 710242 515786 710478
rect 516022 710242 516204 710478
rect 515604 710158 516204 710242
rect 515604 709922 515786 710158
rect 516022 709922 516204 710158
rect 512004 708598 512604 709560
rect 512004 708362 512186 708598
rect 512422 708362 512604 708598
rect 512004 708278 512604 708362
rect 512004 708042 512186 708278
rect 512422 708042 512604 708278
rect 508404 706718 509004 707680
rect 508404 706482 508586 706718
rect 508822 706482 509004 706718
rect 508404 706398 509004 706482
rect 508404 706162 508586 706398
rect 508822 706162 509004 706398
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 554964 498204 570698
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 554964 505404 577898
rect 508404 690054 509004 706162
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 554964 509004 581498
rect 512004 693654 512604 708042
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 485438 542454 485758 542476
rect 485438 542218 485480 542454
rect 485716 542218 485758 542454
rect 485438 542134 485758 542218
rect 485438 541898 485480 542134
rect 485716 541898 485758 542134
rect 485438 541876 485758 541898
rect 490498 524454 490818 524476
rect 490498 524218 490540 524454
rect 490776 524218 490818 524454
rect 490498 524134 490818 524218
rect 490498 523898 490540 524134
rect 490776 523898 490818 524134
rect 490498 523876 490818 523898
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 387749 476604 405098
rect 479604 517254 480204 519800
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 387749 480204 408698
rect 486804 488454 487404 519800
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 387749 487404 415898
rect 490404 492054 491004 519800
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 387749 491004 419498
rect 494004 495654 494604 519800
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387749 494604 423098
rect 497604 499254 498204 519800
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 387749 498204 390698
rect 504804 506454 505404 519800
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 387749 505404 397898
rect 508404 510054 509004 519800
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 479568 380454 479888 380476
rect 479568 380218 479610 380454
rect 479846 380218 479888 380454
rect 479568 380134 479888 380218
rect 479568 379898 479610 380134
rect 479846 379898 479888 380134
rect 479568 379876 479888 379898
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 464208 362454 464528 362476
rect 464208 362218 464250 362454
rect 464486 362218 464528 362454
rect 464208 362134 464528 362218
rect 464208 361898 464250 362134
rect 464486 361898 464528 362134
rect 464208 361876 464528 361898
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 479568 344454 479888 344476
rect 479568 344218 479610 344454
rect 479846 344218 479888 344454
rect 479568 344134 479888 344218
rect 479568 343898 479610 344134
rect 479846 343898 479888 344134
rect 479568 343876 479888 343898
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -5046 458604 27098
rect 458004 -5282 458186 -5046
rect 458422 -5282 458604 -5046
rect 458004 -5366 458604 -5282
rect 458004 -5602 458186 -5366
rect 458422 -5602 458604 -5366
rect 458004 -5624 458604 -5602
rect 461604 319254 462204 339800
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6222 443786 -5986
rect 444022 -6222 444204 -5986
rect 443604 -6306 444204 -6222
rect 443604 -6542 443786 -6306
rect 444022 -6542 444204 -6306
rect 443604 -7504 444204 -6542
rect 461604 -6926 462204 30698
rect 468804 326454 469404 339800
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 472404 330054 473004 339800
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2226 473004 5498
rect 472404 -2462 472586 -2226
rect 472822 -2462 473004 -2226
rect 472404 -2546 473004 -2462
rect 472404 -2782 472586 -2546
rect 472822 -2782 473004 -2546
rect 472404 -3744 473004 -2782
rect 476004 333654 476604 339800
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4106 476604 9098
rect 476004 -4342 476186 -4106
rect 476422 -4342 476604 -4106
rect 476004 -4426 476604 -4342
rect 476004 -4662 476186 -4426
rect 476422 -4662 476604 -4426
rect 476004 -5624 476604 -4662
rect 479604 337254 480204 339800
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7162 461786 -6926
rect 462022 -7162 462204 -6926
rect 461604 -7246 462204 -7162
rect 461604 -7482 461786 -7246
rect 462022 -7482 462204 -7246
rect 461604 -7504 462204 -7482
rect 479604 -5986 480204 12698
rect 486804 308454 487404 339800
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 490404 312054 491004 339800
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3166 491004 23498
rect 490404 -3402 490586 -3166
rect 490822 -3402 491004 -3166
rect 490404 -3486 491004 -3402
rect 490404 -3722 490586 -3486
rect 490822 -3722 491004 -3486
rect 490404 -3744 491004 -3722
rect 494004 315654 494604 339800
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -5046 494604 27098
rect 494004 -5282 494186 -5046
rect 494422 -5282 494604 -5046
rect 494004 -5366 494604 -5282
rect 494004 -5602 494186 -5366
rect 494422 -5602 494604 -5366
rect 494004 -5624 494604 -5602
rect 497604 319254 498204 339800
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6222 479786 -5986
rect 480022 -6222 480204 -5986
rect 479604 -6306 480204 -6222
rect 479604 -6542 479786 -6306
rect 480022 -6542 480204 -6306
rect 479604 -7504 480204 -6542
rect 497604 -6926 498204 30698
rect 504804 326454 505404 339800
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2226 509004 5498
rect 508404 -2462 508586 -2226
rect 508822 -2462 509004 -2226
rect 508404 -2546 509004 -2462
rect 508404 -2782 508586 -2546
rect 508822 -2782 509004 -2546
rect 508404 -3744 509004 -2782
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4106 512604 9098
rect 512004 -4342 512186 -4106
rect 512422 -4342 512604 -4106
rect 512004 -4426 512604 -4342
rect 512004 -4662 512186 -4426
rect 512422 -4662 512604 -4426
rect 512004 -5624 512604 -4662
rect 515604 697254 516204 709922
rect 533604 711418 534204 711440
rect 533604 711182 533786 711418
rect 534022 711182 534204 711418
rect 533604 711098 534204 711182
rect 533604 710862 533786 711098
rect 534022 710862 534204 711098
rect 530004 709538 530604 709560
rect 530004 709302 530186 709538
rect 530422 709302 530604 709538
rect 530004 709218 530604 709302
rect 530004 708982 530186 709218
rect 530422 708982 530604 709218
rect 526404 707658 527004 707680
rect 526404 707422 526586 707658
rect 526822 707422 527004 707658
rect 526404 707338 527004 707422
rect 526404 707102 526586 707338
rect 526822 707102 527004 707338
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7162 497786 -6926
rect 498022 -7162 498204 -6926
rect 497604 -7246 498204 -7162
rect 497604 -7482 497786 -7246
rect 498022 -7482 498204 -7246
rect 497604 -7504 498204 -7482
rect 515604 -5986 516204 12698
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 526404 672054 527004 707102
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3166 527004 23498
rect 526404 -3402 526586 -3166
rect 526822 -3402 527004 -3166
rect 526404 -3486 527004 -3402
rect 526404 -3722 526586 -3486
rect 526822 -3722 527004 -3486
rect 526404 -3744 527004 -3722
rect 530004 675654 530604 708982
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -5046 530604 27098
rect 530004 -5282 530186 -5046
rect 530422 -5282 530604 -5046
rect 530004 -5366 530604 -5282
rect 530004 -5602 530186 -5366
rect 530422 -5602 530604 -5366
rect 530004 -5624 530604 -5602
rect 533604 679254 534204 710862
rect 551604 710478 552204 711440
rect 551604 710242 551786 710478
rect 552022 710242 552204 710478
rect 551604 710158 552204 710242
rect 551604 709922 551786 710158
rect 552022 709922 552204 710158
rect 548004 708598 548604 709560
rect 548004 708362 548186 708598
rect 548422 708362 548604 708598
rect 548004 708278 548604 708362
rect 548004 708042 548186 708278
rect 548422 708042 548604 708278
rect 544404 706718 545004 707680
rect 544404 706482 544586 706718
rect 544822 706482 545004 706718
rect 544404 706398 545004 706482
rect 544404 706162 544586 706398
rect 544822 706162 545004 706398
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6222 515786 -5986
rect 516022 -6222 516204 -5986
rect 515604 -6306 516204 -6222
rect 515604 -6542 515786 -6306
rect 516022 -6542 516204 -6306
rect 515604 -7504 516204 -6542
rect 533604 -6926 534204 30698
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 544404 690054 545004 706162
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2226 545004 5498
rect 544404 -2462 544586 -2226
rect 544822 -2462 545004 -2226
rect 544404 -2546 545004 -2462
rect 544404 -2782 544586 -2546
rect 544822 -2782 545004 -2546
rect 544404 -3744 545004 -2782
rect 548004 693654 548604 708042
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4106 548604 9098
rect 548004 -4342 548186 -4106
rect 548422 -4342 548604 -4106
rect 548004 -4426 548604 -4342
rect 548004 -4662 548186 -4426
rect 548422 -4662 548604 -4426
rect 548004 -5624 548604 -4662
rect 551604 697254 552204 709922
rect 569604 711418 570204 711440
rect 569604 711182 569786 711418
rect 570022 711182 570204 711418
rect 569604 711098 570204 711182
rect 569604 710862 569786 711098
rect 570022 710862 570204 711098
rect 566004 709538 566604 709560
rect 566004 709302 566186 709538
rect 566422 709302 566604 709538
rect 566004 709218 566604 709302
rect 566004 708982 566186 709218
rect 566422 708982 566604 709218
rect 562404 707658 563004 707680
rect 562404 707422 562586 707658
rect 562822 707422 563004 707658
rect 562404 707338 563004 707422
rect 562404 707102 562586 707338
rect 562822 707102 563004 707338
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7162 533786 -6926
rect 534022 -7162 534204 -6926
rect 533604 -7246 534204 -7162
rect 533604 -7482 533786 -7246
rect 534022 -7482 534204 -7246
rect 533604 -7504 534204 -7482
rect 551604 -5986 552204 12698
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 562404 672054 563004 707102
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3166 563004 23498
rect 562404 -3402 562586 -3166
rect 562822 -3402 563004 -3166
rect 562404 -3486 563004 -3402
rect 562404 -3722 562586 -3486
rect 562822 -3722 563004 -3486
rect 562404 -3744 563004 -3722
rect 566004 675654 566604 708982
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -5046 566604 27098
rect 566004 -5282 566186 -5046
rect 566422 -5282 566604 -5046
rect 566004 -5366 566604 -5282
rect 566004 -5602 566186 -5366
rect 566422 -5602 566604 -5366
rect 566004 -5624 566604 -5602
rect 569604 679254 570204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 580404 706718 581004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 580404 706482 580586 706718
rect 580822 706482 581004 706718
rect 580404 706398 581004 706482
rect 580404 706162 580586 706398
rect 580822 706162 581004 706398
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6222 551786 -5986
rect 552022 -6222 552204 -5986
rect 551604 -6306 552204 -6222
rect 551604 -6542 551786 -6306
rect 552022 -6542 552204 -6306
rect 551604 -7504 552204 -6542
rect 569604 -6926 570204 30698
rect 576804 704838 577404 705800
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 580404 690054 581004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2226 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 690054 587800 706162
rect 587200 689818 587382 690054
rect 587618 689818 587800 690054
rect 587200 689734 587800 689818
rect 587200 689498 587382 689734
rect 587618 689498 587800 689734
rect 587200 654054 587800 689498
rect 587200 653818 587382 654054
rect 587618 653818 587800 654054
rect 587200 653734 587800 653818
rect 587200 653498 587382 653734
rect 587618 653498 587800 653734
rect 587200 618054 587800 653498
rect 587200 617818 587382 618054
rect 587618 617818 587800 618054
rect 587200 617734 587800 617818
rect 587200 617498 587382 617734
rect 587618 617498 587800 617734
rect 587200 582054 587800 617498
rect 587200 581818 587382 582054
rect 587618 581818 587800 582054
rect 587200 581734 587800 581818
rect 587200 581498 587382 581734
rect 587618 581498 587800 581734
rect 587200 546054 587800 581498
rect 587200 545818 587382 546054
rect 587618 545818 587800 546054
rect 587200 545734 587800 545818
rect 587200 545498 587382 545734
rect 587618 545498 587800 545734
rect 587200 510054 587800 545498
rect 587200 509818 587382 510054
rect 587618 509818 587800 510054
rect 587200 509734 587800 509818
rect 587200 509498 587382 509734
rect 587618 509498 587800 509734
rect 587200 474054 587800 509498
rect 587200 473818 587382 474054
rect 587618 473818 587800 474054
rect 587200 473734 587800 473818
rect 587200 473498 587382 473734
rect 587618 473498 587800 473734
rect 587200 438054 587800 473498
rect 587200 437818 587382 438054
rect 587618 437818 587800 438054
rect 587200 437734 587800 437818
rect 587200 437498 587382 437734
rect 587618 437498 587800 437734
rect 587200 402054 587800 437498
rect 587200 401818 587382 402054
rect 587618 401818 587800 402054
rect 587200 401734 587800 401818
rect 587200 401498 587382 401734
rect 587618 401498 587800 401734
rect 587200 366054 587800 401498
rect 587200 365818 587382 366054
rect 587618 365818 587800 366054
rect 587200 365734 587800 365818
rect 587200 365498 587382 365734
rect 587618 365498 587800 365734
rect 587200 330054 587800 365498
rect 587200 329818 587382 330054
rect 587618 329818 587800 330054
rect 587200 329734 587800 329818
rect 587200 329498 587382 329734
rect 587618 329498 587800 329734
rect 587200 294054 587800 329498
rect 587200 293818 587382 294054
rect 587618 293818 587800 294054
rect 587200 293734 587800 293818
rect 587200 293498 587382 293734
rect 587618 293498 587800 293734
rect 587200 258054 587800 293498
rect 587200 257818 587382 258054
rect 587618 257818 587800 258054
rect 587200 257734 587800 257818
rect 587200 257498 587382 257734
rect 587618 257498 587800 257734
rect 587200 222054 587800 257498
rect 587200 221818 587382 222054
rect 587618 221818 587800 222054
rect 587200 221734 587800 221818
rect 587200 221498 587382 221734
rect 587618 221498 587800 221734
rect 587200 186054 587800 221498
rect 587200 185818 587382 186054
rect 587618 185818 587800 186054
rect 587200 185734 587800 185818
rect 587200 185498 587382 185734
rect 587618 185498 587800 185734
rect 587200 150054 587800 185498
rect 587200 149818 587382 150054
rect 587618 149818 587800 150054
rect 587200 149734 587800 149818
rect 587200 149498 587382 149734
rect 587618 149498 587800 149734
rect 587200 114054 587800 149498
rect 587200 113818 587382 114054
rect 587618 113818 587800 114054
rect 587200 113734 587800 113818
rect 587200 113498 587382 113734
rect 587618 113498 587800 113734
rect 587200 78054 587800 113498
rect 587200 77818 587382 78054
rect 587618 77818 587800 78054
rect 587200 77734 587800 77818
rect 587200 77498 587382 77734
rect 587618 77498 587800 77734
rect 587200 42054 587800 77498
rect 587200 41818 587382 42054
rect 587618 41818 587800 42054
rect 587200 41734 587800 41818
rect 587200 41498 587382 41734
rect 587618 41498 587800 41734
rect 587200 6054 587800 41498
rect 587200 5818 587382 6054
rect 587618 5818 587800 6054
rect 587200 5734 587800 5818
rect 587200 5498 587382 5734
rect 587618 5498 587800 5734
rect 580404 -2462 580586 -2226
rect 580822 -2462 581004 -2226
rect 580404 -2546 581004 -2462
rect 580404 -2782 580586 -2546
rect 580822 -2782 581004 -2546
rect 580404 -3744 581004 -2782
rect 587200 -2226 587800 5498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 672054 588740 707102
rect 588140 671818 588322 672054
rect 588558 671818 588740 672054
rect 588140 671734 588740 671818
rect 588140 671498 588322 671734
rect 588558 671498 588740 671734
rect 588140 636054 588740 671498
rect 588140 635818 588322 636054
rect 588558 635818 588740 636054
rect 588140 635734 588740 635818
rect 588140 635498 588322 635734
rect 588558 635498 588740 635734
rect 588140 600054 588740 635498
rect 588140 599818 588322 600054
rect 588558 599818 588740 600054
rect 588140 599734 588740 599818
rect 588140 599498 588322 599734
rect 588558 599498 588740 599734
rect 588140 564054 588740 599498
rect 588140 563818 588322 564054
rect 588558 563818 588740 564054
rect 588140 563734 588740 563818
rect 588140 563498 588322 563734
rect 588558 563498 588740 563734
rect 588140 528054 588740 563498
rect 588140 527818 588322 528054
rect 588558 527818 588740 528054
rect 588140 527734 588740 527818
rect 588140 527498 588322 527734
rect 588558 527498 588740 527734
rect 588140 492054 588740 527498
rect 588140 491818 588322 492054
rect 588558 491818 588740 492054
rect 588140 491734 588740 491818
rect 588140 491498 588322 491734
rect 588558 491498 588740 491734
rect 588140 456054 588740 491498
rect 588140 455818 588322 456054
rect 588558 455818 588740 456054
rect 588140 455734 588740 455818
rect 588140 455498 588322 455734
rect 588558 455498 588740 455734
rect 588140 420054 588740 455498
rect 588140 419818 588322 420054
rect 588558 419818 588740 420054
rect 588140 419734 588740 419818
rect 588140 419498 588322 419734
rect 588558 419498 588740 419734
rect 588140 384054 588740 419498
rect 588140 383818 588322 384054
rect 588558 383818 588740 384054
rect 588140 383734 588740 383818
rect 588140 383498 588322 383734
rect 588558 383498 588740 383734
rect 588140 348054 588740 383498
rect 588140 347818 588322 348054
rect 588558 347818 588740 348054
rect 588140 347734 588740 347818
rect 588140 347498 588322 347734
rect 588558 347498 588740 347734
rect 588140 312054 588740 347498
rect 588140 311818 588322 312054
rect 588558 311818 588740 312054
rect 588140 311734 588740 311818
rect 588140 311498 588322 311734
rect 588558 311498 588740 311734
rect 588140 276054 588740 311498
rect 588140 275818 588322 276054
rect 588558 275818 588740 276054
rect 588140 275734 588740 275818
rect 588140 275498 588322 275734
rect 588558 275498 588740 275734
rect 588140 240054 588740 275498
rect 588140 239818 588322 240054
rect 588558 239818 588740 240054
rect 588140 239734 588740 239818
rect 588140 239498 588322 239734
rect 588558 239498 588740 239734
rect 588140 204054 588740 239498
rect 588140 203818 588322 204054
rect 588558 203818 588740 204054
rect 588140 203734 588740 203818
rect 588140 203498 588322 203734
rect 588558 203498 588740 203734
rect 588140 168054 588740 203498
rect 588140 167818 588322 168054
rect 588558 167818 588740 168054
rect 588140 167734 588740 167818
rect 588140 167498 588322 167734
rect 588558 167498 588740 167734
rect 588140 132054 588740 167498
rect 588140 131818 588322 132054
rect 588558 131818 588740 132054
rect 588140 131734 588740 131818
rect 588140 131498 588322 131734
rect 588558 131498 588740 131734
rect 588140 96054 588740 131498
rect 588140 95818 588322 96054
rect 588558 95818 588740 96054
rect 588140 95734 588740 95818
rect 588140 95498 588322 95734
rect 588558 95498 588740 95734
rect 588140 60054 588740 95498
rect 588140 59818 588322 60054
rect 588558 59818 588740 60054
rect 588140 59734 588740 59818
rect 588140 59498 588322 59734
rect 588558 59498 588740 59734
rect 588140 24054 588740 59498
rect 588140 23818 588322 24054
rect 588558 23818 588740 24054
rect 588140 23734 588740 23818
rect 588140 23498 588322 23734
rect 588558 23498 588740 23734
rect 588140 -3166 588740 23498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 693654 589680 708042
rect 589080 693418 589262 693654
rect 589498 693418 589680 693654
rect 589080 693334 589680 693418
rect 589080 693098 589262 693334
rect 589498 693098 589680 693334
rect 589080 657654 589680 693098
rect 589080 657418 589262 657654
rect 589498 657418 589680 657654
rect 589080 657334 589680 657418
rect 589080 657098 589262 657334
rect 589498 657098 589680 657334
rect 589080 621654 589680 657098
rect 589080 621418 589262 621654
rect 589498 621418 589680 621654
rect 589080 621334 589680 621418
rect 589080 621098 589262 621334
rect 589498 621098 589680 621334
rect 589080 585654 589680 621098
rect 589080 585418 589262 585654
rect 589498 585418 589680 585654
rect 589080 585334 589680 585418
rect 589080 585098 589262 585334
rect 589498 585098 589680 585334
rect 589080 549654 589680 585098
rect 589080 549418 589262 549654
rect 589498 549418 589680 549654
rect 589080 549334 589680 549418
rect 589080 549098 589262 549334
rect 589498 549098 589680 549334
rect 589080 513654 589680 549098
rect 589080 513418 589262 513654
rect 589498 513418 589680 513654
rect 589080 513334 589680 513418
rect 589080 513098 589262 513334
rect 589498 513098 589680 513334
rect 589080 477654 589680 513098
rect 589080 477418 589262 477654
rect 589498 477418 589680 477654
rect 589080 477334 589680 477418
rect 589080 477098 589262 477334
rect 589498 477098 589680 477334
rect 589080 441654 589680 477098
rect 589080 441418 589262 441654
rect 589498 441418 589680 441654
rect 589080 441334 589680 441418
rect 589080 441098 589262 441334
rect 589498 441098 589680 441334
rect 589080 405654 589680 441098
rect 589080 405418 589262 405654
rect 589498 405418 589680 405654
rect 589080 405334 589680 405418
rect 589080 405098 589262 405334
rect 589498 405098 589680 405334
rect 589080 369654 589680 405098
rect 589080 369418 589262 369654
rect 589498 369418 589680 369654
rect 589080 369334 589680 369418
rect 589080 369098 589262 369334
rect 589498 369098 589680 369334
rect 589080 333654 589680 369098
rect 589080 333418 589262 333654
rect 589498 333418 589680 333654
rect 589080 333334 589680 333418
rect 589080 333098 589262 333334
rect 589498 333098 589680 333334
rect 589080 297654 589680 333098
rect 589080 297418 589262 297654
rect 589498 297418 589680 297654
rect 589080 297334 589680 297418
rect 589080 297098 589262 297334
rect 589498 297098 589680 297334
rect 589080 261654 589680 297098
rect 589080 261418 589262 261654
rect 589498 261418 589680 261654
rect 589080 261334 589680 261418
rect 589080 261098 589262 261334
rect 589498 261098 589680 261334
rect 589080 225654 589680 261098
rect 589080 225418 589262 225654
rect 589498 225418 589680 225654
rect 589080 225334 589680 225418
rect 589080 225098 589262 225334
rect 589498 225098 589680 225334
rect 589080 189654 589680 225098
rect 589080 189418 589262 189654
rect 589498 189418 589680 189654
rect 589080 189334 589680 189418
rect 589080 189098 589262 189334
rect 589498 189098 589680 189334
rect 589080 153654 589680 189098
rect 589080 153418 589262 153654
rect 589498 153418 589680 153654
rect 589080 153334 589680 153418
rect 589080 153098 589262 153334
rect 589498 153098 589680 153334
rect 589080 117654 589680 153098
rect 589080 117418 589262 117654
rect 589498 117418 589680 117654
rect 589080 117334 589680 117418
rect 589080 117098 589262 117334
rect 589498 117098 589680 117334
rect 589080 81654 589680 117098
rect 589080 81418 589262 81654
rect 589498 81418 589680 81654
rect 589080 81334 589680 81418
rect 589080 81098 589262 81334
rect 589498 81098 589680 81334
rect 589080 45654 589680 81098
rect 589080 45418 589262 45654
rect 589498 45418 589680 45654
rect 589080 45334 589680 45418
rect 589080 45098 589262 45334
rect 589498 45098 589680 45334
rect 589080 9654 589680 45098
rect 589080 9418 589262 9654
rect 589498 9418 589680 9654
rect 589080 9334 589680 9418
rect 589080 9098 589262 9334
rect 589498 9098 589680 9334
rect 589080 -4106 589680 9098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 675654 590620 708982
rect 590020 675418 590202 675654
rect 590438 675418 590620 675654
rect 590020 675334 590620 675418
rect 590020 675098 590202 675334
rect 590438 675098 590620 675334
rect 590020 639654 590620 675098
rect 590020 639418 590202 639654
rect 590438 639418 590620 639654
rect 590020 639334 590620 639418
rect 590020 639098 590202 639334
rect 590438 639098 590620 639334
rect 590020 603654 590620 639098
rect 590020 603418 590202 603654
rect 590438 603418 590620 603654
rect 590020 603334 590620 603418
rect 590020 603098 590202 603334
rect 590438 603098 590620 603334
rect 590020 567654 590620 603098
rect 590020 567418 590202 567654
rect 590438 567418 590620 567654
rect 590020 567334 590620 567418
rect 590020 567098 590202 567334
rect 590438 567098 590620 567334
rect 590020 531654 590620 567098
rect 590020 531418 590202 531654
rect 590438 531418 590620 531654
rect 590020 531334 590620 531418
rect 590020 531098 590202 531334
rect 590438 531098 590620 531334
rect 590020 495654 590620 531098
rect 590020 495418 590202 495654
rect 590438 495418 590620 495654
rect 590020 495334 590620 495418
rect 590020 495098 590202 495334
rect 590438 495098 590620 495334
rect 590020 459654 590620 495098
rect 590020 459418 590202 459654
rect 590438 459418 590620 459654
rect 590020 459334 590620 459418
rect 590020 459098 590202 459334
rect 590438 459098 590620 459334
rect 590020 423654 590620 459098
rect 590020 423418 590202 423654
rect 590438 423418 590620 423654
rect 590020 423334 590620 423418
rect 590020 423098 590202 423334
rect 590438 423098 590620 423334
rect 590020 387654 590620 423098
rect 590020 387418 590202 387654
rect 590438 387418 590620 387654
rect 590020 387334 590620 387418
rect 590020 387098 590202 387334
rect 590438 387098 590620 387334
rect 590020 351654 590620 387098
rect 590020 351418 590202 351654
rect 590438 351418 590620 351654
rect 590020 351334 590620 351418
rect 590020 351098 590202 351334
rect 590438 351098 590620 351334
rect 590020 315654 590620 351098
rect 590020 315418 590202 315654
rect 590438 315418 590620 315654
rect 590020 315334 590620 315418
rect 590020 315098 590202 315334
rect 590438 315098 590620 315334
rect 590020 279654 590620 315098
rect 590020 279418 590202 279654
rect 590438 279418 590620 279654
rect 590020 279334 590620 279418
rect 590020 279098 590202 279334
rect 590438 279098 590620 279334
rect 590020 243654 590620 279098
rect 590020 243418 590202 243654
rect 590438 243418 590620 243654
rect 590020 243334 590620 243418
rect 590020 243098 590202 243334
rect 590438 243098 590620 243334
rect 590020 207654 590620 243098
rect 590020 207418 590202 207654
rect 590438 207418 590620 207654
rect 590020 207334 590620 207418
rect 590020 207098 590202 207334
rect 590438 207098 590620 207334
rect 590020 171654 590620 207098
rect 590020 171418 590202 171654
rect 590438 171418 590620 171654
rect 590020 171334 590620 171418
rect 590020 171098 590202 171334
rect 590438 171098 590620 171334
rect 590020 135654 590620 171098
rect 590020 135418 590202 135654
rect 590438 135418 590620 135654
rect 590020 135334 590620 135418
rect 590020 135098 590202 135334
rect 590438 135098 590620 135334
rect 590020 99654 590620 135098
rect 590020 99418 590202 99654
rect 590438 99418 590620 99654
rect 590020 99334 590620 99418
rect 590020 99098 590202 99334
rect 590438 99098 590620 99334
rect 590020 63654 590620 99098
rect 590020 63418 590202 63654
rect 590438 63418 590620 63654
rect 590020 63334 590620 63418
rect 590020 63098 590202 63334
rect 590438 63098 590620 63334
rect 590020 27654 590620 63098
rect 590020 27418 590202 27654
rect 590438 27418 590620 27654
rect 590020 27334 590620 27418
rect 590020 27098 590202 27334
rect 590438 27098 590620 27334
rect 590020 -5046 590620 27098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 697254 591560 709922
rect 590960 697018 591142 697254
rect 591378 697018 591560 697254
rect 590960 696934 591560 697018
rect 590960 696698 591142 696934
rect 591378 696698 591560 696934
rect 590960 661254 591560 696698
rect 590960 661018 591142 661254
rect 591378 661018 591560 661254
rect 590960 660934 591560 661018
rect 590960 660698 591142 660934
rect 591378 660698 591560 660934
rect 590960 625254 591560 660698
rect 590960 625018 591142 625254
rect 591378 625018 591560 625254
rect 590960 624934 591560 625018
rect 590960 624698 591142 624934
rect 591378 624698 591560 624934
rect 590960 589254 591560 624698
rect 590960 589018 591142 589254
rect 591378 589018 591560 589254
rect 590960 588934 591560 589018
rect 590960 588698 591142 588934
rect 591378 588698 591560 588934
rect 590960 553254 591560 588698
rect 590960 553018 591142 553254
rect 591378 553018 591560 553254
rect 590960 552934 591560 553018
rect 590960 552698 591142 552934
rect 591378 552698 591560 552934
rect 590960 517254 591560 552698
rect 590960 517018 591142 517254
rect 591378 517018 591560 517254
rect 590960 516934 591560 517018
rect 590960 516698 591142 516934
rect 591378 516698 591560 516934
rect 590960 481254 591560 516698
rect 590960 481018 591142 481254
rect 591378 481018 591560 481254
rect 590960 480934 591560 481018
rect 590960 480698 591142 480934
rect 591378 480698 591560 480934
rect 590960 445254 591560 480698
rect 590960 445018 591142 445254
rect 591378 445018 591560 445254
rect 590960 444934 591560 445018
rect 590960 444698 591142 444934
rect 591378 444698 591560 444934
rect 590960 409254 591560 444698
rect 590960 409018 591142 409254
rect 591378 409018 591560 409254
rect 590960 408934 591560 409018
rect 590960 408698 591142 408934
rect 591378 408698 591560 408934
rect 590960 373254 591560 408698
rect 590960 373018 591142 373254
rect 591378 373018 591560 373254
rect 590960 372934 591560 373018
rect 590960 372698 591142 372934
rect 591378 372698 591560 372934
rect 590960 337254 591560 372698
rect 590960 337018 591142 337254
rect 591378 337018 591560 337254
rect 590960 336934 591560 337018
rect 590960 336698 591142 336934
rect 591378 336698 591560 336934
rect 590960 301254 591560 336698
rect 590960 301018 591142 301254
rect 591378 301018 591560 301254
rect 590960 300934 591560 301018
rect 590960 300698 591142 300934
rect 591378 300698 591560 300934
rect 590960 265254 591560 300698
rect 590960 265018 591142 265254
rect 591378 265018 591560 265254
rect 590960 264934 591560 265018
rect 590960 264698 591142 264934
rect 591378 264698 591560 264934
rect 590960 229254 591560 264698
rect 590960 229018 591142 229254
rect 591378 229018 591560 229254
rect 590960 228934 591560 229018
rect 590960 228698 591142 228934
rect 591378 228698 591560 228934
rect 590960 193254 591560 228698
rect 590960 193018 591142 193254
rect 591378 193018 591560 193254
rect 590960 192934 591560 193018
rect 590960 192698 591142 192934
rect 591378 192698 591560 192934
rect 590960 157254 591560 192698
rect 590960 157018 591142 157254
rect 591378 157018 591560 157254
rect 590960 156934 591560 157018
rect 590960 156698 591142 156934
rect 591378 156698 591560 156934
rect 590960 121254 591560 156698
rect 590960 121018 591142 121254
rect 591378 121018 591560 121254
rect 590960 120934 591560 121018
rect 590960 120698 591142 120934
rect 591378 120698 591560 120934
rect 590960 85254 591560 120698
rect 590960 85018 591142 85254
rect 591378 85018 591560 85254
rect 590960 84934 591560 85018
rect 590960 84698 591142 84934
rect 591378 84698 591560 84934
rect 590960 49254 591560 84698
rect 590960 49018 591142 49254
rect 591378 49018 591560 49254
rect 590960 48934 591560 49018
rect 590960 48698 591142 48934
rect 591378 48698 591560 48934
rect 590960 13254 591560 48698
rect 590960 13018 591142 13254
rect 591378 13018 591560 13254
rect 590960 12934 591560 13018
rect 590960 12698 591142 12934
rect 591378 12698 591560 12934
rect 590960 -5986 591560 12698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 679254 592500 710862
rect 591900 679018 592082 679254
rect 592318 679018 592500 679254
rect 591900 678934 592500 679018
rect 591900 678698 592082 678934
rect 592318 678698 592500 678934
rect 591900 643254 592500 678698
rect 591900 643018 592082 643254
rect 592318 643018 592500 643254
rect 591900 642934 592500 643018
rect 591900 642698 592082 642934
rect 592318 642698 592500 642934
rect 591900 607254 592500 642698
rect 591900 607018 592082 607254
rect 592318 607018 592500 607254
rect 591900 606934 592500 607018
rect 591900 606698 592082 606934
rect 592318 606698 592500 606934
rect 591900 571254 592500 606698
rect 591900 571018 592082 571254
rect 592318 571018 592500 571254
rect 591900 570934 592500 571018
rect 591900 570698 592082 570934
rect 592318 570698 592500 570934
rect 591900 535254 592500 570698
rect 591900 535018 592082 535254
rect 592318 535018 592500 535254
rect 591900 534934 592500 535018
rect 591900 534698 592082 534934
rect 592318 534698 592500 534934
rect 591900 499254 592500 534698
rect 591900 499018 592082 499254
rect 592318 499018 592500 499254
rect 591900 498934 592500 499018
rect 591900 498698 592082 498934
rect 592318 498698 592500 498934
rect 591900 463254 592500 498698
rect 591900 463018 592082 463254
rect 592318 463018 592500 463254
rect 591900 462934 592500 463018
rect 591900 462698 592082 462934
rect 592318 462698 592500 462934
rect 591900 427254 592500 462698
rect 591900 427018 592082 427254
rect 592318 427018 592500 427254
rect 591900 426934 592500 427018
rect 591900 426698 592082 426934
rect 592318 426698 592500 426934
rect 591900 391254 592500 426698
rect 591900 391018 592082 391254
rect 592318 391018 592500 391254
rect 591900 390934 592500 391018
rect 591900 390698 592082 390934
rect 592318 390698 592500 390934
rect 591900 355254 592500 390698
rect 591900 355018 592082 355254
rect 592318 355018 592500 355254
rect 591900 354934 592500 355018
rect 591900 354698 592082 354934
rect 592318 354698 592500 354934
rect 591900 319254 592500 354698
rect 591900 319018 592082 319254
rect 592318 319018 592500 319254
rect 591900 318934 592500 319018
rect 591900 318698 592082 318934
rect 592318 318698 592500 318934
rect 591900 283254 592500 318698
rect 591900 283018 592082 283254
rect 592318 283018 592500 283254
rect 591900 282934 592500 283018
rect 591900 282698 592082 282934
rect 592318 282698 592500 282934
rect 591900 247254 592500 282698
rect 591900 247018 592082 247254
rect 592318 247018 592500 247254
rect 591900 246934 592500 247018
rect 591900 246698 592082 246934
rect 592318 246698 592500 246934
rect 591900 211254 592500 246698
rect 591900 211018 592082 211254
rect 592318 211018 592500 211254
rect 591900 210934 592500 211018
rect 591900 210698 592082 210934
rect 592318 210698 592500 210934
rect 591900 175254 592500 210698
rect 591900 175018 592082 175254
rect 592318 175018 592500 175254
rect 591900 174934 592500 175018
rect 591900 174698 592082 174934
rect 592318 174698 592500 174934
rect 591900 139254 592500 174698
rect 591900 139018 592082 139254
rect 592318 139018 592500 139254
rect 591900 138934 592500 139018
rect 591900 138698 592082 138934
rect 592318 138698 592500 138934
rect 591900 103254 592500 138698
rect 591900 103018 592082 103254
rect 592318 103018 592500 103254
rect 591900 102934 592500 103018
rect 591900 102698 592082 102934
rect 592318 102698 592500 102934
rect 591900 67254 592500 102698
rect 591900 67018 592082 67254
rect 592318 67018 592500 67254
rect 591900 66934 592500 67018
rect 591900 66698 592082 66934
rect 592318 66698 592500 66934
rect 591900 31254 592500 66698
rect 591900 31018 592082 31254
rect 592318 31018 592500 31254
rect 591900 30934 592500 31018
rect 591900 30698 592082 30934
rect 592318 30698 592500 30934
rect 569604 -7162 569786 -6926
rect 570022 -7162 570204 -6926
rect 569604 -7246 570204 -7162
rect 569604 -7482 569786 -7246
rect 570022 -7482 570204 -7246
rect 569604 -7504 570204 -7482
rect 591900 -6926 592500 30698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 679018 -8158 679254
rect -8394 678698 -8158 678934
rect -8394 643018 -8158 643254
rect -8394 642698 -8158 642934
rect -8394 607018 -8158 607254
rect -8394 606698 -8158 606934
rect -8394 571018 -8158 571254
rect -8394 570698 -8158 570934
rect -8394 535018 -8158 535254
rect -8394 534698 -8158 534934
rect -8394 499018 -8158 499254
rect -8394 498698 -8158 498934
rect -8394 463018 -8158 463254
rect -8394 462698 -8158 462934
rect -8394 427018 -8158 427254
rect -8394 426698 -8158 426934
rect -8394 391018 -8158 391254
rect -8394 390698 -8158 390934
rect -8394 355018 -8158 355254
rect -8394 354698 -8158 354934
rect -8394 319018 -8158 319254
rect -8394 318698 -8158 318934
rect -8394 283018 -8158 283254
rect -8394 282698 -8158 282934
rect -8394 247018 -8158 247254
rect -8394 246698 -8158 246934
rect -8394 211018 -8158 211254
rect -8394 210698 -8158 210934
rect -8394 175018 -8158 175254
rect -8394 174698 -8158 174934
rect -8394 139018 -8158 139254
rect -8394 138698 -8158 138934
rect -8394 103018 -8158 103254
rect -8394 102698 -8158 102934
rect -8394 67018 -8158 67254
rect -8394 66698 -8158 66934
rect -8394 31018 -8158 31254
rect -8394 30698 -8158 30934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 11786 710242 12022 710478
rect 11786 709922 12022 710158
rect -7454 697018 -7218 697254
rect -7454 696698 -7218 696934
rect -7454 661018 -7218 661254
rect -7454 660698 -7218 660934
rect -7454 625018 -7218 625254
rect -7454 624698 -7218 624934
rect -7454 589018 -7218 589254
rect -7454 588698 -7218 588934
rect -7454 553018 -7218 553254
rect -7454 552698 -7218 552934
rect -7454 517018 -7218 517254
rect -7454 516698 -7218 516934
rect -7454 481018 -7218 481254
rect -7454 480698 -7218 480934
rect -7454 445018 -7218 445254
rect -7454 444698 -7218 444934
rect -7454 409018 -7218 409254
rect -7454 408698 -7218 408934
rect -7454 373018 -7218 373254
rect -7454 372698 -7218 372934
rect -7454 337018 -7218 337254
rect -7454 336698 -7218 336934
rect -7454 301018 -7218 301254
rect -7454 300698 -7218 300934
rect -7454 265018 -7218 265254
rect -7454 264698 -7218 264934
rect -7454 229018 -7218 229254
rect -7454 228698 -7218 228934
rect -7454 193018 -7218 193254
rect -7454 192698 -7218 192934
rect -7454 157018 -7218 157254
rect -7454 156698 -7218 156934
rect -7454 121018 -7218 121254
rect -7454 120698 -7218 120934
rect -7454 85018 -7218 85254
rect -7454 84698 -7218 84934
rect -7454 49018 -7218 49254
rect -7454 48698 -7218 48934
rect -7454 13018 -7218 13254
rect -7454 12698 -7218 12934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 675418 -6278 675654
rect -6514 675098 -6278 675334
rect -6514 639418 -6278 639654
rect -6514 639098 -6278 639334
rect -6514 603418 -6278 603654
rect -6514 603098 -6278 603334
rect -6514 567418 -6278 567654
rect -6514 567098 -6278 567334
rect -6514 531418 -6278 531654
rect -6514 531098 -6278 531334
rect -6514 495418 -6278 495654
rect -6514 495098 -6278 495334
rect -6514 459418 -6278 459654
rect -6514 459098 -6278 459334
rect -6514 423418 -6278 423654
rect -6514 423098 -6278 423334
rect -6514 387418 -6278 387654
rect -6514 387098 -6278 387334
rect -6514 351418 -6278 351654
rect -6514 351098 -6278 351334
rect -6514 315418 -6278 315654
rect -6514 315098 -6278 315334
rect -6514 279418 -6278 279654
rect -6514 279098 -6278 279334
rect -6514 243418 -6278 243654
rect -6514 243098 -6278 243334
rect -6514 207418 -6278 207654
rect -6514 207098 -6278 207334
rect -6514 171418 -6278 171654
rect -6514 171098 -6278 171334
rect -6514 135418 -6278 135654
rect -6514 135098 -6278 135334
rect -6514 99418 -6278 99654
rect -6514 99098 -6278 99334
rect -6514 63418 -6278 63654
rect -6514 63098 -6278 63334
rect -6514 27418 -6278 27654
rect -6514 27098 -6278 27334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 8186 708362 8422 708598
rect 8186 708042 8422 708278
rect -5574 693418 -5338 693654
rect -5574 693098 -5338 693334
rect -5574 657418 -5338 657654
rect -5574 657098 -5338 657334
rect -5574 621418 -5338 621654
rect -5574 621098 -5338 621334
rect -5574 585418 -5338 585654
rect -5574 585098 -5338 585334
rect -5574 549418 -5338 549654
rect -5574 549098 -5338 549334
rect -5574 513418 -5338 513654
rect -5574 513098 -5338 513334
rect -5574 477418 -5338 477654
rect -5574 477098 -5338 477334
rect -5574 441418 -5338 441654
rect -5574 441098 -5338 441334
rect -5574 405418 -5338 405654
rect -5574 405098 -5338 405334
rect -5574 369418 -5338 369654
rect -5574 369098 -5338 369334
rect -5574 333418 -5338 333654
rect -5574 333098 -5338 333334
rect -5574 297418 -5338 297654
rect -5574 297098 -5338 297334
rect -5574 261418 -5338 261654
rect -5574 261098 -5338 261334
rect -5574 225418 -5338 225654
rect -5574 225098 -5338 225334
rect -5574 189418 -5338 189654
rect -5574 189098 -5338 189334
rect -5574 153418 -5338 153654
rect -5574 153098 -5338 153334
rect -5574 117418 -5338 117654
rect -5574 117098 -5338 117334
rect -5574 81418 -5338 81654
rect -5574 81098 -5338 81334
rect -5574 45418 -5338 45654
rect -5574 45098 -5338 45334
rect -5574 9418 -5338 9654
rect -5574 9098 -5338 9334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 671818 -4398 672054
rect -4634 671498 -4398 671734
rect -4634 635818 -4398 636054
rect -4634 635498 -4398 635734
rect -4634 599818 -4398 600054
rect -4634 599498 -4398 599734
rect -4634 563818 -4398 564054
rect -4634 563498 -4398 563734
rect -4634 527818 -4398 528054
rect -4634 527498 -4398 527734
rect -4634 491818 -4398 492054
rect -4634 491498 -4398 491734
rect -4634 455818 -4398 456054
rect -4634 455498 -4398 455734
rect -4634 419818 -4398 420054
rect -4634 419498 -4398 419734
rect -4634 383818 -4398 384054
rect -4634 383498 -4398 383734
rect -4634 347818 -4398 348054
rect -4634 347498 -4398 347734
rect -4634 311818 -4398 312054
rect -4634 311498 -4398 311734
rect -4634 275818 -4398 276054
rect -4634 275498 -4398 275734
rect -4634 239818 -4398 240054
rect -4634 239498 -4398 239734
rect -4634 203818 -4398 204054
rect -4634 203498 -4398 203734
rect -4634 167818 -4398 168054
rect -4634 167498 -4398 167734
rect -4634 131818 -4398 132054
rect -4634 131498 -4398 131734
rect -4634 95818 -4398 96054
rect -4634 95498 -4398 95734
rect -4634 59818 -4398 60054
rect -4634 59498 -4398 59734
rect -4634 23818 -4398 24054
rect -4634 23498 -4398 23734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 4586 706482 4822 706718
rect 4586 706162 4822 706398
rect -3694 689818 -3458 690054
rect -3694 689498 -3458 689734
rect -3694 653818 -3458 654054
rect -3694 653498 -3458 653734
rect -3694 617818 -3458 618054
rect -3694 617498 -3458 617734
rect -3694 581818 -3458 582054
rect -3694 581498 -3458 581734
rect -3694 545818 -3458 546054
rect -3694 545498 -3458 545734
rect -3694 509818 -3458 510054
rect -3694 509498 -3458 509734
rect -3694 473818 -3458 474054
rect -3694 473498 -3458 473734
rect -3694 437818 -3458 438054
rect -3694 437498 -3458 437734
rect -3694 401818 -3458 402054
rect -3694 401498 -3458 401734
rect -3694 365818 -3458 366054
rect -3694 365498 -3458 365734
rect -3694 329818 -3458 330054
rect -3694 329498 -3458 329734
rect -3694 293818 -3458 294054
rect -3694 293498 -3458 293734
rect -3694 257818 -3458 258054
rect -3694 257498 -3458 257734
rect -3694 221818 -3458 222054
rect -3694 221498 -3458 221734
rect -3694 185818 -3458 186054
rect -3694 185498 -3458 185734
rect -3694 149818 -3458 150054
rect -3694 149498 -3458 149734
rect -3694 113818 -3458 114054
rect -3694 113498 -3458 113734
rect -3694 77818 -3458 78054
rect -3694 77498 -3458 77734
rect -3694 41818 -3458 42054
rect -3694 41498 -3458 41734
rect -3694 5818 -3458 6054
rect -3694 5498 -3458 5734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 4586 -2462 4822 -2226
rect 4586 -2782 4822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 8186 -4342 8422 -4106
rect 8186 -4662 8422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 29786 711182 30022 711418
rect 29786 710862 30022 711098
rect 26186 709302 26422 709538
rect 26186 708982 26422 709218
rect 22586 707422 22822 707658
rect 22586 707102 22822 707338
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3402 22822 -3166
rect 22586 -3722 22822 -3486
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5282 26422 -5046
rect 26186 -5602 26422 -5366
rect 47786 710242 48022 710478
rect 47786 709922 48022 710158
rect 44186 708362 44422 708598
rect 44186 708042 44422 708278
rect 40586 706482 40822 706718
rect 40586 706162 40822 706398
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6222 12022 -5986
rect 11786 -6542 12022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2462 40822 -2226
rect 40586 -2782 40822 -2546
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4342 44422 -4106
rect 44186 -4662 44422 -4426
rect 65786 711182 66022 711418
rect 65786 710862 66022 711098
rect 62186 709302 62422 709538
rect 62186 708982 62422 709218
rect 58586 707422 58822 707658
rect 58586 707102 58822 707338
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7162 30022 -6926
rect 29786 -7482 30022 -7246
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3402 58822 -3166
rect 58586 -3722 58822 -3486
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5282 62422 -5046
rect 62186 -5602 62422 -5366
rect 83786 710242 84022 710478
rect 83786 709922 84022 710158
rect 80186 708362 80422 708598
rect 80186 708042 80422 708278
rect 76586 706482 76822 706718
rect 76586 706162 76822 706398
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 101786 711182 102022 711418
rect 101786 710862 102022 711098
rect 98186 709302 98422 709538
rect 98186 708982 98422 709218
rect 94586 707422 94822 707658
rect 94586 707102 94822 707338
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 119786 710242 120022 710478
rect 119786 709922 120022 710158
rect 116186 708362 116422 708598
rect 116186 708042 116422 708278
rect 112586 706482 112822 706718
rect 112586 706162 112822 706398
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 91571 542218 91807 542454
rect 91571 541898 91807 542134
rect 96155 524218 96391 524454
rect 96155 523898 96391 524134
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 137786 711182 138022 711418
rect 137786 710862 138022 711098
rect 134186 709302 134422 709538
rect 134186 708982 134422 709218
rect 130586 707422 130822 707658
rect 130586 707102 130822 707338
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 91610 380218 91846 380454
rect 91610 379898 91846 380134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 76250 362218 76486 362454
rect 76250 361898 76486 362134
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 91610 344218 91846 344454
rect 91610 343898 91846 344134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6222 48022 -5986
rect 47786 -6542 48022 -6306
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2462 76822 -2226
rect 76586 -2782 76822 -2546
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4342 80422 -4106
rect 80186 -4662 80422 -4426
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7162 66022 -6926
rect 65786 -7482 66022 -7246
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3402 94822 -3166
rect 94586 -3722 94822 -3486
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5282 98422 -5046
rect 98186 -5602 98422 -5366
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6222 84022 -5986
rect 83786 -6542 84022 -6306
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2462 112822 -2226
rect 112586 -2782 112822 -2546
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4342 116422 -4106
rect 116186 -4662 116422 -4426
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7162 102022 -6926
rect 101786 -7482 102022 -7246
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 155786 710242 156022 710478
rect 155786 709922 156022 710158
rect 152186 708362 152422 708598
rect 152186 708042 152422 708278
rect 148586 706482 148822 706718
rect 148586 706162 148822 706398
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 173786 711182 174022 711418
rect 173786 710862 174022 711098
rect 170186 709302 170422 709538
rect 170186 708982 170422 709218
rect 166586 707422 166822 707658
rect 166586 707102 166822 707338
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 155786 409018 156022 409254
rect 155786 408698 156022 408934
rect 155786 373018 156022 373254
rect 155786 372698 156022 372934
rect 155786 337018 156022 337254
rect 155786 336698 156022 336934
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 166586 383818 166822 384054
rect 166586 383498 166822 383734
rect 166586 347818 166822 348054
rect 166586 347498 166822 347734
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 170186 387418 170422 387654
rect 170186 387098 170422 387334
rect 170186 351418 170422 351654
rect 170186 351098 170422 351334
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 191786 710242 192022 710478
rect 191786 709922 192022 710158
rect 188186 708362 188422 708598
rect 188186 708042 188422 708278
rect 184586 706482 184822 706718
rect 184586 706162 184822 706398
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 173786 391018 174022 391254
rect 173786 390698 174022 390934
rect 173786 355018 174022 355254
rect 173786 354698 174022 354934
rect 173786 319018 174022 319254
rect 173786 318698 174022 318934
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 184586 401818 184822 402054
rect 184586 401498 184822 401734
rect 184586 365818 184822 366054
rect 184586 365498 184822 365734
rect 184586 329818 184822 330054
rect 184586 329498 184822 329734
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 188186 405418 188422 405654
rect 188186 405098 188422 405334
rect 188186 369418 188422 369654
rect 188186 369098 188422 369334
rect 188186 333418 188422 333654
rect 188186 333098 188422 333334
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 209786 711182 210022 711418
rect 209786 710862 210022 711098
rect 206186 709302 206422 709538
rect 206186 708982 206422 709218
rect 202586 707422 202822 707658
rect 202586 707102 202822 707338
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 191786 409018 192022 409254
rect 191786 408698 192022 408934
rect 191786 373018 192022 373254
rect 191786 372698 192022 372934
rect 191786 337018 192022 337254
rect 191786 336698 192022 336934
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 198986 560218 199222 560454
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 227786 710242 228022 710478
rect 227786 709922 228022 710158
rect 224186 708362 224422 708598
rect 224186 708042 224422 708278
rect 220586 706482 220822 706718
rect 220586 706162 220822 706398
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 198986 559898 199222 560134
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 203951 542218 204187 542454
rect 203951 541898 204187 542134
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 206917 524218 207153 524454
rect 206917 523898 207153 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 245786 711182 246022 711418
rect 245786 710862 246022 711098
rect 242186 709302 242422 709538
rect 242186 708982 242422 709218
rect 238586 707422 238822 707658
rect 238586 707102 238822 707338
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 238586 419818 238822 420054
rect 238586 419498 238822 419734
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 242186 423418 242422 423654
rect 242186 423098 242422 423334
rect 263786 710242 264022 710478
rect 263786 709922 264022 710158
rect 260186 708362 260422 708598
rect 260186 708042 260422 708278
rect 256586 706482 256822 706718
rect 256586 706162 256822 706398
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 260186 477418 260422 477654
rect 260186 477098 260422 477334
rect 260186 441418 260422 441654
rect 260186 441098 260422 441334
rect 281786 711182 282022 711418
rect 281786 710862 282022 711098
rect 278186 709302 278422 709538
rect 278186 708982 278422 709218
rect 274586 707422 274822 707658
rect 274586 707102 274822 707338
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 263786 481018 264022 481254
rect 263786 480698 264022 480934
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 204250 398218 204486 398454
rect 204250 397898 204486 398134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 219610 380218 219846 380454
rect 219610 379898 219846 380134
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 204250 362218 204486 362454
rect 204250 361898 204486 362134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 219610 344218 219846 344454
rect 219610 343898 219846 344134
rect 270986 344218 271222 344454
rect 270986 343898 271222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 209786 319018 210022 319254
rect 209786 318698 210022 318934
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 220586 329818 220822 330054
rect 220586 329498 220822 329734
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 224186 333418 224422 333654
rect 224186 333098 224422 333334
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 227786 337018 228022 337254
rect 227786 336698 228022 336934
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 245786 319018 246022 319254
rect 245786 318698 246022 318934
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 256586 329818 256822 330054
rect 256586 329498 256822 329734
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 260186 333418 260422 333654
rect 260186 333098 260422 333334
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 263786 337018 264022 337254
rect 263786 336698 264022 336934
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 274586 419818 274822 420054
rect 274586 419498 274822 419734
rect 274586 383818 274822 384054
rect 274586 383498 274822 383734
rect 274586 347818 274822 348054
rect 274586 347498 274822 347734
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 278186 459418 278422 459654
rect 278186 459098 278422 459334
rect 278186 423418 278422 423654
rect 278186 423098 278422 423334
rect 278186 387418 278422 387654
rect 278186 387098 278422 387334
rect 278186 351418 278422 351654
rect 278186 351098 278422 351334
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 299786 710242 300022 710478
rect 299786 709922 300022 710158
rect 296186 708362 296422 708598
rect 296186 708042 296422 708278
rect 292586 706482 292822 706718
rect 292586 706162 292822 706398
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 281786 463018 282022 463254
rect 281786 462698 282022 462934
rect 281786 427018 282022 427254
rect 281786 426698 282022 426934
rect 281786 391018 282022 391254
rect 281786 390698 282022 390934
rect 281786 355018 282022 355254
rect 281786 354698 282022 354934
rect 281786 319018 282022 319254
rect 281786 318698 282022 318934
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 317786 711182 318022 711418
rect 317786 710862 318022 711098
rect 314186 709302 314422 709538
rect 314186 708982 314422 709218
rect 310586 707422 310822 707658
rect 310586 707102 310822 707338
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 335786 710242 336022 710478
rect 335786 709922 336022 710158
rect 332186 708362 332422 708598
rect 332186 708042 332422 708278
rect 328586 706482 328822 706718
rect 328586 706162 328822 706398
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 353786 711182 354022 711418
rect 353786 710862 354022 711098
rect 350186 709302 350422 709538
rect 350186 708982 350422 709218
rect 346586 707422 346822 707658
rect 346586 707102 346822 707338
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 371786 710242 372022 710478
rect 371786 709922 372022 710158
rect 368186 708362 368422 708598
rect 368186 708042 368422 708278
rect 364586 706482 364822 706718
rect 364586 706162 364822 706398
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 389786 711182 390022 711418
rect 389786 710862 390022 711098
rect 386186 709302 386422 709538
rect 386186 708982 386422 709218
rect 382586 707422 382822 707658
rect 382586 707102 382822 707338
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 319610 560218 319846 560454
rect 319610 559898 319846 560134
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 304250 542218 304486 542454
rect 304250 541898 304486 542134
rect 319610 524218 319846 524454
rect 319610 523898 319846 524134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 304250 506218 304486 506454
rect 304250 505898 304486 506134
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 346586 383818 346822 384054
rect 346586 383498 346822 383734
rect 346586 347818 346822 348054
rect 346586 347498 346822 347734
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 350186 387418 350422 387654
rect 350186 387098 350422 387334
rect 350186 351418 350422 351654
rect 350186 351098 350422 351334
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 353786 391018 354022 391254
rect 353786 390698 354022 390934
rect 353786 355018 354022 355254
rect 353786 354698 354022 354934
rect 353786 319018 354022 319254
rect 353786 318698 354022 318934
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 364586 401818 364822 402054
rect 364586 401498 364822 401734
rect 364586 365818 364822 366054
rect 364586 365498 364822 365734
rect 364586 329818 364822 330054
rect 364586 329498 364822 329734
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 368186 405418 368422 405654
rect 368186 405098 368422 405334
rect 368186 369418 368422 369654
rect 368186 369098 368422 369334
rect 368186 333418 368422 333654
rect 368186 333098 368422 333334
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 371786 409018 372022 409254
rect 371786 408698 372022 408934
rect 371786 373018 372022 373254
rect 371786 372698 372022 372934
rect 371786 337018 372022 337254
rect 371786 336698 372022 336934
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 382586 383818 382822 384054
rect 382586 383498 382822 383734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 386186 387418 386422 387654
rect 386186 387098 386422 387334
rect 407786 710242 408022 710478
rect 407786 709922 408022 710158
rect 404186 708362 404422 708598
rect 404186 708042 404422 708278
rect 400586 706482 400822 706718
rect 400586 706162 400822 706398
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 389786 391018 390022 391254
rect 389786 390698 390022 390934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 425786 711182 426022 711418
rect 425786 710862 426022 711098
rect 422186 709302 422422 709538
rect 422186 708982 422422 709218
rect 418586 707422 418822 707658
rect 418586 707102 418822 707338
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 394646 380218 394882 380454
rect 394646 379898 394882 380134
rect 389816 362218 390052 362454
rect 389816 361898 390052 362134
rect 382586 347818 382822 348054
rect 382586 347498 382822 347734
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 389786 319018 390022 319254
rect 389786 318698 390022 318934
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 443786 710242 444022 710478
rect 443786 709922 444022 710158
rect 440186 708362 440422 708598
rect 440186 708042 440422 708278
rect 436586 706482 436822 706718
rect 436586 706162 436822 706398
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 138250 182218 138486 182454
rect 138250 181898 138486 182134
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 153610 164218 153846 164454
rect 153610 163898 153846 164134
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 138250 146218 138486 146454
rect 138250 145898 138486 146134
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 153610 128218 153846 128454
rect 153610 127898 153846 128134
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3402 130822 -3166
rect 130586 -3722 130822 -3486
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5282 134422 -5046
rect 134186 -5602 134422 -5366
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6222 120022 -5986
rect 119786 -6542 120022 -6306
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2462 148822 -2226
rect 148586 -2782 148822 -2546
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4342 152422 -4106
rect 152186 -4662 152422 -4426
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7162 138022 -6926
rect 137786 -7482 138022 -7246
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3402 166822 -3166
rect 166586 -3722 166822 -3486
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5282 170422 -5046
rect 170186 -5602 170422 -5366
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6222 156022 -5986
rect 155786 -6542 156022 -6306
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2462 184822 -2226
rect 184586 -2782 184822 -2546
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4342 188422 -4106
rect 188186 -4662 188422 -4426
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7162 174022 -6926
rect 173786 -7482 174022 -7246
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3402 202822 -3166
rect 202586 -3722 202822 -3486
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5282 206422 -5046
rect 206186 -5602 206422 -5366
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6222 192022 -5986
rect 191786 -6542 192022 -6306
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2462 220822 -2226
rect 220586 -2782 220822 -2546
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4342 224422 -4106
rect 224186 -4662 224422 -4426
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7162 210022 -6926
rect 209786 -7482 210022 -7246
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3402 238822 -3166
rect 238586 -3722 238822 -3486
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5282 242422 -5046
rect 242186 -5602 242422 -5366
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6222 228022 -5986
rect 227786 -6542 228022 -6306
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2462 256822 -2226
rect 256586 -2782 256822 -2546
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4342 260422 -4106
rect 260186 -4662 260422 -4426
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7162 246022 -6926
rect 245786 -7482 246022 -7246
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3402 274822 -3166
rect 274586 -3722 274822 -3486
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5282 278422 -5046
rect 278186 -5602 278422 -5366
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6222 264022 -5986
rect 263786 -6542 264022 -6306
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2462 292822 -2226
rect 292586 -2782 292822 -2546
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4342 296422 -4106
rect 296186 -4662 296422 -4426
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7162 282022 -6926
rect 281786 -7482 282022 -7246
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3402 310822 -3166
rect 310586 -3722 310822 -3486
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5282 314422 -5046
rect 314186 -5602 314422 -5366
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6222 300022 -5986
rect 299786 -6542 300022 -6306
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2462 328822 -2226
rect 328586 -2782 328822 -2546
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4342 332422 -4106
rect 332186 -4662 332422 -4426
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7162 318022 -6926
rect 317786 -7482 318022 -7246
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3402 346822 -3166
rect 346586 -3722 346822 -3486
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5282 350422 -5046
rect 350186 -5602 350422 -5366
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6222 336022 -5986
rect 335786 -6542 336022 -6306
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2462 364822 -2226
rect 364586 -2782 364822 -2546
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4342 368422 -4106
rect 368186 -4662 368422 -4426
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7162 354022 -6926
rect 353786 -7482 354022 -7246
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 382586 -3402 382822 -3166
rect 382586 -3722 382822 -3486
rect 386186 -5282 386422 -5046
rect 386186 -5602 386422 -5366
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6222 372022 -5986
rect 371786 -6542 372022 -6306
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2462 400822 -2226
rect 400586 -2782 400822 -2546
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4342 404422 -4106
rect 404186 -4662 404422 -4426
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7162 390022 -6926
rect 389786 -7482 390022 -7246
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3402 418822 -3166
rect 418586 -3722 418822 -3486
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5282 422422 -5046
rect 422186 -5602 422422 -5366
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6222 408022 -5986
rect 407786 -6542 408022 -6306
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2462 436822 -2226
rect 436586 -2782 436822 -2546
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4342 440422 -4106
rect 440186 -4662 440422 -4426
rect 461786 711182 462022 711418
rect 461786 710862 462022 711098
rect 458186 709302 458422 709538
rect 458186 708982 458422 709218
rect 454586 707422 454822 707658
rect 454586 707102 454822 707338
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7162 426022 -6926
rect 425786 -7482 426022 -7246
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3402 454822 -3166
rect 454586 -3722 454822 -3486
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 479786 710242 480022 710478
rect 479786 709922 480022 710158
rect 476186 708362 476422 708598
rect 476186 708042 476422 708278
rect 472586 706482 472822 706718
rect 472586 706162 472822 706398
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 497786 711182 498022 711418
rect 497786 710862 498022 711098
rect 494186 709302 494422 709538
rect 494186 708982 494422 709218
rect 490586 707422 490822 707658
rect 490586 707102 490822 707338
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 515786 710242 516022 710478
rect 515786 709922 516022 710158
rect 512186 708362 512422 708598
rect 512186 708042 512422 708278
rect 508586 706482 508822 706718
rect 508586 706162 508822 706398
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 485480 542218 485716 542454
rect 485480 541898 485716 542134
rect 490540 524218 490776 524454
rect 490540 523898 490776 524134
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 479610 380218 479846 380454
rect 479610 379898 479846 380134
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 464250 362218 464486 362454
rect 464250 361898 464486 362134
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 479610 344218 479846 344454
rect 479610 343898 479846 344134
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5282 458422 -5046
rect 458186 -5602 458422 -5366
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6222 444022 -5986
rect 443786 -6542 444022 -6306
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2462 472822 -2226
rect 472586 -2782 472822 -2546
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4342 476422 -4106
rect 476186 -4662 476422 -4426
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7162 462022 -6926
rect 461786 -7482 462022 -7246
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3402 490822 -3166
rect 490586 -3722 490822 -3486
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5282 494422 -5046
rect 494186 -5602 494422 -5366
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6222 480022 -5986
rect 479786 -6542 480022 -6306
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2462 508822 -2226
rect 508586 -2782 508822 -2546
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4342 512422 -4106
rect 512186 -4662 512422 -4426
rect 533786 711182 534022 711418
rect 533786 710862 534022 711098
rect 530186 709302 530422 709538
rect 530186 708982 530422 709218
rect 526586 707422 526822 707658
rect 526586 707102 526822 707338
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7162 498022 -6926
rect 497786 -7482 498022 -7246
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3402 526822 -3166
rect 526586 -3722 526822 -3486
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5282 530422 -5046
rect 530186 -5602 530422 -5366
rect 551786 710242 552022 710478
rect 551786 709922 552022 710158
rect 548186 708362 548422 708598
rect 548186 708042 548422 708278
rect 544586 706482 544822 706718
rect 544586 706162 544822 706398
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6222 516022 -5986
rect 515786 -6542 516022 -6306
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2462 544822 -2226
rect 544586 -2782 544822 -2546
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4342 548422 -4106
rect 548186 -4662 548422 -4426
rect 569786 711182 570022 711418
rect 569786 710862 570022 711098
rect 566186 709302 566422 709538
rect 566186 708982 566422 709218
rect 562586 707422 562822 707658
rect 562586 707102 562822 707338
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7162 534022 -6926
rect 533786 -7482 534022 -7246
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3402 562822 -3166
rect 562586 -3722 562822 -3486
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5282 566422 -5046
rect 566186 -5602 566422 -5366
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 580586 706482 580822 706718
rect 580586 706162 580822 706398
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6222 552022 -5986
rect 551786 -6542 552022 -6306
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 689818 587618 690054
rect 587382 689498 587618 689734
rect 587382 653818 587618 654054
rect 587382 653498 587618 653734
rect 587382 617818 587618 618054
rect 587382 617498 587618 617734
rect 587382 581818 587618 582054
rect 587382 581498 587618 581734
rect 587382 545818 587618 546054
rect 587382 545498 587618 545734
rect 587382 509818 587618 510054
rect 587382 509498 587618 509734
rect 587382 473818 587618 474054
rect 587382 473498 587618 473734
rect 587382 437818 587618 438054
rect 587382 437498 587618 437734
rect 587382 401818 587618 402054
rect 587382 401498 587618 401734
rect 587382 365818 587618 366054
rect 587382 365498 587618 365734
rect 587382 329818 587618 330054
rect 587382 329498 587618 329734
rect 587382 293818 587618 294054
rect 587382 293498 587618 293734
rect 587382 257818 587618 258054
rect 587382 257498 587618 257734
rect 587382 221818 587618 222054
rect 587382 221498 587618 221734
rect 587382 185818 587618 186054
rect 587382 185498 587618 185734
rect 587382 149818 587618 150054
rect 587382 149498 587618 149734
rect 587382 113818 587618 114054
rect 587382 113498 587618 113734
rect 587382 77818 587618 78054
rect 587382 77498 587618 77734
rect 587382 41818 587618 42054
rect 587382 41498 587618 41734
rect 587382 5818 587618 6054
rect 587382 5498 587618 5734
rect 580586 -2462 580822 -2226
rect 580586 -2782 580822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 671818 588558 672054
rect 588322 671498 588558 671734
rect 588322 635818 588558 636054
rect 588322 635498 588558 635734
rect 588322 599818 588558 600054
rect 588322 599498 588558 599734
rect 588322 563818 588558 564054
rect 588322 563498 588558 563734
rect 588322 527818 588558 528054
rect 588322 527498 588558 527734
rect 588322 491818 588558 492054
rect 588322 491498 588558 491734
rect 588322 455818 588558 456054
rect 588322 455498 588558 455734
rect 588322 419818 588558 420054
rect 588322 419498 588558 419734
rect 588322 383818 588558 384054
rect 588322 383498 588558 383734
rect 588322 347818 588558 348054
rect 588322 347498 588558 347734
rect 588322 311818 588558 312054
rect 588322 311498 588558 311734
rect 588322 275818 588558 276054
rect 588322 275498 588558 275734
rect 588322 239818 588558 240054
rect 588322 239498 588558 239734
rect 588322 203818 588558 204054
rect 588322 203498 588558 203734
rect 588322 167818 588558 168054
rect 588322 167498 588558 167734
rect 588322 131818 588558 132054
rect 588322 131498 588558 131734
rect 588322 95818 588558 96054
rect 588322 95498 588558 95734
rect 588322 59818 588558 60054
rect 588322 59498 588558 59734
rect 588322 23818 588558 24054
rect 588322 23498 588558 23734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 693418 589498 693654
rect 589262 693098 589498 693334
rect 589262 657418 589498 657654
rect 589262 657098 589498 657334
rect 589262 621418 589498 621654
rect 589262 621098 589498 621334
rect 589262 585418 589498 585654
rect 589262 585098 589498 585334
rect 589262 549418 589498 549654
rect 589262 549098 589498 549334
rect 589262 513418 589498 513654
rect 589262 513098 589498 513334
rect 589262 477418 589498 477654
rect 589262 477098 589498 477334
rect 589262 441418 589498 441654
rect 589262 441098 589498 441334
rect 589262 405418 589498 405654
rect 589262 405098 589498 405334
rect 589262 369418 589498 369654
rect 589262 369098 589498 369334
rect 589262 333418 589498 333654
rect 589262 333098 589498 333334
rect 589262 297418 589498 297654
rect 589262 297098 589498 297334
rect 589262 261418 589498 261654
rect 589262 261098 589498 261334
rect 589262 225418 589498 225654
rect 589262 225098 589498 225334
rect 589262 189418 589498 189654
rect 589262 189098 589498 189334
rect 589262 153418 589498 153654
rect 589262 153098 589498 153334
rect 589262 117418 589498 117654
rect 589262 117098 589498 117334
rect 589262 81418 589498 81654
rect 589262 81098 589498 81334
rect 589262 45418 589498 45654
rect 589262 45098 589498 45334
rect 589262 9418 589498 9654
rect 589262 9098 589498 9334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 675418 590438 675654
rect 590202 675098 590438 675334
rect 590202 639418 590438 639654
rect 590202 639098 590438 639334
rect 590202 603418 590438 603654
rect 590202 603098 590438 603334
rect 590202 567418 590438 567654
rect 590202 567098 590438 567334
rect 590202 531418 590438 531654
rect 590202 531098 590438 531334
rect 590202 495418 590438 495654
rect 590202 495098 590438 495334
rect 590202 459418 590438 459654
rect 590202 459098 590438 459334
rect 590202 423418 590438 423654
rect 590202 423098 590438 423334
rect 590202 387418 590438 387654
rect 590202 387098 590438 387334
rect 590202 351418 590438 351654
rect 590202 351098 590438 351334
rect 590202 315418 590438 315654
rect 590202 315098 590438 315334
rect 590202 279418 590438 279654
rect 590202 279098 590438 279334
rect 590202 243418 590438 243654
rect 590202 243098 590438 243334
rect 590202 207418 590438 207654
rect 590202 207098 590438 207334
rect 590202 171418 590438 171654
rect 590202 171098 590438 171334
rect 590202 135418 590438 135654
rect 590202 135098 590438 135334
rect 590202 99418 590438 99654
rect 590202 99098 590438 99334
rect 590202 63418 590438 63654
rect 590202 63098 590438 63334
rect 590202 27418 590438 27654
rect 590202 27098 590438 27334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 697018 591378 697254
rect 591142 696698 591378 696934
rect 591142 661018 591378 661254
rect 591142 660698 591378 660934
rect 591142 625018 591378 625254
rect 591142 624698 591378 624934
rect 591142 589018 591378 589254
rect 591142 588698 591378 588934
rect 591142 553018 591378 553254
rect 591142 552698 591378 552934
rect 591142 517018 591378 517254
rect 591142 516698 591378 516934
rect 591142 481018 591378 481254
rect 591142 480698 591378 480934
rect 591142 445018 591378 445254
rect 591142 444698 591378 444934
rect 591142 409018 591378 409254
rect 591142 408698 591378 408934
rect 591142 373018 591378 373254
rect 591142 372698 591378 372934
rect 591142 337018 591378 337254
rect 591142 336698 591378 336934
rect 591142 301018 591378 301254
rect 591142 300698 591378 300934
rect 591142 265018 591378 265254
rect 591142 264698 591378 264934
rect 591142 229018 591378 229254
rect 591142 228698 591378 228934
rect 591142 193018 591378 193254
rect 591142 192698 591378 192934
rect 591142 157018 591378 157254
rect 591142 156698 591378 156934
rect 591142 121018 591378 121254
rect 591142 120698 591378 120934
rect 591142 85018 591378 85254
rect 591142 84698 591378 84934
rect 591142 49018 591378 49254
rect 591142 48698 591378 48934
rect 591142 13018 591378 13254
rect 591142 12698 591378 12934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 679018 592318 679254
rect 592082 678698 592318 678934
rect 592082 643018 592318 643254
rect 592082 642698 592318 642934
rect 592082 607018 592318 607254
rect 592082 606698 592318 606934
rect 592082 571018 592318 571254
rect 592082 570698 592318 570934
rect 592082 535018 592318 535254
rect 592082 534698 592318 534934
rect 592082 499018 592318 499254
rect 592082 498698 592318 498934
rect 592082 463018 592318 463254
rect 592082 462698 592318 462934
rect 592082 427018 592318 427254
rect 592082 426698 592318 426934
rect 592082 391018 592318 391254
rect 592082 390698 592318 390934
rect 592082 355018 592318 355254
rect 592082 354698 592318 354934
rect 592082 319018 592318 319254
rect 592082 318698 592318 318934
rect 592082 283018 592318 283254
rect 592082 282698 592318 282934
rect 592082 247018 592318 247254
rect 592082 246698 592318 246934
rect 592082 211018 592318 211254
rect 592082 210698 592318 210934
rect 592082 175018 592318 175254
rect 592082 174698 592318 174934
rect 592082 139018 592318 139254
rect 592082 138698 592318 138934
rect 592082 103018 592318 103254
rect 592082 102698 592318 102934
rect 592082 67018 592318 67254
rect 592082 66698 592318 66934
rect 592082 31018 592318 31254
rect 592082 30698 592318 30934
rect 569786 -7162 570022 -6926
rect 569786 -7482 570022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 29786 711418
rect 30022 711182 65786 711418
rect 66022 711182 101786 711418
rect 102022 711182 137786 711418
rect 138022 711182 173786 711418
rect 174022 711182 209786 711418
rect 210022 711182 245786 711418
rect 246022 711182 281786 711418
rect 282022 711182 317786 711418
rect 318022 711182 353786 711418
rect 354022 711182 389786 711418
rect 390022 711182 425786 711418
rect 426022 711182 461786 711418
rect 462022 711182 497786 711418
rect 498022 711182 533786 711418
rect 534022 711182 569786 711418
rect 570022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 29786 711098
rect 30022 710862 65786 711098
rect 66022 710862 101786 711098
rect 102022 710862 137786 711098
rect 138022 710862 173786 711098
rect 174022 710862 209786 711098
rect 210022 710862 245786 711098
rect 246022 710862 281786 711098
rect 282022 710862 317786 711098
rect 318022 710862 353786 711098
rect 354022 710862 389786 711098
rect 390022 710862 425786 711098
rect 426022 710862 461786 711098
rect 462022 710862 497786 711098
rect 498022 710862 533786 711098
rect 534022 710862 569786 711098
rect 570022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 11786 710478
rect 12022 710242 47786 710478
rect 48022 710242 83786 710478
rect 84022 710242 119786 710478
rect 120022 710242 155786 710478
rect 156022 710242 191786 710478
rect 192022 710242 227786 710478
rect 228022 710242 263786 710478
rect 264022 710242 299786 710478
rect 300022 710242 335786 710478
rect 336022 710242 371786 710478
rect 372022 710242 407786 710478
rect 408022 710242 443786 710478
rect 444022 710242 479786 710478
rect 480022 710242 515786 710478
rect 516022 710242 551786 710478
rect 552022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 11786 710158
rect 12022 709922 47786 710158
rect 48022 709922 83786 710158
rect 84022 709922 119786 710158
rect 120022 709922 155786 710158
rect 156022 709922 191786 710158
rect 192022 709922 227786 710158
rect 228022 709922 263786 710158
rect 264022 709922 299786 710158
rect 300022 709922 335786 710158
rect 336022 709922 371786 710158
rect 372022 709922 407786 710158
rect 408022 709922 443786 710158
rect 444022 709922 479786 710158
rect 480022 709922 515786 710158
rect 516022 709922 551786 710158
rect 552022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 26186 709538
rect 26422 709302 62186 709538
rect 62422 709302 98186 709538
rect 98422 709302 134186 709538
rect 134422 709302 170186 709538
rect 170422 709302 206186 709538
rect 206422 709302 242186 709538
rect 242422 709302 278186 709538
rect 278422 709302 314186 709538
rect 314422 709302 350186 709538
rect 350422 709302 386186 709538
rect 386422 709302 422186 709538
rect 422422 709302 458186 709538
rect 458422 709302 494186 709538
rect 494422 709302 530186 709538
rect 530422 709302 566186 709538
rect 566422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 26186 709218
rect 26422 708982 62186 709218
rect 62422 708982 98186 709218
rect 98422 708982 134186 709218
rect 134422 708982 170186 709218
rect 170422 708982 206186 709218
rect 206422 708982 242186 709218
rect 242422 708982 278186 709218
rect 278422 708982 314186 709218
rect 314422 708982 350186 709218
rect 350422 708982 386186 709218
rect 386422 708982 422186 709218
rect 422422 708982 458186 709218
rect 458422 708982 494186 709218
rect 494422 708982 530186 709218
rect 530422 708982 566186 709218
rect 566422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 8186 708598
rect 8422 708362 44186 708598
rect 44422 708362 80186 708598
rect 80422 708362 116186 708598
rect 116422 708362 152186 708598
rect 152422 708362 188186 708598
rect 188422 708362 224186 708598
rect 224422 708362 260186 708598
rect 260422 708362 296186 708598
rect 296422 708362 332186 708598
rect 332422 708362 368186 708598
rect 368422 708362 404186 708598
rect 404422 708362 440186 708598
rect 440422 708362 476186 708598
rect 476422 708362 512186 708598
rect 512422 708362 548186 708598
rect 548422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 8186 708278
rect 8422 708042 44186 708278
rect 44422 708042 80186 708278
rect 80422 708042 116186 708278
rect 116422 708042 152186 708278
rect 152422 708042 188186 708278
rect 188422 708042 224186 708278
rect 224422 708042 260186 708278
rect 260422 708042 296186 708278
rect 296422 708042 332186 708278
rect 332422 708042 368186 708278
rect 368422 708042 404186 708278
rect 404422 708042 440186 708278
rect 440422 708042 476186 708278
rect 476422 708042 512186 708278
rect 512422 708042 548186 708278
rect 548422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 22586 707658
rect 22822 707422 58586 707658
rect 58822 707422 94586 707658
rect 94822 707422 130586 707658
rect 130822 707422 166586 707658
rect 166822 707422 202586 707658
rect 202822 707422 238586 707658
rect 238822 707422 274586 707658
rect 274822 707422 310586 707658
rect 310822 707422 346586 707658
rect 346822 707422 382586 707658
rect 382822 707422 418586 707658
rect 418822 707422 454586 707658
rect 454822 707422 490586 707658
rect 490822 707422 526586 707658
rect 526822 707422 562586 707658
rect 562822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 22586 707338
rect 22822 707102 58586 707338
rect 58822 707102 94586 707338
rect 94822 707102 130586 707338
rect 130822 707102 166586 707338
rect 166822 707102 202586 707338
rect 202822 707102 238586 707338
rect 238822 707102 274586 707338
rect 274822 707102 310586 707338
rect 310822 707102 346586 707338
rect 346822 707102 382586 707338
rect 382822 707102 418586 707338
rect 418822 707102 454586 707338
rect 454822 707102 490586 707338
rect 490822 707102 526586 707338
rect 526822 707102 562586 707338
rect 562822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 4586 706718
rect 4822 706482 40586 706718
rect 40822 706482 76586 706718
rect 76822 706482 112586 706718
rect 112822 706482 148586 706718
rect 148822 706482 184586 706718
rect 184822 706482 220586 706718
rect 220822 706482 256586 706718
rect 256822 706482 292586 706718
rect 292822 706482 328586 706718
rect 328822 706482 364586 706718
rect 364822 706482 400586 706718
rect 400822 706482 436586 706718
rect 436822 706482 472586 706718
rect 472822 706482 508586 706718
rect 508822 706482 544586 706718
rect 544822 706482 580586 706718
rect 580822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 4586 706398
rect 4822 706162 40586 706398
rect 40822 706162 76586 706398
rect 76822 706162 112586 706398
rect 112822 706162 148586 706398
rect 148822 706162 184586 706398
rect 184822 706162 220586 706398
rect 220822 706162 256586 706398
rect 256822 706162 292586 706398
rect 292822 706162 328586 706398
rect 328822 706162 364586 706398
rect 364822 706162 400586 706398
rect 400822 706162 436586 706398
rect 436822 706162 472586 706398
rect 472822 706162 508586 706398
rect 508822 706162 544586 706398
rect 544822 706162 580586 706398
rect 580822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7636 697276 -7036 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590960 697276 591560 697278
rect -8576 697254 592500 697276
rect -8576 697018 -7454 697254
rect -7218 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591142 697254
rect 591378 697018 592500 697254
rect -8576 696934 592500 697018
rect -8576 696698 -7454 696934
rect -7218 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591142 696934
rect 591378 696698 592500 696934
rect -8576 696676 592500 696698
rect -7636 696674 -7036 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590960 696674 591560 696676
rect -5756 693676 -5156 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589080 693676 589680 693678
rect -6696 693654 590620 693676
rect -6696 693418 -5574 693654
rect -5338 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589262 693654
rect 589498 693418 590620 693654
rect -6696 693334 590620 693418
rect -6696 693098 -5574 693334
rect -5338 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589262 693334
rect 589498 693098 590620 693334
rect -6696 693076 590620 693098
rect -5756 693074 -5156 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589080 693074 589680 693076
rect -3876 690076 -3276 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587200 690076 587800 690078
rect -4816 690054 588740 690076
rect -4816 689818 -3694 690054
rect -3458 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587382 690054
rect 587618 689818 588740 690054
rect -4816 689734 588740 689818
rect -4816 689498 -3694 689734
rect -3458 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587382 689734
rect 587618 689498 588740 689734
rect -4816 689476 588740 689498
rect -3876 689474 -3276 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587200 689474 587800 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8576 679276 -7976 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591900 679276 592500 679278
rect -8576 679254 592500 679276
rect -8576 679018 -8394 679254
rect -8158 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 592082 679254
rect 592318 679018 592500 679254
rect -8576 678934 592500 679018
rect -8576 678698 -8394 678934
rect -8158 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 592082 678934
rect 592318 678698 592500 678934
rect -8576 678676 592500 678698
rect -8576 678674 -7976 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591900 678674 592500 678676
rect -6696 675676 -6096 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 590020 675676 590620 675678
rect -6696 675654 590620 675676
rect -6696 675418 -6514 675654
rect -6278 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590202 675654
rect 590438 675418 590620 675654
rect -6696 675334 590620 675418
rect -6696 675098 -6514 675334
rect -6278 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590202 675334
rect 590438 675098 590620 675334
rect -6696 675076 590620 675098
rect -6696 675074 -6096 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 590020 675074 590620 675076
rect -4816 672076 -4216 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588140 672076 588740 672078
rect -4816 672054 588740 672076
rect -4816 671818 -4634 672054
rect -4398 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588322 672054
rect 588558 671818 588740 672054
rect -4816 671734 588740 671818
rect -4816 671498 -4634 671734
rect -4398 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588322 671734
rect 588558 671498 588740 671734
rect -4816 671476 588740 671498
rect -4816 671474 -4216 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588140 671474 588740 671476
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -7636 661276 -7036 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590960 661276 591560 661278
rect -8576 661254 592500 661276
rect -8576 661018 -7454 661254
rect -7218 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591142 661254
rect 591378 661018 592500 661254
rect -8576 660934 592500 661018
rect -8576 660698 -7454 660934
rect -7218 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591142 660934
rect 591378 660698 592500 660934
rect -8576 660676 592500 660698
rect -7636 660674 -7036 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590960 660674 591560 660676
rect -5756 657676 -5156 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589080 657676 589680 657678
rect -6696 657654 590620 657676
rect -6696 657418 -5574 657654
rect -5338 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589262 657654
rect 589498 657418 590620 657654
rect -6696 657334 590620 657418
rect -6696 657098 -5574 657334
rect -5338 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589262 657334
rect 589498 657098 590620 657334
rect -6696 657076 590620 657098
rect -5756 657074 -5156 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589080 657074 589680 657076
rect -3876 654076 -3276 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587200 654076 587800 654078
rect -4816 654054 588740 654076
rect -4816 653818 -3694 654054
rect -3458 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587382 654054
rect 587618 653818 588740 654054
rect -4816 653734 588740 653818
rect -4816 653498 -3694 653734
rect -3458 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587382 653734
rect 587618 653498 588740 653734
rect -4816 653476 588740 653498
rect -3876 653474 -3276 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587200 653474 587800 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8576 643276 -7976 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591900 643276 592500 643278
rect -8576 643254 592500 643276
rect -8576 643018 -8394 643254
rect -8158 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 592082 643254
rect 592318 643018 592500 643254
rect -8576 642934 592500 643018
rect -8576 642698 -8394 642934
rect -8158 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 592082 642934
rect 592318 642698 592500 642934
rect -8576 642676 592500 642698
rect -8576 642674 -7976 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591900 642674 592500 642676
rect -6696 639676 -6096 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 590020 639676 590620 639678
rect -6696 639654 590620 639676
rect -6696 639418 -6514 639654
rect -6278 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590202 639654
rect 590438 639418 590620 639654
rect -6696 639334 590620 639418
rect -6696 639098 -6514 639334
rect -6278 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590202 639334
rect 590438 639098 590620 639334
rect -6696 639076 590620 639098
rect -6696 639074 -6096 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 590020 639074 590620 639076
rect -4816 636076 -4216 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588140 636076 588740 636078
rect -4816 636054 588740 636076
rect -4816 635818 -4634 636054
rect -4398 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588322 636054
rect 588558 635818 588740 636054
rect -4816 635734 588740 635818
rect -4816 635498 -4634 635734
rect -4398 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588322 635734
rect 588558 635498 588740 635734
rect -4816 635476 588740 635498
rect -4816 635474 -4216 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588140 635474 588740 635476
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -7636 625276 -7036 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590960 625276 591560 625278
rect -8576 625254 592500 625276
rect -8576 625018 -7454 625254
rect -7218 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591142 625254
rect 591378 625018 592500 625254
rect -8576 624934 592500 625018
rect -8576 624698 -7454 624934
rect -7218 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591142 624934
rect 591378 624698 592500 624934
rect -8576 624676 592500 624698
rect -7636 624674 -7036 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590960 624674 591560 624676
rect -5756 621676 -5156 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589080 621676 589680 621678
rect -6696 621654 590620 621676
rect -6696 621418 -5574 621654
rect -5338 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589262 621654
rect 589498 621418 590620 621654
rect -6696 621334 590620 621418
rect -6696 621098 -5574 621334
rect -5338 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589262 621334
rect 589498 621098 590620 621334
rect -6696 621076 590620 621098
rect -5756 621074 -5156 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589080 621074 589680 621076
rect -3876 618076 -3276 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587200 618076 587800 618078
rect -4816 618054 588740 618076
rect -4816 617818 -3694 618054
rect -3458 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587382 618054
rect 587618 617818 588740 618054
rect -4816 617734 588740 617818
rect -4816 617498 -3694 617734
rect -3458 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587382 617734
rect 587618 617498 588740 617734
rect -4816 617476 588740 617498
rect -3876 617474 -3276 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587200 617474 587800 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8576 607276 -7976 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591900 607276 592500 607278
rect -8576 607254 592500 607276
rect -8576 607018 -8394 607254
rect -8158 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 592082 607254
rect 592318 607018 592500 607254
rect -8576 606934 592500 607018
rect -8576 606698 -8394 606934
rect -8158 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 592082 606934
rect 592318 606698 592500 606934
rect -8576 606676 592500 606698
rect -8576 606674 -7976 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591900 606674 592500 606676
rect -6696 603676 -6096 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 590020 603676 590620 603678
rect -6696 603654 590620 603676
rect -6696 603418 -6514 603654
rect -6278 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590202 603654
rect 590438 603418 590620 603654
rect -6696 603334 590620 603418
rect -6696 603098 -6514 603334
rect -6278 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590202 603334
rect 590438 603098 590620 603334
rect -6696 603076 590620 603098
rect -6696 603074 -6096 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 590020 603074 590620 603076
rect -4816 600076 -4216 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588140 600076 588740 600078
rect -4816 600054 588740 600076
rect -4816 599818 -4634 600054
rect -4398 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588322 600054
rect 588558 599818 588740 600054
rect -4816 599734 588740 599818
rect -4816 599498 -4634 599734
rect -4398 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588322 599734
rect 588558 599498 588740 599734
rect -4816 599476 588740 599498
rect -4816 599474 -4216 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588140 599474 588740 599476
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -7636 589276 -7036 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590960 589276 591560 589278
rect -8576 589254 592500 589276
rect -8576 589018 -7454 589254
rect -7218 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591142 589254
rect 591378 589018 592500 589254
rect -8576 588934 592500 589018
rect -8576 588698 -7454 588934
rect -7218 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591142 588934
rect 591378 588698 592500 588934
rect -8576 588676 592500 588698
rect -7636 588674 -7036 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590960 588674 591560 588676
rect -5756 585676 -5156 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589080 585676 589680 585678
rect -6696 585654 590620 585676
rect -6696 585418 -5574 585654
rect -5338 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589262 585654
rect 589498 585418 590620 585654
rect -6696 585334 590620 585418
rect -6696 585098 -5574 585334
rect -5338 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589262 585334
rect 589498 585098 590620 585334
rect -6696 585076 590620 585098
rect -5756 585074 -5156 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589080 585074 589680 585076
rect -3876 582076 -3276 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587200 582076 587800 582078
rect -4816 582054 588740 582076
rect -4816 581818 -3694 582054
rect -3458 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587382 582054
rect 587618 581818 588740 582054
rect -4816 581734 588740 581818
rect -4816 581498 -3694 581734
rect -3458 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587382 581734
rect 587618 581498 588740 581734
rect -4816 581476 588740 581498
rect -3876 581474 -3276 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587200 581474 587800 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8576 571276 -7976 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591900 571276 592500 571278
rect -8576 571254 592500 571276
rect -8576 571018 -8394 571254
rect -8158 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 592082 571254
rect 592318 571018 592500 571254
rect -8576 570934 592500 571018
rect -8576 570698 -8394 570934
rect -8158 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 592082 570934
rect 592318 570698 592500 570934
rect -8576 570676 592500 570698
rect -8576 570674 -7976 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591900 570674 592500 570676
rect -6696 567676 -6096 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 590020 567676 590620 567678
rect -6696 567654 590620 567676
rect -6696 567418 -6514 567654
rect -6278 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590202 567654
rect 590438 567418 590620 567654
rect -6696 567334 590620 567418
rect -6696 567098 -6514 567334
rect -6278 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590202 567334
rect 590438 567098 590620 567334
rect -6696 567076 590620 567098
rect -6696 567074 -6096 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 590020 567074 590620 567076
rect -4816 564076 -4216 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588140 564076 588740 564078
rect -4816 564054 588740 564076
rect -4816 563818 -4634 564054
rect -4398 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588322 564054
rect 588558 563818 588740 564054
rect -4816 563734 588740 563818
rect -4816 563498 -4634 563734
rect -4398 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588322 563734
rect 588558 563498 588740 563734
rect -4816 563476 588740 563498
rect -4816 563474 -4216 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588140 563474 588740 563476
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 319568 560476 319888 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 319610 560454
rect 319846 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 319610 560134
rect 319846 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 319568 559874 319888 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -7636 553276 -7036 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590960 553276 591560 553278
rect -8576 553254 592500 553276
rect -8576 553018 -7454 553254
rect -7218 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591142 553254
rect 591378 553018 592500 553254
rect -8576 552934 592500 553018
rect -8576 552698 -7454 552934
rect -7218 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591142 552934
rect 591378 552698 592500 552934
rect -8576 552676 592500 552698
rect -7636 552674 -7036 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590960 552674 591560 552676
rect -5756 549676 -5156 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589080 549676 589680 549678
rect -6696 549654 590620 549676
rect -6696 549418 -5574 549654
rect -5338 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589262 549654
rect 589498 549418 590620 549654
rect -6696 549334 590620 549418
rect -6696 549098 -5574 549334
rect -5338 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589262 549334
rect 589498 549098 590620 549334
rect -6696 549076 590620 549098
rect -5756 549074 -5156 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589080 549074 589680 549076
rect -3876 546076 -3276 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587200 546076 587800 546078
rect -4816 546054 588740 546076
rect -4816 545818 -3694 546054
rect -3458 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587382 546054
rect 587618 545818 588740 546054
rect -4816 545734 588740 545818
rect -4816 545498 -3694 545734
rect -3458 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587382 545734
rect 587618 545498 588740 545734
rect -4816 545476 588740 545498
rect -3876 545474 -3276 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587200 545474 587800 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 91529 542476 91849 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 203909 542476 204229 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 304208 542476 304528 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 485438 542476 485758 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 91571 542454
rect 91807 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 203951 542454
rect 204187 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 304250 542454
rect 304486 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 485480 542454
rect 485716 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 91571 542134
rect 91807 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 203951 542134
rect 204187 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 304250 542134
rect 304486 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 485480 542134
rect 485716 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 91529 541874 91849 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 203909 541874 204229 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 304208 541874 304528 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 485438 541874 485758 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8576 535276 -7976 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591900 535276 592500 535278
rect -8576 535254 592500 535276
rect -8576 535018 -8394 535254
rect -8158 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 592082 535254
rect 592318 535018 592500 535254
rect -8576 534934 592500 535018
rect -8576 534698 -8394 534934
rect -8158 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 592082 534934
rect 592318 534698 592500 534934
rect -8576 534676 592500 534698
rect -8576 534674 -7976 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591900 534674 592500 534676
rect -6696 531676 -6096 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 590020 531676 590620 531678
rect -6696 531654 590620 531676
rect -6696 531418 -6514 531654
rect -6278 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590202 531654
rect 590438 531418 590620 531654
rect -6696 531334 590620 531418
rect -6696 531098 -6514 531334
rect -6278 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590202 531334
rect 590438 531098 590620 531334
rect -6696 531076 590620 531098
rect -6696 531074 -6096 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 590020 531074 590620 531076
rect -4816 528076 -4216 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588140 528076 588740 528078
rect -4816 528054 588740 528076
rect -4816 527818 -4634 528054
rect -4398 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588322 528054
rect 588558 527818 588740 528054
rect -4816 527734 588740 527818
rect -4816 527498 -4634 527734
rect -4398 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588322 527734
rect 588558 527498 588740 527734
rect -4816 527476 588740 527498
rect -4816 527474 -4216 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588140 527474 588740 527476
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 96113 524476 96433 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 206875 524476 207195 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 319568 524476 319888 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 490498 524476 490818 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 96155 524454
rect 96391 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 206917 524454
rect 207153 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 319610 524454
rect 319846 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 490540 524454
rect 490776 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 96155 524134
rect 96391 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 206917 524134
rect 207153 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 319610 524134
rect 319846 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 490540 524134
rect 490776 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 96113 523874 96433 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 206875 523874 207195 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 319568 523874 319888 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 490498 523874 490818 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586260 523874 586860 523876
rect -7636 517276 -7036 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590960 517276 591560 517278
rect -8576 517254 592500 517276
rect -8576 517018 -7454 517254
rect -7218 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591142 517254
rect 591378 517018 592500 517254
rect -8576 516934 592500 517018
rect -8576 516698 -7454 516934
rect -7218 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591142 516934
rect 591378 516698 592500 516934
rect -8576 516676 592500 516698
rect -7636 516674 -7036 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590960 516674 591560 516676
rect -5756 513676 -5156 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589080 513676 589680 513678
rect -6696 513654 590620 513676
rect -6696 513418 -5574 513654
rect -5338 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589262 513654
rect 589498 513418 590620 513654
rect -6696 513334 590620 513418
rect -6696 513098 -5574 513334
rect -5338 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589262 513334
rect 589498 513098 590620 513334
rect -6696 513076 590620 513098
rect -5756 513074 -5156 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589080 513074 589680 513076
rect -3876 510076 -3276 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587200 510076 587800 510078
rect -4816 510054 588740 510076
rect -4816 509818 -3694 510054
rect -3458 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587382 510054
rect 587618 509818 588740 510054
rect -4816 509734 588740 509818
rect -4816 509498 -3694 509734
rect -3458 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587382 509734
rect 587618 509498 588740 509734
rect -4816 509476 588740 509498
rect -3876 509474 -3276 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587200 509474 587800 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 304208 506476 304528 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 304250 506454
rect 304486 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 304250 506134
rect 304486 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 304208 505874 304528 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8576 499276 -7976 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591900 499276 592500 499278
rect -8576 499254 592500 499276
rect -8576 499018 -8394 499254
rect -8158 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 592082 499254
rect 592318 499018 592500 499254
rect -8576 498934 592500 499018
rect -8576 498698 -8394 498934
rect -8158 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 592082 498934
rect 592318 498698 592500 498934
rect -8576 498676 592500 498698
rect -8576 498674 -7976 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591900 498674 592500 498676
rect -6696 495676 -6096 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 590020 495676 590620 495678
rect -6696 495654 590620 495676
rect -6696 495418 -6514 495654
rect -6278 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590202 495654
rect 590438 495418 590620 495654
rect -6696 495334 590620 495418
rect -6696 495098 -6514 495334
rect -6278 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590202 495334
rect 590438 495098 590620 495334
rect -6696 495076 590620 495098
rect -6696 495074 -6096 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 590020 495074 590620 495076
rect -4816 492076 -4216 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588140 492076 588740 492078
rect -4816 492054 588740 492076
rect -4816 491818 -4634 492054
rect -4398 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588322 492054
rect 588558 491818 588740 492054
rect -4816 491734 588740 491818
rect -4816 491498 -4634 491734
rect -4398 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588322 491734
rect 588558 491498 588740 491734
rect -4816 491476 588740 491498
rect -4816 491474 -4216 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588140 491474 588740 491476
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -7636 481276 -7036 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 263604 481276 264204 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590960 481276 591560 481278
rect -8576 481254 592500 481276
rect -8576 481018 -7454 481254
rect -7218 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 263786 481254
rect 264022 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591142 481254
rect 591378 481018 592500 481254
rect -8576 480934 592500 481018
rect -8576 480698 -7454 480934
rect -7218 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 263786 480934
rect 264022 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591142 480934
rect 591378 480698 592500 480934
rect -8576 480676 592500 480698
rect -7636 480674 -7036 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 263604 480674 264204 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590960 480674 591560 480676
rect -5756 477676 -5156 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 260004 477676 260604 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589080 477676 589680 477678
rect -6696 477654 590620 477676
rect -6696 477418 -5574 477654
rect -5338 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 260186 477654
rect 260422 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589262 477654
rect 589498 477418 590620 477654
rect -6696 477334 590620 477418
rect -6696 477098 -5574 477334
rect -5338 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 260186 477334
rect 260422 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589262 477334
rect 589498 477098 590620 477334
rect -6696 477076 590620 477098
rect -5756 477074 -5156 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 260004 477074 260604 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589080 477074 589680 477076
rect -3876 474076 -3276 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587200 474076 587800 474078
rect -4816 474054 588740 474076
rect -4816 473818 -3694 474054
rect -3458 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587382 474054
rect 587618 473818 588740 474054
rect -4816 473734 588740 473818
rect -4816 473498 -3694 473734
rect -3458 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587382 473734
rect 587618 473498 588740 473734
rect -4816 473476 588740 473498
rect -3876 473474 -3276 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587200 473474 587800 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8576 463276 -7976 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 281604 463276 282204 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591900 463276 592500 463278
rect -8576 463254 592500 463276
rect -8576 463018 -8394 463254
rect -8158 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 281786 463254
rect 282022 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 592082 463254
rect 592318 463018 592500 463254
rect -8576 462934 592500 463018
rect -8576 462698 -8394 462934
rect -8158 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 281786 462934
rect 282022 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 592082 462934
rect 592318 462698 592500 462934
rect -8576 462676 592500 462698
rect -8576 462674 -7976 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 281604 462674 282204 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591900 462674 592500 462676
rect -6696 459676 -6096 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 278004 459676 278604 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 590020 459676 590620 459678
rect -6696 459654 590620 459676
rect -6696 459418 -6514 459654
rect -6278 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 278186 459654
rect 278422 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590202 459654
rect 590438 459418 590620 459654
rect -6696 459334 590620 459418
rect -6696 459098 -6514 459334
rect -6278 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 278186 459334
rect 278422 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590202 459334
rect 590438 459098 590620 459334
rect -6696 459076 590620 459098
rect -6696 459074 -6096 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 278004 459074 278604 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 590020 459074 590620 459076
rect -4816 456076 -4216 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588140 456076 588740 456078
rect -4816 456054 588740 456076
rect -4816 455818 -4634 456054
rect -4398 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588322 456054
rect 588558 455818 588740 456054
rect -4816 455734 588740 455818
rect -4816 455498 -4634 455734
rect -4398 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588322 455734
rect 588558 455498 588740 455734
rect -4816 455476 588740 455498
rect -4816 455474 -4216 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588140 455474 588740 455476
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -7636 445276 -7036 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590960 445276 591560 445278
rect -8576 445254 592500 445276
rect -8576 445018 -7454 445254
rect -7218 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591142 445254
rect 591378 445018 592500 445254
rect -8576 444934 592500 445018
rect -8576 444698 -7454 444934
rect -7218 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591142 444934
rect 591378 444698 592500 444934
rect -8576 444676 592500 444698
rect -7636 444674 -7036 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590960 444674 591560 444676
rect -5756 441676 -5156 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 260004 441676 260604 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589080 441676 589680 441678
rect -6696 441654 590620 441676
rect -6696 441418 -5574 441654
rect -5338 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 260186 441654
rect 260422 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589262 441654
rect 589498 441418 590620 441654
rect -6696 441334 590620 441418
rect -6696 441098 -5574 441334
rect -5338 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 260186 441334
rect 260422 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589262 441334
rect 589498 441098 590620 441334
rect -6696 441076 590620 441098
rect -5756 441074 -5156 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 260004 441074 260604 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589080 441074 589680 441076
rect -3876 438076 -3276 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587200 438076 587800 438078
rect -4816 438054 588740 438076
rect -4816 437818 -3694 438054
rect -3458 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587382 438054
rect 587618 437818 588740 438054
rect -4816 437734 588740 437818
rect -4816 437498 -3694 437734
rect -3458 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587382 437734
rect 587618 437498 588740 437734
rect -4816 437476 588740 437498
rect -3876 437474 -3276 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587200 437474 587800 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8576 427276 -7976 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 281604 427276 282204 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591900 427276 592500 427278
rect -8576 427254 592500 427276
rect -8576 427018 -8394 427254
rect -8158 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 281786 427254
rect 282022 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 592082 427254
rect 592318 427018 592500 427254
rect -8576 426934 592500 427018
rect -8576 426698 -8394 426934
rect -8158 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 281786 426934
rect 282022 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 592082 426934
rect 592318 426698 592500 426934
rect -8576 426676 592500 426698
rect -8576 426674 -7976 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 281604 426674 282204 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591900 426674 592500 426676
rect -6696 423676 -6096 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 278004 423676 278604 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 590020 423676 590620 423678
rect -6696 423654 590620 423676
rect -6696 423418 -6514 423654
rect -6278 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 278186 423654
rect 278422 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590202 423654
rect 590438 423418 590620 423654
rect -6696 423334 590620 423418
rect -6696 423098 -6514 423334
rect -6278 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 278186 423334
rect 278422 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590202 423334
rect 590438 423098 590620 423334
rect -6696 423076 590620 423098
rect -6696 423074 -6096 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 278004 423074 278604 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 590020 423074 590620 423076
rect -4816 420076 -4216 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 238404 420076 239004 420078
rect 274404 420076 275004 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588140 420076 588740 420078
rect -4816 420054 588740 420076
rect -4816 419818 -4634 420054
rect -4398 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 238586 420054
rect 238822 419818 274586 420054
rect 274822 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588322 420054
rect 588558 419818 588740 420054
rect -4816 419734 588740 419818
rect -4816 419498 -4634 419734
rect -4398 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 238586 419734
rect 238822 419498 274586 419734
rect 274822 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588322 419734
rect 588558 419498 588740 419734
rect -4816 419476 588740 419498
rect -4816 419474 -4216 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 238404 419474 239004 419476
rect 274404 419474 275004 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588140 419474 588740 419476
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect -7636 409276 -7036 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 155604 409276 156204 409278
rect 191604 409276 192204 409278
rect 299604 409276 300204 409278
rect 335604 409276 336204 409278
rect 371604 409276 372204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590960 409276 591560 409278
rect -8576 409254 592500 409276
rect -8576 409018 -7454 409254
rect -7218 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 155786 409254
rect 156022 409018 191786 409254
rect 192022 409018 299786 409254
rect 300022 409018 335786 409254
rect 336022 409018 371786 409254
rect 372022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591142 409254
rect 591378 409018 592500 409254
rect -8576 408934 592500 409018
rect -8576 408698 -7454 408934
rect -7218 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 155786 408934
rect 156022 408698 191786 408934
rect 192022 408698 299786 408934
rect 300022 408698 335786 408934
rect 336022 408698 371786 408934
rect 372022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591142 408934
rect 591378 408698 592500 408934
rect -8576 408676 592500 408698
rect -7636 408674 -7036 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 155604 408674 156204 408676
rect 191604 408674 192204 408676
rect 299604 408674 300204 408676
rect 335604 408674 336204 408676
rect 371604 408674 372204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590960 408674 591560 408676
rect -5756 405676 -5156 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 188004 405676 188604 405678
rect 296004 405676 296604 405678
rect 332004 405676 332604 405678
rect 368004 405676 368604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589080 405676 589680 405678
rect -6696 405654 590620 405676
rect -6696 405418 -5574 405654
rect -5338 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 188186 405654
rect 188422 405418 296186 405654
rect 296422 405418 332186 405654
rect 332422 405418 368186 405654
rect 368422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589262 405654
rect 589498 405418 590620 405654
rect -6696 405334 590620 405418
rect -6696 405098 -5574 405334
rect -5338 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 188186 405334
rect 188422 405098 296186 405334
rect 296422 405098 332186 405334
rect 332422 405098 368186 405334
rect 368422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589262 405334
rect 589498 405098 590620 405334
rect -6696 405076 590620 405098
rect -5756 405074 -5156 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 188004 405074 188604 405076
rect 296004 405074 296604 405076
rect 332004 405074 332604 405076
rect 368004 405074 368604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589080 405074 589680 405076
rect -3876 402076 -3276 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 184404 402076 185004 402078
rect 292404 402076 293004 402078
rect 328404 402076 329004 402078
rect 364404 402076 365004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587200 402076 587800 402078
rect -4816 402054 588740 402076
rect -4816 401818 -3694 402054
rect -3458 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 184586 402054
rect 184822 401818 292586 402054
rect 292822 401818 328586 402054
rect 328822 401818 364586 402054
rect 364822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587382 402054
rect 587618 401818 588740 402054
rect -4816 401734 588740 401818
rect -4816 401498 -3694 401734
rect -3458 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 184586 401734
rect 184822 401498 292586 401734
rect 292822 401498 328586 401734
rect 328822 401498 364586 401734
rect 364822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587382 401734
rect 587618 401498 588740 401734
rect -4816 401476 588740 401498
rect -3876 401474 -3276 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 184404 401474 185004 401476
rect 292404 401474 293004 401476
rect 328404 401474 329004 401476
rect 364404 401474 365004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587200 401474 587800 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 204208 398476 204528 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 204250 398454
rect 204486 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 204250 398134
rect 204486 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 204208 397874 204528 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8576 391276 -7976 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 137604 391276 138204 391278
rect 173604 391276 174204 391278
rect 281604 391276 282204 391278
rect 317604 391276 318204 391278
rect 353604 391276 354204 391278
rect 389604 391276 390204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591900 391276 592500 391278
rect -8576 391254 592500 391276
rect -8576 391018 -8394 391254
rect -8158 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 137786 391254
rect 138022 391018 173786 391254
rect 174022 391018 281786 391254
rect 282022 391018 317786 391254
rect 318022 391018 353786 391254
rect 354022 391018 389786 391254
rect 390022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 592082 391254
rect 592318 391018 592500 391254
rect -8576 390934 592500 391018
rect -8576 390698 -8394 390934
rect -8158 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 137786 390934
rect 138022 390698 173786 390934
rect 174022 390698 281786 390934
rect 282022 390698 317786 390934
rect 318022 390698 353786 390934
rect 354022 390698 389786 390934
rect 390022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 592082 390934
rect 592318 390698 592500 390934
rect -8576 390676 592500 390698
rect -8576 390674 -7976 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 137604 390674 138204 390676
rect 173604 390674 174204 390676
rect 281604 390674 282204 390676
rect 317604 390674 318204 390676
rect 353604 390674 354204 390676
rect 389604 390674 390204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591900 390674 592500 390676
rect -6696 387676 -6096 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 134004 387676 134604 387678
rect 170004 387676 170604 387678
rect 278004 387676 278604 387678
rect 314004 387676 314604 387678
rect 350004 387676 350604 387678
rect 386004 387676 386604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 590020 387676 590620 387678
rect -6696 387654 590620 387676
rect -6696 387418 -6514 387654
rect -6278 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 134186 387654
rect 134422 387418 170186 387654
rect 170422 387418 278186 387654
rect 278422 387418 314186 387654
rect 314422 387418 350186 387654
rect 350422 387418 386186 387654
rect 386422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590202 387654
rect 590438 387418 590620 387654
rect -6696 387334 590620 387418
rect -6696 387098 -6514 387334
rect -6278 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 134186 387334
rect 134422 387098 170186 387334
rect 170422 387098 278186 387334
rect 278422 387098 314186 387334
rect 314422 387098 350186 387334
rect 350422 387098 386186 387334
rect 386422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590202 387334
rect 590438 387098 590620 387334
rect -6696 387076 590620 387098
rect -6696 387074 -6096 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 134004 387074 134604 387076
rect 170004 387074 170604 387076
rect 278004 387074 278604 387076
rect 314004 387074 314604 387076
rect 350004 387074 350604 387076
rect 386004 387074 386604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 590020 387074 590620 387076
rect -4816 384076 -4216 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 130404 384076 131004 384078
rect 166404 384076 167004 384078
rect 274404 384076 275004 384078
rect 310404 384076 311004 384078
rect 346404 384076 347004 384078
rect 382404 384076 383004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588140 384076 588740 384078
rect -4816 384054 588740 384076
rect -4816 383818 -4634 384054
rect -4398 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 130586 384054
rect 130822 383818 166586 384054
rect 166822 383818 274586 384054
rect 274822 383818 310586 384054
rect 310822 383818 346586 384054
rect 346822 383818 382586 384054
rect 382822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588322 384054
rect 588558 383818 588740 384054
rect -4816 383734 588740 383818
rect -4816 383498 -4634 383734
rect -4398 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 130586 383734
rect 130822 383498 166586 383734
rect 166822 383498 274586 383734
rect 274822 383498 310586 383734
rect 310822 383498 346586 383734
rect 346822 383498 382586 383734
rect 382822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588322 383734
rect 588558 383498 588740 383734
rect -4816 383476 588740 383498
rect -4816 383474 -4216 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 130404 383474 131004 383476
rect 166404 383474 167004 383476
rect 274404 383474 275004 383476
rect 310404 383474 311004 383476
rect 346404 383474 347004 383476
rect 382404 383474 383004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588140 383474 588740 383476
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 91568 380476 91888 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 219568 380476 219888 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 394604 380476 394924 380478
rect 450804 380476 451404 380478
rect 479568 380476 479888 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 91610 380454
rect 91846 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 219610 380454
rect 219846 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 394646 380454
rect 394882 380218 450986 380454
rect 451222 380218 479610 380454
rect 479846 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 91610 380134
rect 91846 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 219610 380134
rect 219846 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 394646 380134
rect 394882 379898 450986 380134
rect 451222 379898 479610 380134
rect 479846 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 91568 379874 91888 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 219568 379874 219888 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 394604 379874 394924 379876
rect 450804 379874 451404 379876
rect 479568 379874 479888 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -7636 373276 -7036 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 155604 373276 156204 373278
rect 191604 373276 192204 373278
rect 299604 373276 300204 373278
rect 335604 373276 336204 373278
rect 371604 373276 372204 373278
rect 443604 373276 444204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590960 373276 591560 373278
rect -8576 373254 592500 373276
rect -8576 373018 -7454 373254
rect -7218 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 155786 373254
rect 156022 373018 191786 373254
rect 192022 373018 299786 373254
rect 300022 373018 335786 373254
rect 336022 373018 371786 373254
rect 372022 373018 443786 373254
rect 444022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591142 373254
rect 591378 373018 592500 373254
rect -8576 372934 592500 373018
rect -8576 372698 -7454 372934
rect -7218 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 155786 372934
rect 156022 372698 191786 372934
rect 192022 372698 299786 372934
rect 300022 372698 335786 372934
rect 336022 372698 371786 372934
rect 372022 372698 443786 372934
rect 444022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591142 372934
rect 591378 372698 592500 372934
rect -8576 372676 592500 372698
rect -7636 372674 -7036 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 155604 372674 156204 372676
rect 191604 372674 192204 372676
rect 299604 372674 300204 372676
rect 335604 372674 336204 372676
rect 371604 372674 372204 372676
rect 443604 372674 444204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590960 372674 591560 372676
rect -5756 369676 -5156 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 152004 369676 152604 369678
rect 188004 369676 188604 369678
rect 296004 369676 296604 369678
rect 332004 369676 332604 369678
rect 368004 369676 368604 369678
rect 440004 369676 440604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589080 369676 589680 369678
rect -6696 369654 590620 369676
rect -6696 369418 -5574 369654
rect -5338 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 152186 369654
rect 152422 369418 188186 369654
rect 188422 369418 296186 369654
rect 296422 369418 332186 369654
rect 332422 369418 368186 369654
rect 368422 369418 440186 369654
rect 440422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589262 369654
rect 589498 369418 590620 369654
rect -6696 369334 590620 369418
rect -6696 369098 -5574 369334
rect -5338 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 152186 369334
rect 152422 369098 188186 369334
rect 188422 369098 296186 369334
rect 296422 369098 332186 369334
rect 332422 369098 368186 369334
rect 368422 369098 440186 369334
rect 440422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589262 369334
rect 589498 369098 590620 369334
rect -6696 369076 590620 369098
rect -5756 369074 -5156 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 152004 369074 152604 369076
rect 188004 369074 188604 369076
rect 296004 369074 296604 369076
rect 332004 369074 332604 369076
rect 368004 369074 368604 369076
rect 440004 369074 440604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589080 369074 589680 369076
rect -3876 366076 -3276 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 148404 366076 149004 366078
rect 184404 366076 185004 366078
rect 292404 366076 293004 366078
rect 328404 366076 329004 366078
rect 364404 366076 365004 366078
rect 436404 366076 437004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587200 366076 587800 366078
rect -4816 366054 588740 366076
rect -4816 365818 -3694 366054
rect -3458 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 148586 366054
rect 148822 365818 184586 366054
rect 184822 365818 292586 366054
rect 292822 365818 328586 366054
rect 328822 365818 364586 366054
rect 364822 365818 436586 366054
rect 436822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587382 366054
rect 587618 365818 588740 366054
rect -4816 365734 588740 365818
rect -4816 365498 -3694 365734
rect -3458 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 148586 365734
rect 148822 365498 184586 365734
rect 184822 365498 292586 365734
rect 292822 365498 328586 365734
rect 328822 365498 364586 365734
rect 364822 365498 436586 365734
rect 436822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587382 365734
rect 587618 365498 588740 365734
rect -4816 365476 588740 365498
rect -3876 365474 -3276 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 148404 365474 149004 365476
rect 184404 365474 185004 365476
rect 292404 365474 293004 365476
rect 328404 365474 329004 365476
rect 364404 365474 365004 365476
rect 436404 365474 437004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587200 365474 587800 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 76208 362476 76528 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 204208 362476 204528 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 389774 362476 390094 362478
rect 432804 362476 433404 362478
rect 464208 362476 464528 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 76250 362454
rect 76486 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 204250 362454
rect 204486 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 389816 362454
rect 390052 362218 432986 362454
rect 433222 362218 464250 362454
rect 464486 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 76250 362134
rect 76486 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 204250 362134
rect 204486 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 389816 362134
rect 390052 361898 432986 362134
rect 433222 361898 464250 362134
rect 464486 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 76208 361874 76528 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 204208 361874 204528 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 389774 361874 390094 361876
rect 432804 361874 433404 361876
rect 464208 361874 464528 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8576 355276 -7976 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 137604 355276 138204 355278
rect 173604 355276 174204 355278
rect 281604 355276 282204 355278
rect 317604 355276 318204 355278
rect 353604 355276 354204 355278
rect 425604 355276 426204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591900 355276 592500 355278
rect -8576 355254 592500 355276
rect -8576 355018 -8394 355254
rect -8158 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 137786 355254
rect 138022 355018 173786 355254
rect 174022 355018 281786 355254
rect 282022 355018 317786 355254
rect 318022 355018 353786 355254
rect 354022 355018 425786 355254
rect 426022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 592082 355254
rect 592318 355018 592500 355254
rect -8576 354934 592500 355018
rect -8576 354698 -8394 354934
rect -8158 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 137786 354934
rect 138022 354698 173786 354934
rect 174022 354698 281786 354934
rect 282022 354698 317786 354934
rect 318022 354698 353786 354934
rect 354022 354698 425786 354934
rect 426022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 592082 354934
rect 592318 354698 592500 354934
rect -8576 354676 592500 354698
rect -8576 354674 -7976 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 137604 354674 138204 354676
rect 173604 354674 174204 354676
rect 281604 354674 282204 354676
rect 317604 354674 318204 354676
rect 353604 354674 354204 354676
rect 425604 354674 426204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591900 354674 592500 354676
rect -6696 351676 -6096 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 134004 351676 134604 351678
rect 170004 351676 170604 351678
rect 278004 351676 278604 351678
rect 314004 351676 314604 351678
rect 350004 351676 350604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 590020 351676 590620 351678
rect -6696 351654 590620 351676
rect -6696 351418 -6514 351654
rect -6278 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 134186 351654
rect 134422 351418 170186 351654
rect 170422 351418 278186 351654
rect 278422 351418 314186 351654
rect 314422 351418 350186 351654
rect 350422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590202 351654
rect 590438 351418 590620 351654
rect -6696 351334 590620 351418
rect -6696 351098 -6514 351334
rect -6278 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 134186 351334
rect 134422 351098 170186 351334
rect 170422 351098 278186 351334
rect 278422 351098 314186 351334
rect 314422 351098 350186 351334
rect 350422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590202 351334
rect 590438 351098 590620 351334
rect -6696 351076 590620 351098
rect -6696 351074 -6096 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 134004 351074 134604 351076
rect 170004 351074 170604 351076
rect 278004 351074 278604 351076
rect 314004 351074 314604 351076
rect 350004 351074 350604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 590020 351074 590620 351076
rect -4816 348076 -4216 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 130404 348076 131004 348078
rect 166404 348076 167004 348078
rect 274404 348076 275004 348078
rect 310404 348076 311004 348078
rect 346404 348076 347004 348078
rect 382404 348076 383004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588140 348076 588740 348078
rect -4816 348054 588740 348076
rect -4816 347818 -4634 348054
rect -4398 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 130586 348054
rect 130822 347818 166586 348054
rect 166822 347818 274586 348054
rect 274822 347818 310586 348054
rect 310822 347818 346586 348054
rect 346822 347818 382586 348054
rect 382822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588322 348054
rect 588558 347818 588740 348054
rect -4816 347734 588740 347818
rect -4816 347498 -4634 347734
rect -4398 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 130586 347734
rect 130822 347498 166586 347734
rect 166822 347498 274586 347734
rect 274822 347498 310586 347734
rect 310822 347498 346586 347734
rect 346822 347498 382586 347734
rect 382822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588322 347734
rect 588558 347498 588740 347734
rect -4816 347476 588740 347498
rect -4816 347474 -4216 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 130404 347474 131004 347476
rect 166404 347474 167004 347476
rect 274404 347474 275004 347476
rect 310404 347474 311004 347476
rect 346404 347474 347004 347476
rect 382404 347474 383004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588140 347474 588740 347476
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 91568 344476 91888 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 219568 344476 219888 344478
rect 270804 344476 271404 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 479568 344476 479888 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 91610 344454
rect 91846 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 219610 344454
rect 219846 344218 270986 344454
rect 271222 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 479610 344454
rect 479846 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 91610 344134
rect 91846 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 219610 344134
rect 219846 343898 270986 344134
rect 271222 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 479610 344134
rect 479846 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 91568 343874 91888 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 219568 343874 219888 343876
rect 270804 343874 271404 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 479568 343874 479888 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -7636 337276 -7036 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 155604 337276 156204 337278
rect 191604 337276 192204 337278
rect 227604 337276 228204 337278
rect 263604 337276 264204 337278
rect 299604 337276 300204 337278
rect 335604 337276 336204 337278
rect 371604 337276 372204 337278
rect 407604 337276 408204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590960 337276 591560 337278
rect -8576 337254 592500 337276
rect -8576 337018 -7454 337254
rect -7218 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 155786 337254
rect 156022 337018 191786 337254
rect 192022 337018 227786 337254
rect 228022 337018 263786 337254
rect 264022 337018 299786 337254
rect 300022 337018 335786 337254
rect 336022 337018 371786 337254
rect 372022 337018 407786 337254
rect 408022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591142 337254
rect 591378 337018 592500 337254
rect -8576 336934 592500 337018
rect -8576 336698 -7454 336934
rect -7218 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 155786 336934
rect 156022 336698 191786 336934
rect 192022 336698 227786 336934
rect 228022 336698 263786 336934
rect 264022 336698 299786 336934
rect 300022 336698 335786 336934
rect 336022 336698 371786 336934
rect 372022 336698 407786 336934
rect 408022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591142 336934
rect 591378 336698 592500 336934
rect -8576 336676 592500 336698
rect -7636 336674 -7036 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 155604 336674 156204 336676
rect 191604 336674 192204 336676
rect 227604 336674 228204 336676
rect 263604 336674 264204 336676
rect 299604 336674 300204 336676
rect 335604 336674 336204 336676
rect 371604 336674 372204 336676
rect 407604 336674 408204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590960 336674 591560 336676
rect -5756 333676 -5156 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 188004 333676 188604 333678
rect 224004 333676 224604 333678
rect 260004 333676 260604 333678
rect 296004 333676 296604 333678
rect 332004 333676 332604 333678
rect 368004 333676 368604 333678
rect 404004 333676 404604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589080 333676 589680 333678
rect -6696 333654 590620 333676
rect -6696 333418 -5574 333654
rect -5338 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 188186 333654
rect 188422 333418 224186 333654
rect 224422 333418 260186 333654
rect 260422 333418 296186 333654
rect 296422 333418 332186 333654
rect 332422 333418 368186 333654
rect 368422 333418 404186 333654
rect 404422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589262 333654
rect 589498 333418 590620 333654
rect -6696 333334 590620 333418
rect -6696 333098 -5574 333334
rect -5338 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 188186 333334
rect 188422 333098 224186 333334
rect 224422 333098 260186 333334
rect 260422 333098 296186 333334
rect 296422 333098 332186 333334
rect 332422 333098 368186 333334
rect 368422 333098 404186 333334
rect 404422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589262 333334
rect 589498 333098 590620 333334
rect -6696 333076 590620 333098
rect -5756 333074 -5156 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 188004 333074 188604 333076
rect 224004 333074 224604 333076
rect 260004 333074 260604 333076
rect 296004 333074 296604 333076
rect 332004 333074 332604 333076
rect 368004 333074 368604 333076
rect 404004 333074 404604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589080 333074 589680 333076
rect -3876 330076 -3276 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 184404 330076 185004 330078
rect 220404 330076 221004 330078
rect 256404 330076 257004 330078
rect 292404 330076 293004 330078
rect 328404 330076 329004 330078
rect 364404 330076 365004 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587200 330076 587800 330078
rect -4816 330054 588740 330076
rect -4816 329818 -3694 330054
rect -3458 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 184586 330054
rect 184822 329818 220586 330054
rect 220822 329818 256586 330054
rect 256822 329818 292586 330054
rect 292822 329818 328586 330054
rect 328822 329818 364586 330054
rect 364822 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587382 330054
rect 587618 329818 588740 330054
rect -4816 329734 588740 329818
rect -4816 329498 -3694 329734
rect -3458 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 184586 329734
rect 184822 329498 220586 329734
rect 220822 329498 256586 329734
rect 256822 329498 292586 329734
rect 292822 329498 328586 329734
rect 328822 329498 364586 329734
rect 364822 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587382 329734
rect 587618 329498 588740 329734
rect -4816 329476 588740 329498
rect -3876 329474 -3276 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 184404 329474 185004 329476
rect 220404 329474 221004 329476
rect 256404 329474 257004 329476
rect 292404 329474 293004 329476
rect 328404 329474 329004 329476
rect 364404 329474 365004 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587200 329474 587800 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8576 319276 -7976 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 173604 319276 174204 319278
rect 209604 319276 210204 319278
rect 245604 319276 246204 319278
rect 281604 319276 282204 319278
rect 317604 319276 318204 319278
rect 353604 319276 354204 319278
rect 389604 319276 390204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591900 319276 592500 319278
rect -8576 319254 592500 319276
rect -8576 319018 -8394 319254
rect -8158 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 173786 319254
rect 174022 319018 209786 319254
rect 210022 319018 245786 319254
rect 246022 319018 281786 319254
rect 282022 319018 317786 319254
rect 318022 319018 353786 319254
rect 354022 319018 389786 319254
rect 390022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 592082 319254
rect 592318 319018 592500 319254
rect -8576 318934 592500 319018
rect -8576 318698 -8394 318934
rect -8158 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 173786 318934
rect 174022 318698 209786 318934
rect 210022 318698 245786 318934
rect 246022 318698 281786 318934
rect 282022 318698 317786 318934
rect 318022 318698 353786 318934
rect 354022 318698 389786 318934
rect 390022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 592082 318934
rect 592318 318698 592500 318934
rect -8576 318676 592500 318698
rect -8576 318674 -7976 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 173604 318674 174204 318676
rect 209604 318674 210204 318676
rect 245604 318674 246204 318676
rect 281604 318674 282204 318676
rect 317604 318674 318204 318676
rect 353604 318674 354204 318676
rect 389604 318674 390204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591900 318674 592500 318676
rect -6696 315676 -6096 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 590020 315676 590620 315678
rect -6696 315654 590620 315676
rect -6696 315418 -6514 315654
rect -6278 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590202 315654
rect 590438 315418 590620 315654
rect -6696 315334 590620 315418
rect -6696 315098 -6514 315334
rect -6278 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590202 315334
rect 590438 315098 590620 315334
rect -6696 315076 590620 315098
rect -6696 315074 -6096 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 590020 315074 590620 315076
rect -4816 312076 -4216 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588140 312076 588740 312078
rect -4816 312054 588740 312076
rect -4816 311818 -4634 312054
rect -4398 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588322 312054
rect 588558 311818 588740 312054
rect -4816 311734 588740 311818
rect -4816 311498 -4634 311734
rect -4398 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588322 311734
rect 588558 311498 588740 311734
rect -4816 311476 588740 311498
rect -4816 311474 -4216 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588140 311474 588740 311476
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -7636 301276 -7036 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590960 301276 591560 301278
rect -8576 301254 592500 301276
rect -8576 301018 -7454 301254
rect -7218 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591142 301254
rect 591378 301018 592500 301254
rect -8576 300934 592500 301018
rect -8576 300698 -7454 300934
rect -7218 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591142 300934
rect 591378 300698 592500 300934
rect -8576 300676 592500 300698
rect -7636 300674 -7036 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590960 300674 591560 300676
rect -5756 297676 -5156 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589080 297676 589680 297678
rect -6696 297654 590620 297676
rect -6696 297418 -5574 297654
rect -5338 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589262 297654
rect 589498 297418 590620 297654
rect -6696 297334 590620 297418
rect -6696 297098 -5574 297334
rect -5338 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589262 297334
rect 589498 297098 590620 297334
rect -6696 297076 590620 297098
rect -5756 297074 -5156 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589080 297074 589680 297076
rect -3876 294076 -3276 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587200 294076 587800 294078
rect -4816 294054 588740 294076
rect -4816 293818 -3694 294054
rect -3458 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587382 294054
rect 587618 293818 588740 294054
rect -4816 293734 588740 293818
rect -4816 293498 -3694 293734
rect -3458 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587382 293734
rect 587618 293498 588740 293734
rect -4816 293476 588740 293498
rect -3876 293474 -3276 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587200 293474 587800 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8576 283276 -7976 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591900 283276 592500 283278
rect -8576 283254 592500 283276
rect -8576 283018 -8394 283254
rect -8158 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 592082 283254
rect 592318 283018 592500 283254
rect -8576 282934 592500 283018
rect -8576 282698 -8394 282934
rect -8158 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 592082 282934
rect 592318 282698 592500 282934
rect -8576 282676 592500 282698
rect -8576 282674 -7976 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591900 282674 592500 282676
rect -6696 279676 -6096 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 590020 279676 590620 279678
rect -6696 279654 590620 279676
rect -6696 279418 -6514 279654
rect -6278 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590202 279654
rect 590438 279418 590620 279654
rect -6696 279334 590620 279418
rect -6696 279098 -6514 279334
rect -6278 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590202 279334
rect 590438 279098 590620 279334
rect -6696 279076 590620 279098
rect -6696 279074 -6096 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 590020 279074 590620 279076
rect -4816 276076 -4216 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588140 276076 588740 276078
rect -4816 276054 588740 276076
rect -4816 275818 -4634 276054
rect -4398 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588322 276054
rect 588558 275818 588740 276054
rect -4816 275734 588740 275818
rect -4816 275498 -4634 275734
rect -4398 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588322 275734
rect 588558 275498 588740 275734
rect -4816 275476 588740 275498
rect -4816 275474 -4216 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588140 275474 588740 275476
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -7636 265276 -7036 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590960 265276 591560 265278
rect -8576 265254 592500 265276
rect -8576 265018 -7454 265254
rect -7218 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591142 265254
rect 591378 265018 592500 265254
rect -8576 264934 592500 265018
rect -8576 264698 -7454 264934
rect -7218 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591142 264934
rect 591378 264698 592500 264934
rect -8576 264676 592500 264698
rect -7636 264674 -7036 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590960 264674 591560 264676
rect -5756 261676 -5156 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589080 261676 589680 261678
rect -6696 261654 590620 261676
rect -6696 261418 -5574 261654
rect -5338 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589262 261654
rect 589498 261418 590620 261654
rect -6696 261334 590620 261418
rect -6696 261098 -5574 261334
rect -5338 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589262 261334
rect 589498 261098 590620 261334
rect -6696 261076 590620 261098
rect -5756 261074 -5156 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589080 261074 589680 261076
rect -3876 258076 -3276 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587200 258076 587800 258078
rect -4816 258054 588740 258076
rect -4816 257818 -3694 258054
rect -3458 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587382 258054
rect 587618 257818 588740 258054
rect -4816 257734 588740 257818
rect -4816 257498 -3694 257734
rect -3458 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587382 257734
rect 587618 257498 588740 257734
rect -4816 257476 588740 257498
rect -3876 257474 -3276 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587200 257474 587800 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8576 247276 -7976 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591900 247276 592500 247278
rect -8576 247254 592500 247276
rect -8576 247018 -8394 247254
rect -8158 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 592082 247254
rect 592318 247018 592500 247254
rect -8576 246934 592500 247018
rect -8576 246698 -8394 246934
rect -8158 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 592082 246934
rect 592318 246698 592500 246934
rect -8576 246676 592500 246698
rect -8576 246674 -7976 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591900 246674 592500 246676
rect -6696 243676 -6096 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 590020 243676 590620 243678
rect -6696 243654 590620 243676
rect -6696 243418 -6514 243654
rect -6278 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590202 243654
rect 590438 243418 590620 243654
rect -6696 243334 590620 243418
rect -6696 243098 -6514 243334
rect -6278 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590202 243334
rect 590438 243098 590620 243334
rect -6696 243076 590620 243098
rect -6696 243074 -6096 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 590020 243074 590620 243076
rect -4816 240076 -4216 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588140 240076 588740 240078
rect -4816 240054 588740 240076
rect -4816 239818 -4634 240054
rect -4398 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588322 240054
rect 588558 239818 588740 240054
rect -4816 239734 588740 239818
rect -4816 239498 -4634 239734
rect -4398 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588322 239734
rect 588558 239498 588740 239734
rect -4816 239476 588740 239498
rect -4816 239474 -4216 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588140 239474 588740 239476
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -7636 229276 -7036 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590960 229276 591560 229278
rect -8576 229254 592500 229276
rect -8576 229018 -7454 229254
rect -7218 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591142 229254
rect 591378 229018 592500 229254
rect -8576 228934 592500 229018
rect -8576 228698 -7454 228934
rect -7218 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591142 228934
rect 591378 228698 592500 228934
rect -8576 228676 592500 228698
rect -7636 228674 -7036 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590960 228674 591560 228676
rect -5756 225676 -5156 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589080 225676 589680 225678
rect -6696 225654 590620 225676
rect -6696 225418 -5574 225654
rect -5338 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589262 225654
rect 589498 225418 590620 225654
rect -6696 225334 590620 225418
rect -6696 225098 -5574 225334
rect -5338 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589262 225334
rect 589498 225098 590620 225334
rect -6696 225076 590620 225098
rect -5756 225074 -5156 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589080 225074 589680 225076
rect -3876 222076 -3276 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587200 222076 587800 222078
rect -4816 222054 588740 222076
rect -4816 221818 -3694 222054
rect -3458 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587382 222054
rect 587618 221818 588740 222054
rect -4816 221734 588740 221818
rect -4816 221498 -3694 221734
rect -3458 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587382 221734
rect 587618 221498 588740 221734
rect -4816 221476 588740 221498
rect -3876 221474 -3276 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587200 221474 587800 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8576 211276 -7976 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591900 211276 592500 211278
rect -8576 211254 592500 211276
rect -8576 211018 -8394 211254
rect -8158 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 592082 211254
rect 592318 211018 592500 211254
rect -8576 210934 592500 211018
rect -8576 210698 -8394 210934
rect -8158 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 592082 210934
rect 592318 210698 592500 210934
rect -8576 210676 592500 210698
rect -8576 210674 -7976 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591900 210674 592500 210676
rect -6696 207676 -6096 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 590020 207676 590620 207678
rect -6696 207654 590620 207676
rect -6696 207418 -6514 207654
rect -6278 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590202 207654
rect 590438 207418 590620 207654
rect -6696 207334 590620 207418
rect -6696 207098 -6514 207334
rect -6278 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590202 207334
rect 590438 207098 590620 207334
rect -6696 207076 590620 207098
rect -6696 207074 -6096 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 590020 207074 590620 207076
rect -4816 204076 -4216 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588140 204076 588740 204078
rect -4816 204054 588740 204076
rect -4816 203818 -4634 204054
rect -4398 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588322 204054
rect 588558 203818 588740 204054
rect -4816 203734 588740 203818
rect -4816 203498 -4634 203734
rect -4398 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588322 203734
rect 588558 203498 588740 203734
rect -4816 203476 588740 203498
rect -4816 203474 -4216 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588140 203474 588740 203476
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -7636 193276 -7036 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590960 193276 591560 193278
rect -8576 193254 592500 193276
rect -8576 193018 -7454 193254
rect -7218 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591142 193254
rect 591378 193018 592500 193254
rect -8576 192934 592500 193018
rect -8576 192698 -7454 192934
rect -7218 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591142 192934
rect 591378 192698 592500 192934
rect -8576 192676 592500 192698
rect -7636 192674 -7036 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590960 192674 591560 192676
rect -5756 189676 -5156 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589080 189676 589680 189678
rect -6696 189654 590620 189676
rect -6696 189418 -5574 189654
rect -5338 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589262 189654
rect 589498 189418 590620 189654
rect -6696 189334 590620 189418
rect -6696 189098 -5574 189334
rect -5338 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589262 189334
rect 589498 189098 590620 189334
rect -6696 189076 590620 189098
rect -5756 189074 -5156 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589080 189074 589680 189076
rect -3876 186076 -3276 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587200 186076 587800 186078
rect -4816 186054 588740 186076
rect -4816 185818 -3694 186054
rect -3458 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587382 186054
rect 587618 185818 588740 186054
rect -4816 185734 588740 185818
rect -4816 185498 -3694 185734
rect -3458 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587382 185734
rect 587618 185498 588740 185734
rect -4816 185476 588740 185498
rect -3876 185474 -3276 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587200 185474 587800 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 138208 182476 138528 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 138250 182454
rect 138486 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 138250 182134
rect 138486 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 138208 181874 138528 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8576 175276 -7976 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591900 175276 592500 175278
rect -8576 175254 592500 175276
rect -8576 175018 -8394 175254
rect -8158 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 592082 175254
rect 592318 175018 592500 175254
rect -8576 174934 592500 175018
rect -8576 174698 -8394 174934
rect -8158 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 592082 174934
rect 592318 174698 592500 174934
rect -8576 174676 592500 174698
rect -8576 174674 -7976 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591900 174674 592500 174676
rect -6696 171676 -6096 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 590020 171676 590620 171678
rect -6696 171654 590620 171676
rect -6696 171418 -6514 171654
rect -6278 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590202 171654
rect 590438 171418 590620 171654
rect -6696 171334 590620 171418
rect -6696 171098 -6514 171334
rect -6278 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590202 171334
rect 590438 171098 590620 171334
rect -6696 171076 590620 171098
rect -6696 171074 -6096 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 590020 171074 590620 171076
rect -4816 168076 -4216 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588140 168076 588740 168078
rect -4816 168054 588740 168076
rect -4816 167818 -4634 168054
rect -4398 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588322 168054
rect 588558 167818 588740 168054
rect -4816 167734 588740 167818
rect -4816 167498 -4634 167734
rect -4398 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588322 167734
rect 588558 167498 588740 167734
rect -4816 167476 588740 167498
rect -4816 167474 -4216 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588140 167474 588740 167476
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 153568 164476 153888 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 153610 164454
rect 153846 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 153610 164134
rect 153846 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 153568 163874 153888 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -7636 157276 -7036 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590960 157276 591560 157278
rect -8576 157254 592500 157276
rect -8576 157018 -7454 157254
rect -7218 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591142 157254
rect 591378 157018 592500 157254
rect -8576 156934 592500 157018
rect -8576 156698 -7454 156934
rect -7218 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591142 156934
rect 591378 156698 592500 156934
rect -8576 156676 592500 156698
rect -7636 156674 -7036 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590960 156674 591560 156676
rect -5756 153676 -5156 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589080 153676 589680 153678
rect -6696 153654 590620 153676
rect -6696 153418 -5574 153654
rect -5338 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589262 153654
rect 589498 153418 590620 153654
rect -6696 153334 590620 153418
rect -6696 153098 -5574 153334
rect -5338 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589262 153334
rect 589498 153098 590620 153334
rect -6696 153076 590620 153098
rect -5756 153074 -5156 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589080 153074 589680 153076
rect -3876 150076 -3276 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587200 150076 587800 150078
rect -4816 150054 588740 150076
rect -4816 149818 -3694 150054
rect -3458 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587382 150054
rect 587618 149818 588740 150054
rect -4816 149734 588740 149818
rect -4816 149498 -3694 149734
rect -3458 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587382 149734
rect 587618 149498 588740 149734
rect -4816 149476 588740 149498
rect -3876 149474 -3276 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587200 149474 587800 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 138208 146476 138528 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 138250 146454
rect 138486 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 138250 146134
rect 138486 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 138208 145874 138528 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8576 139276 -7976 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591900 139276 592500 139278
rect -8576 139254 592500 139276
rect -8576 139018 -8394 139254
rect -8158 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 592082 139254
rect 592318 139018 592500 139254
rect -8576 138934 592500 139018
rect -8576 138698 -8394 138934
rect -8158 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 592082 138934
rect 592318 138698 592500 138934
rect -8576 138676 592500 138698
rect -8576 138674 -7976 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591900 138674 592500 138676
rect -6696 135676 -6096 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 590020 135676 590620 135678
rect -6696 135654 590620 135676
rect -6696 135418 -6514 135654
rect -6278 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590202 135654
rect 590438 135418 590620 135654
rect -6696 135334 590620 135418
rect -6696 135098 -6514 135334
rect -6278 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590202 135334
rect 590438 135098 590620 135334
rect -6696 135076 590620 135098
rect -6696 135074 -6096 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 590020 135074 590620 135076
rect -4816 132076 -4216 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588140 132076 588740 132078
rect -4816 132054 588740 132076
rect -4816 131818 -4634 132054
rect -4398 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588322 132054
rect 588558 131818 588740 132054
rect -4816 131734 588740 131818
rect -4816 131498 -4634 131734
rect -4398 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588322 131734
rect 588558 131498 588740 131734
rect -4816 131476 588740 131498
rect -4816 131474 -4216 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588140 131474 588740 131476
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 153568 128476 153888 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 153610 128454
rect 153846 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 153610 128134
rect 153846 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 153568 127874 153888 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -7636 121276 -7036 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590960 121276 591560 121278
rect -8576 121254 592500 121276
rect -8576 121018 -7454 121254
rect -7218 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591142 121254
rect 591378 121018 592500 121254
rect -8576 120934 592500 121018
rect -8576 120698 -7454 120934
rect -7218 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591142 120934
rect 591378 120698 592500 120934
rect -8576 120676 592500 120698
rect -7636 120674 -7036 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590960 120674 591560 120676
rect -5756 117676 -5156 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589080 117676 589680 117678
rect -6696 117654 590620 117676
rect -6696 117418 -5574 117654
rect -5338 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589262 117654
rect 589498 117418 590620 117654
rect -6696 117334 590620 117418
rect -6696 117098 -5574 117334
rect -5338 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589262 117334
rect 589498 117098 590620 117334
rect -6696 117076 590620 117098
rect -5756 117074 -5156 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589080 117074 589680 117076
rect -3876 114076 -3276 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587200 114076 587800 114078
rect -4816 114054 588740 114076
rect -4816 113818 -3694 114054
rect -3458 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587382 114054
rect 587618 113818 588740 114054
rect -4816 113734 588740 113818
rect -4816 113498 -3694 113734
rect -3458 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587382 113734
rect 587618 113498 588740 113734
rect -4816 113476 588740 113498
rect -3876 113474 -3276 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587200 113474 587800 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8576 103276 -7976 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591900 103276 592500 103278
rect -8576 103254 592500 103276
rect -8576 103018 -8394 103254
rect -8158 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 592082 103254
rect 592318 103018 592500 103254
rect -8576 102934 592500 103018
rect -8576 102698 -8394 102934
rect -8158 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 592082 102934
rect 592318 102698 592500 102934
rect -8576 102676 592500 102698
rect -8576 102674 -7976 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591900 102674 592500 102676
rect -6696 99676 -6096 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 590020 99676 590620 99678
rect -6696 99654 590620 99676
rect -6696 99418 -6514 99654
rect -6278 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590202 99654
rect 590438 99418 590620 99654
rect -6696 99334 590620 99418
rect -6696 99098 -6514 99334
rect -6278 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590202 99334
rect 590438 99098 590620 99334
rect -6696 99076 590620 99098
rect -6696 99074 -6096 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 590020 99074 590620 99076
rect -4816 96076 -4216 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588140 96076 588740 96078
rect -4816 96054 588740 96076
rect -4816 95818 -4634 96054
rect -4398 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588322 96054
rect 588558 95818 588740 96054
rect -4816 95734 588740 95818
rect -4816 95498 -4634 95734
rect -4398 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588322 95734
rect 588558 95498 588740 95734
rect -4816 95476 588740 95498
rect -4816 95474 -4216 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588140 95474 588740 95476
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -7636 85276 -7036 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590960 85276 591560 85278
rect -8576 85254 592500 85276
rect -8576 85018 -7454 85254
rect -7218 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591142 85254
rect 591378 85018 592500 85254
rect -8576 84934 592500 85018
rect -8576 84698 -7454 84934
rect -7218 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591142 84934
rect 591378 84698 592500 84934
rect -8576 84676 592500 84698
rect -7636 84674 -7036 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590960 84674 591560 84676
rect -5756 81676 -5156 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589080 81676 589680 81678
rect -6696 81654 590620 81676
rect -6696 81418 -5574 81654
rect -5338 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589262 81654
rect 589498 81418 590620 81654
rect -6696 81334 590620 81418
rect -6696 81098 -5574 81334
rect -5338 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589262 81334
rect 589498 81098 590620 81334
rect -6696 81076 590620 81098
rect -5756 81074 -5156 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589080 81074 589680 81076
rect -3876 78076 -3276 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587200 78076 587800 78078
rect -4816 78054 588740 78076
rect -4816 77818 -3694 78054
rect -3458 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587382 78054
rect 587618 77818 588740 78054
rect -4816 77734 588740 77818
rect -4816 77498 -3694 77734
rect -3458 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587382 77734
rect 587618 77498 588740 77734
rect -4816 77476 588740 77498
rect -3876 77474 -3276 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587200 77474 587800 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8576 67276 -7976 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591900 67276 592500 67278
rect -8576 67254 592500 67276
rect -8576 67018 -8394 67254
rect -8158 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 592082 67254
rect 592318 67018 592500 67254
rect -8576 66934 592500 67018
rect -8576 66698 -8394 66934
rect -8158 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 592082 66934
rect 592318 66698 592500 66934
rect -8576 66676 592500 66698
rect -8576 66674 -7976 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591900 66674 592500 66676
rect -6696 63676 -6096 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 590020 63676 590620 63678
rect -6696 63654 590620 63676
rect -6696 63418 -6514 63654
rect -6278 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590202 63654
rect 590438 63418 590620 63654
rect -6696 63334 590620 63418
rect -6696 63098 -6514 63334
rect -6278 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590202 63334
rect 590438 63098 590620 63334
rect -6696 63076 590620 63098
rect -6696 63074 -6096 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 590020 63074 590620 63076
rect -4816 60076 -4216 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588140 60076 588740 60078
rect -4816 60054 588740 60076
rect -4816 59818 -4634 60054
rect -4398 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588322 60054
rect 588558 59818 588740 60054
rect -4816 59734 588740 59818
rect -4816 59498 -4634 59734
rect -4398 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588322 59734
rect 588558 59498 588740 59734
rect -4816 59476 588740 59498
rect -4816 59474 -4216 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588140 59474 588740 59476
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -7636 49276 -7036 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590960 49276 591560 49278
rect -8576 49254 592500 49276
rect -8576 49018 -7454 49254
rect -7218 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591142 49254
rect 591378 49018 592500 49254
rect -8576 48934 592500 49018
rect -8576 48698 -7454 48934
rect -7218 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591142 48934
rect 591378 48698 592500 48934
rect -8576 48676 592500 48698
rect -7636 48674 -7036 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590960 48674 591560 48676
rect -5756 45676 -5156 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589080 45676 589680 45678
rect -6696 45654 590620 45676
rect -6696 45418 -5574 45654
rect -5338 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589262 45654
rect 589498 45418 590620 45654
rect -6696 45334 590620 45418
rect -6696 45098 -5574 45334
rect -5338 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589262 45334
rect 589498 45098 590620 45334
rect -6696 45076 590620 45098
rect -5756 45074 -5156 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589080 45074 589680 45076
rect -3876 42076 -3276 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587200 42076 587800 42078
rect -4816 42054 588740 42076
rect -4816 41818 -3694 42054
rect -3458 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587382 42054
rect 587618 41818 588740 42054
rect -4816 41734 588740 41818
rect -4816 41498 -3694 41734
rect -3458 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587382 41734
rect 587618 41498 588740 41734
rect -4816 41476 588740 41498
rect -3876 41474 -3276 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587200 41474 587800 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8576 31276 -7976 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591900 31276 592500 31278
rect -8576 31254 592500 31276
rect -8576 31018 -8394 31254
rect -8158 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 592082 31254
rect 592318 31018 592500 31254
rect -8576 30934 592500 31018
rect -8576 30698 -8394 30934
rect -8158 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 592082 30934
rect 592318 30698 592500 30934
rect -8576 30676 592500 30698
rect -8576 30674 -7976 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591900 30674 592500 30676
rect -6696 27676 -6096 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 590020 27676 590620 27678
rect -6696 27654 590620 27676
rect -6696 27418 -6514 27654
rect -6278 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590202 27654
rect 590438 27418 590620 27654
rect -6696 27334 590620 27418
rect -6696 27098 -6514 27334
rect -6278 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590202 27334
rect 590438 27098 590620 27334
rect -6696 27076 590620 27098
rect -6696 27074 -6096 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 590020 27074 590620 27076
rect -4816 24076 -4216 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588140 24076 588740 24078
rect -4816 24054 588740 24076
rect -4816 23818 -4634 24054
rect -4398 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588322 24054
rect 588558 23818 588740 24054
rect -4816 23734 588740 23818
rect -4816 23498 -4634 23734
rect -4398 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588322 23734
rect 588558 23498 588740 23734
rect -4816 23476 588740 23498
rect -4816 23474 -4216 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588140 23474 588740 23476
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -7636 13276 -7036 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590960 13276 591560 13278
rect -8576 13254 592500 13276
rect -8576 13018 -7454 13254
rect -7218 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591142 13254
rect 591378 13018 592500 13254
rect -8576 12934 592500 13018
rect -8576 12698 -7454 12934
rect -7218 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591142 12934
rect 591378 12698 592500 12934
rect -8576 12676 592500 12698
rect -7636 12674 -7036 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590960 12674 591560 12676
rect -5756 9676 -5156 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589080 9676 589680 9678
rect -6696 9654 590620 9676
rect -6696 9418 -5574 9654
rect -5338 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589262 9654
rect 589498 9418 590620 9654
rect -6696 9334 590620 9418
rect -6696 9098 -5574 9334
rect -5338 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589262 9334
rect 589498 9098 590620 9334
rect -6696 9076 590620 9098
rect -5756 9074 -5156 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589080 9074 589680 9076
rect -3876 6076 -3276 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587200 6076 587800 6078
rect -4816 6054 588740 6076
rect -4816 5818 -3694 6054
rect -3458 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587382 6054
rect 587618 5818 588740 6054
rect -4816 5734 588740 5818
rect -4816 5498 -3694 5734
rect -3458 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587382 5734
rect 587618 5498 588740 5734
rect -4816 5476 588740 5498
rect -3876 5474 -3276 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587200 5474 587800 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 4586 -2226
rect 4822 -2462 40586 -2226
rect 40822 -2462 76586 -2226
rect 76822 -2462 112586 -2226
rect 112822 -2462 148586 -2226
rect 148822 -2462 184586 -2226
rect 184822 -2462 220586 -2226
rect 220822 -2462 256586 -2226
rect 256822 -2462 292586 -2226
rect 292822 -2462 328586 -2226
rect 328822 -2462 364586 -2226
rect 364822 -2462 400586 -2226
rect 400822 -2462 436586 -2226
rect 436822 -2462 472586 -2226
rect 472822 -2462 508586 -2226
rect 508822 -2462 544586 -2226
rect 544822 -2462 580586 -2226
rect 580822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 4586 -2546
rect 4822 -2782 40586 -2546
rect 40822 -2782 76586 -2546
rect 76822 -2782 112586 -2546
rect 112822 -2782 148586 -2546
rect 148822 -2782 184586 -2546
rect 184822 -2782 220586 -2546
rect 220822 -2782 256586 -2546
rect 256822 -2782 292586 -2546
rect 292822 -2782 328586 -2546
rect 328822 -2782 364586 -2546
rect 364822 -2782 400586 -2546
rect 400822 -2782 436586 -2546
rect 436822 -2782 472586 -2546
rect 472822 -2782 508586 -2546
rect 508822 -2782 544586 -2546
rect 544822 -2782 580586 -2546
rect 580822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 22586 -3166
rect 22822 -3402 58586 -3166
rect 58822 -3402 94586 -3166
rect 94822 -3402 130586 -3166
rect 130822 -3402 166586 -3166
rect 166822 -3402 202586 -3166
rect 202822 -3402 238586 -3166
rect 238822 -3402 274586 -3166
rect 274822 -3402 310586 -3166
rect 310822 -3402 346586 -3166
rect 346822 -3402 382586 -3166
rect 382822 -3402 418586 -3166
rect 418822 -3402 454586 -3166
rect 454822 -3402 490586 -3166
rect 490822 -3402 526586 -3166
rect 526822 -3402 562586 -3166
rect 562822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 22586 -3486
rect 22822 -3722 58586 -3486
rect 58822 -3722 94586 -3486
rect 94822 -3722 130586 -3486
rect 130822 -3722 166586 -3486
rect 166822 -3722 202586 -3486
rect 202822 -3722 238586 -3486
rect 238822 -3722 274586 -3486
rect 274822 -3722 310586 -3486
rect 310822 -3722 346586 -3486
rect 346822 -3722 382586 -3486
rect 382822 -3722 418586 -3486
rect 418822 -3722 454586 -3486
rect 454822 -3722 490586 -3486
rect 490822 -3722 526586 -3486
rect 526822 -3722 562586 -3486
rect 562822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 8186 -4106
rect 8422 -4342 44186 -4106
rect 44422 -4342 80186 -4106
rect 80422 -4342 116186 -4106
rect 116422 -4342 152186 -4106
rect 152422 -4342 188186 -4106
rect 188422 -4342 224186 -4106
rect 224422 -4342 260186 -4106
rect 260422 -4342 296186 -4106
rect 296422 -4342 332186 -4106
rect 332422 -4342 368186 -4106
rect 368422 -4342 404186 -4106
rect 404422 -4342 440186 -4106
rect 440422 -4342 476186 -4106
rect 476422 -4342 512186 -4106
rect 512422 -4342 548186 -4106
rect 548422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 8186 -4426
rect 8422 -4662 44186 -4426
rect 44422 -4662 80186 -4426
rect 80422 -4662 116186 -4426
rect 116422 -4662 152186 -4426
rect 152422 -4662 188186 -4426
rect 188422 -4662 224186 -4426
rect 224422 -4662 260186 -4426
rect 260422 -4662 296186 -4426
rect 296422 -4662 332186 -4426
rect 332422 -4662 368186 -4426
rect 368422 -4662 404186 -4426
rect 404422 -4662 440186 -4426
rect 440422 -4662 476186 -4426
rect 476422 -4662 512186 -4426
rect 512422 -4662 548186 -4426
rect 548422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 26186 -5046
rect 26422 -5282 62186 -5046
rect 62422 -5282 98186 -5046
rect 98422 -5282 134186 -5046
rect 134422 -5282 170186 -5046
rect 170422 -5282 206186 -5046
rect 206422 -5282 242186 -5046
rect 242422 -5282 278186 -5046
rect 278422 -5282 314186 -5046
rect 314422 -5282 350186 -5046
rect 350422 -5282 386186 -5046
rect 386422 -5282 422186 -5046
rect 422422 -5282 458186 -5046
rect 458422 -5282 494186 -5046
rect 494422 -5282 530186 -5046
rect 530422 -5282 566186 -5046
rect 566422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 26186 -5366
rect 26422 -5602 62186 -5366
rect 62422 -5602 98186 -5366
rect 98422 -5602 134186 -5366
rect 134422 -5602 170186 -5366
rect 170422 -5602 206186 -5366
rect 206422 -5602 242186 -5366
rect 242422 -5602 278186 -5366
rect 278422 -5602 314186 -5366
rect 314422 -5602 350186 -5366
rect 350422 -5602 386186 -5366
rect 386422 -5602 422186 -5366
rect 422422 -5602 458186 -5366
rect 458422 -5602 494186 -5366
rect 494422 -5602 530186 -5366
rect 530422 -5602 566186 -5366
rect 566422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 11786 -5986
rect 12022 -6222 47786 -5986
rect 48022 -6222 83786 -5986
rect 84022 -6222 119786 -5986
rect 120022 -6222 155786 -5986
rect 156022 -6222 191786 -5986
rect 192022 -6222 227786 -5986
rect 228022 -6222 263786 -5986
rect 264022 -6222 299786 -5986
rect 300022 -6222 335786 -5986
rect 336022 -6222 371786 -5986
rect 372022 -6222 407786 -5986
rect 408022 -6222 443786 -5986
rect 444022 -6222 479786 -5986
rect 480022 -6222 515786 -5986
rect 516022 -6222 551786 -5986
rect 552022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 11786 -6306
rect 12022 -6542 47786 -6306
rect 48022 -6542 83786 -6306
rect 84022 -6542 119786 -6306
rect 120022 -6542 155786 -6306
rect 156022 -6542 191786 -6306
rect 192022 -6542 227786 -6306
rect 228022 -6542 263786 -6306
rect 264022 -6542 299786 -6306
rect 300022 -6542 335786 -6306
rect 336022 -6542 371786 -6306
rect 372022 -6542 407786 -6306
rect 408022 -6542 443786 -6306
rect 444022 -6542 479786 -6306
rect 480022 -6542 515786 -6306
rect 516022 -6542 551786 -6306
rect 552022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 29786 -6926
rect 30022 -7162 65786 -6926
rect 66022 -7162 101786 -6926
rect 102022 -7162 137786 -6926
rect 138022 -7162 173786 -6926
rect 174022 -7162 209786 -6926
rect 210022 -7162 245786 -6926
rect 246022 -7162 281786 -6926
rect 282022 -7162 317786 -6926
rect 318022 -7162 353786 -6926
rect 354022 -7162 389786 -6926
rect 390022 -7162 425786 -6926
rect 426022 -7162 461786 -6926
rect 462022 -7162 497786 -6926
rect 498022 -7162 533786 -6926
rect 534022 -7162 569786 -6926
rect 570022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 29786 -7246
rect 30022 -7482 65786 -7246
rect 66022 -7482 101786 -7246
rect 102022 -7482 137786 -7246
rect 138022 -7482 173786 -7246
rect 174022 -7482 209786 -7246
rect 210022 -7482 245786 -7246
rect 246022 -7482 281786 -7246
rect 282022 -7482 317786 -7246
rect 318022 -7482 353786 -7246
rect 354022 -7482 389786 -7246
rect 390022 -7482 425786 -7246
rect 426022 -7482 461786 -7246
rect 462022 -7482 497786 -7246
rect 498022 -7482 533786 -7246
rect 534022 -7482 569786 -7246
rect 570022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
use MM2hdmi  proj_7
timestamp 1608298212
transform 1 0 200000 0 1 520000
box 0 0 20000 40000
use challenge  proj_6
timestamp 1608298212
transform 1 0 480000 0 1 520000
box 0 0 31344 34764
use watch_hhmm  proj_5
timestamp 1608298212
transform 1 0 384000 0 1 350000
box 0 0 31275 33419
use asic_freq  proj_4
timestamp 1608298212
transform 1 0 300000 0 1 500000
box 0 0 77867 80011
use spinet5  proj_3
timestamp 1608298212
transform 1 0 200000 0 1 340000
box 0 0 66678 68822
use vga_clock  proj_2
timestamp 1608298212
transform 1 0 460000 0 1 340000
box 0 0 45405 47549
use ws2812  proj_1
timestamp 1608298212
transform 1 0 72000 0 1 340000
box 0 0 54206 56350
use seven_segment_seconds  proj_0
timestamp 1608298212
transform 1 0 86000 0 1 520000
box 0 0 29760 31904
use multi_project_harness  mprj
timestamp 1608298212
transform 1 0 134000 0 1 120000
box 0 0 300000 80000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
