magic
tech sky130A
magscale 1 2
timestamp 1608124775
<< locali >>
rect 153577 666587 153611 684437
rect 153485 647275 153519 656829
rect 142813 578527 142847 578765
rect 153393 569959 153427 579581
rect 154589 578731 154623 578833
rect 164157 578731 164191 578833
rect 176611 578765 176669 578799
rect 183569 578731 183603 578901
rect 193137 578799 193171 578901
rect 195931 578765 196115 578799
rect 196081 578731 196115 578765
rect 202889 578731 202923 578901
rect 212457 578799 212491 578901
rect 215251 578765 215435 578799
rect 215401 578731 215435 578765
rect 222209 578731 222243 578901
rect 231777 578799 231811 578901
rect 234571 578765 234755 578799
rect 234721 578731 234755 578765
rect 241529 578731 241563 578901
rect 251097 578799 251131 578901
rect 282871 578901 282929 578935
rect 253891 578765 254075 578799
rect 254041 578731 254075 578765
rect 268393 578527 268427 578765
rect 270417 578663 270451 578833
rect 270509 578663 270543 578901
rect 278053 578527 278087 578765
rect 284125 578527 284159 578765
rect 292497 578663 292531 578901
rect 294429 578527 294463 578765
rect 306389 578527 306423 578697
rect 310989 578663 311023 579309
rect 312001 578731 312035 578765
rect 311851 578697 312035 578731
rect 315221 578595 315255 579309
rect 317429 578459 317463 579309
rect 318809 578799 318843 578901
rect 323593 578799 323627 578901
rect 336657 578391 336691 579309
rect 343005 578323 343039 579309
rect 364257 578255 364291 579309
rect 153301 563023 153335 563125
rect 200129 562003 200163 562105
rect 208777 561935 208811 562105
rect 153301 550647 153335 560201
rect 96537 518755 96571 518925
rect 115949 518687 115983 518925
rect 125517 518823 125551 518925
rect 153393 502367 153427 505121
rect 380725 500939 380759 503081
rect 288357 492711 288391 497097
rect 288265 476051 288299 482953
rect 288265 463811 288299 466497
rect 299857 466395 299891 473297
rect 153485 456739 153519 463641
rect 288265 456739 288299 463641
rect 288357 444431 288391 447185
rect 299857 447083 299891 453985
rect 153393 437427 153427 444329
rect 288265 437427 288299 444329
rect 304181 434775 304215 452557
rect 288357 425119 288391 427873
rect 299857 427771 299891 434673
rect 118433 405739 118467 415361
rect 128553 405739 128587 415361
rect 132877 405739 132911 407881
rect 222209 406759 222243 406861
rect 202889 406555 202923 406725
rect 212457 406623 212491 406725
rect 215217 406725 215401 406759
rect 215217 406623 215251 406725
rect 231777 406691 231811 406861
rect 241529 406759 241563 406861
rect 251097 406691 251131 406861
rect 234571 406657 234629 406691
rect 253891 406657 253949 406691
rect 260849 406555 260883 406725
rect 289829 406623 289863 406725
rect 266093 406419 266127 406521
rect 299857 405739 299891 415361
rect 84025 395607 84059 395709
rect 84117 395607 84151 395845
rect 128553 394723 128587 404277
rect 153393 396083 153427 398905
rect 153301 389147 153335 395913
rect 128829 376771 128863 388433
rect 304273 379355 304307 386325
rect 132693 366979 132727 375309
rect 133153 358683 133187 367013
rect 153485 357459 153519 367013
rect 288357 362967 288391 369869
rect 288357 353311 288391 360213
rect 304273 347871 304307 357221
rect 132877 340595 132911 342057
rect 153393 340459 153427 340969
rect 288173 338147 288207 344573
rect 133153 333319 133187 337977
rect 241345 337875 241379 337977
rect 233525 337195 233559 337773
rect 251649 337331 251683 337637
rect 213929 328491 213963 331313
rect 129013 318903 129047 328389
rect 128645 307819 128679 317373
rect 209789 309179 209823 318733
rect 257721 317475 257755 335257
rect 288357 328491 288391 331993
rect 503729 328559 503763 331245
rect 288173 318835 288207 328321
rect 288357 309179 288391 313361
rect 304273 309247 304307 318733
rect 503729 317475 503763 321657
rect 503913 321555 503947 321725
rect 504005 318835 504039 321657
rect 504281 317475 504315 327029
rect 209789 289867 209823 299421
rect 257813 298163 257847 307717
rect 288357 299523 288391 302209
rect 304273 301699 304307 309077
rect 504373 299523 504407 312613
rect 288357 289867 288391 294049
rect 304273 289935 304307 299421
rect 128829 280211 128863 289765
rect 126069 270555 126103 280109
rect 153393 273275 153427 280109
rect 209789 270555 209823 280109
rect 257813 278783 257847 288269
rect 288173 280211 288207 289697
rect 304273 282795 304307 289765
rect 504465 288439 504499 298061
rect 288357 270555 288391 274737
rect 304273 270623 304307 280109
rect 128921 260899 128955 263585
rect 153577 260899 153611 270453
rect 257813 263551 257847 270453
rect 288173 260899 288207 270385
rect 504465 269127 504499 278681
rect 126069 251311 126103 260797
rect 209789 251311 209823 260797
rect 257813 253827 257847 260797
rect 304089 251311 304123 260797
rect 504281 253827 504315 260797
rect 304215 251209 304365 251243
rect 257721 241519 257755 251141
rect 288265 241519 288299 251141
rect 304181 241519 304215 244273
rect 504281 241519 504315 251141
rect 129013 231931 129047 236725
rect 288357 231863 288391 235977
rect 304181 231863 304215 241349
rect 153209 222207 153243 224961
rect 504373 222207 504407 231761
rect 126437 205547 126471 205649
rect 153301 202895 153335 212449
rect 304089 202895 304123 205649
rect 504189 202895 504223 205649
rect 199945 202351 199979 202793
rect 239597 202691 239631 202793
rect 199945 202317 200037 202351
rect 199945 202079 199979 202249
rect 199887 202045 199979 202079
rect 211813 201875 211847 202317
rect 215217 201399 215251 202249
rect 215861 201467 215895 201841
rect 216229 201535 216263 201841
rect 219265 201603 219299 202249
rect 216965 201399 216999 201569
rect 219357 201535 219391 202317
rect 223129 201535 223163 201705
rect 229109 201535 229143 202317
rect 229201 201603 229235 202249
rect 233525 202045 233743 202079
rect 233525 201603 233559 202045
rect 233709 202011 233743 202045
rect 238585 202011 238619 202249
rect 233617 201603 233651 201977
rect 236561 201807 236595 201977
rect 237389 201807 237423 201977
rect 236561 201773 236837 201807
rect 238677 201535 238711 202317
rect 239137 201603 239171 201909
rect 239505 201535 239539 202657
rect 253857 202555 253891 202657
rect 244841 201875 244875 202453
rect 248797 202283 248831 202521
rect 255605 202351 255639 202589
rect 258641 202487 258675 202725
rect 257997 202249 258273 202283
rect 257997 202215 258031 202249
rect 258365 201603 258399 202317
rect 258825 201535 258859 202793
rect 262229 201535 262263 202317
rect 264069 201875 264103 202181
rect 302249 201535 302283 202657
rect 302433 202555 302467 202725
rect 302893 202419 302927 202521
rect 302985 202079 303019 202385
rect 304917 201739 304951 202589
rect 306297 201807 306331 201977
rect 308505 201943 308539 202385
rect 311357 202079 311391 202453
rect 315681 201739 315715 202793
rect 318349 202011 318383 202725
rect 347697 202623 347731 202725
rect 351929 202147 351963 202725
rect 375573 202555 375607 202793
rect 375481 202351 375515 202521
rect 374377 202215 374411 202317
rect 374285 201671 374319 202181
rect 416145 201875 416179 202453
rect 417065 201671 417099 202181
rect 131497 196027 131531 198305
rect 131773 195959 131807 196061
rect 132877 195959 132911 196061
rect 131129 183379 131163 186269
rect 128921 171139 128955 180761
rect 99331 154513 99515 154547
rect 57989 154343 58023 154513
rect 99481 154479 99515 154513
rect 118651 154445 118835 154479
rect 67557 154343 67591 154445
rect 118801 154411 118835 154445
rect 80103 154377 80161 154411
rect 108991 153085 109049 153119
rect 17969 152779 18003 152881
rect 22753 152779 22787 153017
rect 27629 152915 27663 153017
rect 32413 152915 32447 153085
rect 77309 152847 77343 152949
rect 86877 152847 86911 153017
rect 131221 147679 131255 157301
rect 131313 151895 131347 153085
rect 80011 144857 80195 144891
rect 41371 144721 41429 144755
rect 60691 144721 60749 144755
rect 29009 144551 29043 144653
rect 38577 144551 38611 144721
rect 48329 144551 48363 144653
rect 57897 144551 57931 144721
rect 67649 144687 67683 144857
rect 80161 144755 80195 144857
rect 99331 144857 99515 144891
rect 86969 144619 87003 144721
rect 96537 144619 96571 144857
rect 99481 144823 99515 144857
rect 118651 144857 118835 144891
rect 109049 144755 109083 144857
rect 118801 144755 118835 144857
rect 132785 142171 132819 143565
rect 128829 133875 128863 142069
rect 134073 120479 134107 122349
rect 138581 120411 138615 120581
rect 143457 120411 143491 120581
rect 143549 120343 143583 120513
rect 151829 120207 151863 120309
rect 161397 120207 161431 120445
rect 171149 120343 171183 120445
rect 180717 120343 180751 120445
rect 182189 120275 182223 120445
rect 145021 118847 145055 120105
rect 89729 117759 89763 117929
rect 108957 117759 108991 117929
rect 115949 117759 115983 117997
rect 123769 117759 123803 117997
rect 123861 117963 123895 118133
rect 130761 117555 130795 117589
rect 135361 117555 135395 117657
rect 130761 117521 130945 117555
rect 135211 117521 135395 117555
rect 137937 117283 137971 117929
rect 138029 117283 138063 117929
rect 128921 99331 128955 106233
rect 145021 96679 145055 118813
rect 210433 118507 210467 118609
rect 210525 118303 210559 118473
rect 220093 118303 220127 118609
rect 219909 118201 220185 118235
rect 219909 117963 219943 118201
rect 147689 117487 147723 117929
rect 150449 117487 150483 117861
rect 154589 117487 154623 117861
rect 164157 117487 164191 117929
rect 220277 117827 220311 118269
rect 220369 117963 220403 118473
rect 237941 118201 238125 118235
rect 200405 117623 200439 117793
rect 220001 117793 220311 117827
rect 220001 117759 220035 117793
rect 220093 117419 220127 117725
rect 226257 117623 226291 117861
rect 229293 117419 229327 117861
rect 229845 117419 229879 117725
rect 237941 117487 237975 118201
rect 243645 117759 243679 118609
rect 253397 118507 253431 118609
rect 240551 117453 240701 117487
rect 249073 117351 249107 118473
rect 324881 117487 324915 118065
rect 359473 117895 359507 118133
rect 384313 118031 384347 118269
rect 325709 114563 325743 117725
rect 391213 117419 391247 117725
rect 398791 117521 398849 117555
rect 413201 117487 413235 117725
rect 396089 117283 396123 117385
rect 416789 117351 416823 117657
rect 416881 117555 416915 117861
rect 420745 117555 420779 117861
rect 422309 117623 422343 117793
rect 423045 117623 423079 117793
rect 427737 117691 427771 117793
rect 431693 117759 431727 118609
rect 431693 117725 431969 117759
rect 424149 117657 424425 117691
rect 427679 117657 427771 117691
rect 424149 117487 424183 117657
rect 424091 117453 424183 117487
rect 430221 117283 430255 117453
rect 433349 117283 433383 117453
rect 157533 99331 157567 106233
rect 174185 104907 174219 114461
rect 179521 99331 179555 106233
rect 138029 89675 138063 96577
rect 173909 95251 173943 97189
rect 140881 86887 140915 95149
rect 150633 85595 150667 95149
rect 162869 86887 162903 95149
rect 186237 93891 186271 103445
rect 215401 95251 215435 104805
rect 221013 96679 221047 106233
rect 229293 103547 229327 113101
rect 230397 103547 230431 114461
rect 248337 104907 248371 114461
rect 403909 106335 403943 115889
rect 420561 108987 420595 115889
rect 431509 108987 431543 115889
rect 216781 89539 216815 96577
rect 128645 75939 128679 85493
rect 140973 74579 141007 84133
rect 147965 75939 147999 85493
rect 192217 74579 192251 84133
rect 207305 77299 207339 80801
rect 214113 75939 214147 85493
rect 222301 82875 222335 100657
rect 223681 92531 223715 102085
rect 233341 93891 233375 103445
rect 240241 95251 240275 100045
rect 248337 95251 248371 100045
rect 276121 95251 276155 104805
rect 227913 82875 227947 92429
rect 271981 85595 272015 95149
rect 279709 93891 279743 103445
rect 301973 99331 302007 106233
rect 322673 99331 322707 106233
rect 290565 89403 290599 96577
rect 325709 95251 325743 104805
rect 394433 99331 394467 106233
rect 383117 87023 383151 96577
rect 388637 87023 388671 96577
rect 403909 87023 403943 96577
rect 415041 95251 415075 104805
rect 420653 87023 420687 96577
rect 426265 95319 426299 104805
rect 431601 87023 431635 104805
rect 216873 79951 216907 80121
rect 223681 74579 223715 80121
rect 229201 74579 229235 80121
rect 230397 74579 230431 84133
rect 232145 79951 232179 80121
rect 244289 70295 244323 75837
rect 245761 70363 245795 75837
rect 248429 74579 248463 84133
rect 128829 56627 128863 66181
rect 125977 46971 126011 51085
rect 140881 48331 140915 57817
rect 144929 55267 144963 64821
rect 157349 55267 157383 64821
rect 162961 56627 162995 66181
rect 214205 56627 214239 66181
rect 216873 61047 216907 67541
rect 238953 57987 238987 67541
rect 271889 66283 271923 75837
rect 279709 66283 279743 84133
rect 290565 79951 290599 86921
rect 322673 77299 322707 86921
rect 301973 67643 302007 77129
rect 325709 75939 325743 85493
rect 394433 77299 394467 86921
rect 426173 85595 426207 86989
rect 341349 67643 341383 77129
rect 383209 67643 383243 77129
rect 388729 67643 388763 77129
rect 404001 67643 404035 77129
rect 426081 69683 426115 84133
rect 431601 66283 431635 75837
rect 133337 37315 133371 46869
rect 150633 37315 150667 46869
rect 157625 38675 157659 51765
rect 179429 46971 179463 56525
rect 162961 37315 162995 46869
rect 186237 45611 186271 55165
rect 192125 46971 192159 56525
rect 125977 9707 126011 27557
rect 133337 19295 133371 27557
rect 140881 19431 140915 28917
rect 140881 9707 140915 19261
rect 161765 11883 161799 22729
rect 162961 18003 162995 27557
rect 174001 26299 174035 40681
rect 179429 27659 179463 37213
rect 183753 27659 183787 45509
rect 190653 40715 190687 45509
rect 192125 41327 192159 45849
rect 186237 27115 186271 40681
rect 207489 38675 207523 56525
rect 280077 51051 280111 57885
rect 290473 55267 290507 64821
rect 214113 37315 214147 46869
rect 215401 37315 215435 46869
rect 248337 37315 248371 46869
rect 271889 41327 271923 48161
rect 290381 47039 290415 51153
rect 301789 48331 301823 57885
rect 322673 48331 322707 57885
rect 325525 56627 325559 66181
rect 192217 27591 192251 31705
rect 244289 31671 244323 37213
rect 245761 31671 245795 37213
rect 271889 29019 271923 38573
rect 276121 29087 276155 46733
rect 290657 38539 290691 46869
rect 322673 29019 322707 38573
rect 325709 29087 325743 46869
rect 341533 45611 341567 51153
rect 383209 48331 383243 57885
rect 388729 48331 388763 57885
rect 404001 48331 404035 57885
rect 415041 56627 415075 66181
rect 341441 38267 341475 45441
rect 383209 29019 383243 38573
rect 404001 29019 404035 38573
rect 414949 35955 414983 45509
rect 425989 37315 426023 46869
rect 431601 31671 431635 37213
rect 168389 9707 168423 12461
rect 179705 9707 179739 19261
rect 183753 16643 183787 26197
rect 190469 18003 190503 27557
rect 192217 16643 192251 26197
rect 207489 19431 207523 28917
rect 207213 9707 207247 19261
rect 214113 9707 214147 27557
rect 215401 9707 215435 27557
rect 222301 23511 222335 24905
rect 123125 7259 123159 7361
rect 125609 6987 125643 8313
rect 227821 6919 227855 20009
rect 230121 6919 230155 24769
rect 238953 19363 238987 22185
rect 238401 9707 238435 19261
rect 276121 18003 276155 27557
rect 279985 19363 280019 28917
rect 274833 9707 274867 15861
rect 290933 9707 290967 19261
rect 301881 8347 301915 26197
rect 325709 9707 325743 27557
rect 383393 19363 383427 25245
rect 415041 16643 415075 26197
rect 420469 18003 420503 27557
rect 431509 16643 431543 26197
rect 383301 9707 383335 12529
rect 414799 8245 415041 8279
rect 412649 7055 412683 7565
rect 55229 3179 55263 4097
rect 64797 3179 64831 4097
rect 74549 3179 74583 4097
rect 84117 3179 84151 4097
rect 93869 2975 93903 4097
rect 103437 2975 103471 4097
rect 113189 2907 113223 4097
rect 123493 2907 123527 4097
rect 133153 2907 133187 4097
rect 142813 2907 142847 4097
rect 148885 4063 148919 4097
rect 148885 4029 149069 4063
rect 355367 4029 355517 4063
rect 217885 3587 217919 3825
rect 218069 3791 218103 4029
rect 194609 3179 194643 3281
rect 210065 3247 210099 3417
rect 217241 3247 217275 3485
rect 225245 3383 225279 3825
rect 228833 3383 228867 3621
rect 229753 3519 229787 3893
rect 234629 3383 234663 3553
rect 326445 595 326479 3757
rect 340245 3587 340279 3689
rect 355241 3587 355275 3961
rect 398849 3655 398883 3825
rect 407405 3519 407439 3757
rect 417985 3519 418019 3621
rect 418203 3485 418295 3519
rect 418261 2975 418295 3485
rect 427737 2975 427771 3553
rect 422309 2771 422343 2941
rect 432521 2771 432555 3417
rect 437397 2975 437431 3417
rect 442273 2907 442307 3485
rect 482109 3281 482385 3315
rect 480913 3043 480947 3213
rect 463709 2907 463743 3009
rect 473277 2839 473311 3009
rect 481005 2975 481039 3213
rect 482109 2975 482143 3281
rect 485145 2975 485179 3213
rect 481097 2907 481131 2941
rect 480821 2873 481131 2907
rect 480821 2839 480855 2873
rect 485053 2839 485087 2941
rect 485697 2907 485731 3281
rect 489561 3043 489595 3281
rect 489101 2975 489135 3009
rect 489653 2975 489687 3281
rect 496645 3179 496679 3281
rect 504373 3247 504407 3349
rect 504557 3315 504591 4097
rect 489101 2941 489687 2975
rect 483029 2703 483063 2805
<< viali >>
rect 153577 684437 153611 684471
rect 153577 666553 153611 666587
rect 153485 656829 153519 656863
rect 153485 647241 153519 647275
rect 153393 579581 153427 579615
rect 142813 578765 142847 578799
rect 142813 578493 142847 578527
rect 310989 579309 311023 579343
rect 183569 578901 183603 578935
rect 154589 578833 154623 578867
rect 154589 578697 154623 578731
rect 164157 578833 164191 578867
rect 176577 578765 176611 578799
rect 176669 578765 176703 578799
rect 164157 578697 164191 578731
rect 193137 578901 193171 578935
rect 202889 578901 202923 578935
rect 193137 578765 193171 578799
rect 195897 578765 195931 578799
rect 183569 578697 183603 578731
rect 196081 578697 196115 578731
rect 212457 578901 212491 578935
rect 222209 578901 222243 578935
rect 212457 578765 212491 578799
rect 215217 578765 215251 578799
rect 202889 578697 202923 578731
rect 215401 578697 215435 578731
rect 231777 578901 231811 578935
rect 241529 578901 241563 578935
rect 231777 578765 231811 578799
rect 234537 578765 234571 578799
rect 222209 578697 222243 578731
rect 234721 578697 234755 578731
rect 251097 578901 251131 578935
rect 270509 578901 270543 578935
rect 282837 578901 282871 578935
rect 282929 578901 282963 578935
rect 292497 578901 292531 578935
rect 270417 578833 270451 578867
rect 251097 578765 251131 578799
rect 253857 578765 253891 578799
rect 241529 578697 241563 578731
rect 254041 578697 254075 578731
rect 268393 578765 268427 578799
rect 270417 578629 270451 578663
rect 270509 578629 270543 578663
rect 278053 578765 278087 578799
rect 268393 578493 268427 578527
rect 278053 578493 278087 578527
rect 284125 578765 284159 578799
rect 292497 578629 292531 578663
rect 294429 578765 294463 578799
rect 284125 578493 284159 578527
rect 294429 578493 294463 578527
rect 306389 578697 306423 578731
rect 315221 579309 315255 579343
rect 312001 578765 312035 578799
rect 311817 578697 311851 578731
rect 310989 578629 311023 578663
rect 315221 578561 315255 578595
rect 317429 579309 317463 579343
rect 306389 578493 306423 578527
rect 336657 579309 336691 579343
rect 318809 578901 318843 578935
rect 318809 578765 318843 578799
rect 323593 578901 323627 578935
rect 323593 578765 323627 578799
rect 317429 578425 317463 578459
rect 336657 578357 336691 578391
rect 343005 579309 343039 579343
rect 343005 578289 343039 578323
rect 364257 579309 364291 579343
rect 364257 578221 364291 578255
rect 153393 569925 153427 569959
rect 153301 563125 153335 563159
rect 153301 562989 153335 563023
rect 200129 562105 200163 562139
rect 200129 561969 200163 562003
rect 208777 562105 208811 562139
rect 208777 561901 208811 561935
rect 153301 560201 153335 560235
rect 153301 550613 153335 550647
rect 96537 518925 96571 518959
rect 96537 518721 96571 518755
rect 115949 518925 115983 518959
rect 125517 518925 125551 518959
rect 125517 518789 125551 518823
rect 115949 518653 115983 518687
rect 153393 505121 153427 505155
rect 153393 502333 153427 502367
rect 380725 503081 380759 503115
rect 380725 500905 380759 500939
rect 288357 497097 288391 497131
rect 288357 492677 288391 492711
rect 288265 482953 288299 482987
rect 288265 476017 288299 476051
rect 299857 473297 299891 473331
rect 288265 466497 288299 466531
rect 299857 466361 299891 466395
rect 288265 463777 288299 463811
rect 153485 463641 153519 463675
rect 153485 456705 153519 456739
rect 288265 463641 288299 463675
rect 288265 456705 288299 456739
rect 299857 453985 299891 454019
rect 288357 447185 288391 447219
rect 299857 447049 299891 447083
rect 304181 452557 304215 452591
rect 288357 444397 288391 444431
rect 153393 444329 153427 444363
rect 153393 437393 153427 437427
rect 288265 444329 288299 444363
rect 288265 437393 288299 437427
rect 304181 434741 304215 434775
rect 299857 434673 299891 434707
rect 288357 427873 288391 427907
rect 299857 427737 299891 427771
rect 288357 425085 288391 425119
rect 118433 415361 118467 415395
rect 118433 405705 118467 405739
rect 128553 415361 128587 415395
rect 299857 415361 299891 415395
rect 128553 405705 128587 405739
rect 132877 407881 132911 407915
rect 222209 406861 222243 406895
rect 202889 406725 202923 406759
rect 212457 406725 212491 406759
rect 212457 406589 212491 406623
rect 215401 406725 215435 406759
rect 222209 406725 222243 406759
rect 231777 406861 231811 406895
rect 241529 406861 241563 406895
rect 241529 406725 241563 406759
rect 251097 406861 251131 406895
rect 260849 406725 260883 406759
rect 231777 406657 231811 406691
rect 234537 406657 234571 406691
rect 234629 406657 234663 406691
rect 251097 406657 251131 406691
rect 253857 406657 253891 406691
rect 253949 406657 253983 406691
rect 215217 406589 215251 406623
rect 202889 406521 202923 406555
rect 289829 406725 289863 406759
rect 289829 406589 289863 406623
rect 260849 406521 260883 406555
rect 266093 406521 266127 406555
rect 266093 406385 266127 406419
rect 132877 405705 132911 405739
rect 299857 405705 299891 405739
rect 128553 404277 128587 404311
rect 84117 395845 84151 395879
rect 84025 395709 84059 395743
rect 84025 395573 84059 395607
rect 84117 395573 84151 395607
rect 153393 398905 153427 398939
rect 153393 396049 153427 396083
rect 128553 394689 128587 394723
rect 153301 395913 153335 395947
rect 153301 389113 153335 389147
rect 128829 388433 128863 388467
rect 304273 386325 304307 386359
rect 304273 379321 304307 379355
rect 128829 376737 128863 376771
rect 132693 375309 132727 375343
rect 288357 369869 288391 369903
rect 132693 366945 132727 366979
rect 133153 367013 133187 367047
rect 133153 358649 133187 358683
rect 153485 367013 153519 367047
rect 288357 362933 288391 362967
rect 153485 357425 153519 357459
rect 288357 360213 288391 360247
rect 288357 353277 288391 353311
rect 304273 357221 304307 357255
rect 304273 347837 304307 347871
rect 288173 344573 288207 344607
rect 132877 342057 132911 342091
rect 132877 340561 132911 340595
rect 153393 340969 153427 341003
rect 153393 340425 153427 340459
rect 288173 338113 288207 338147
rect 133153 337977 133187 338011
rect 241345 337977 241379 338011
rect 241345 337841 241379 337875
rect 233525 337773 233559 337807
rect 251649 337637 251683 337671
rect 251649 337297 251683 337331
rect 233525 337161 233559 337195
rect 133153 333285 133187 333319
rect 257721 335257 257755 335291
rect 213929 331313 213963 331347
rect 213929 328457 213963 328491
rect 129013 328389 129047 328423
rect 129013 318869 129047 318903
rect 209789 318733 209823 318767
rect 128645 317373 128679 317407
rect 288357 331993 288391 332027
rect 503729 331245 503763 331279
rect 503729 328525 503763 328559
rect 288357 328457 288391 328491
rect 288173 328321 288207 328355
rect 504281 327029 504315 327063
rect 503913 321725 503947 321759
rect 288173 318801 288207 318835
rect 503729 321657 503763 321691
rect 257721 317441 257755 317475
rect 304273 318733 304307 318767
rect 209789 309145 209823 309179
rect 288357 313361 288391 313395
rect 503913 321521 503947 321555
rect 504005 321657 504039 321691
rect 504005 318801 504039 318835
rect 503729 317441 503763 317475
rect 504281 317441 504315 317475
rect 304273 309213 304307 309247
rect 504373 312613 504407 312647
rect 288357 309145 288391 309179
rect 128645 307785 128679 307819
rect 304273 309077 304307 309111
rect 257813 307717 257847 307751
rect 209789 299421 209823 299455
rect 288357 302209 288391 302243
rect 304273 301665 304307 301699
rect 288357 299489 288391 299523
rect 504373 299489 504407 299523
rect 257813 298129 257847 298163
rect 304273 299421 304307 299455
rect 209789 289833 209823 289867
rect 288357 294049 288391 294083
rect 304273 289901 304307 289935
rect 504465 298061 504499 298095
rect 288357 289833 288391 289867
rect 128829 289765 128863 289799
rect 304273 289765 304307 289799
rect 288173 289697 288207 289731
rect 128829 280177 128863 280211
rect 257813 288269 257847 288303
rect 126069 280109 126103 280143
rect 153393 280109 153427 280143
rect 153393 273241 153427 273275
rect 209789 280109 209823 280143
rect 126069 270521 126103 270555
rect 504465 288405 504499 288439
rect 304273 282761 304307 282795
rect 288173 280177 288207 280211
rect 257813 278749 257847 278783
rect 304273 280109 304307 280143
rect 209789 270521 209823 270555
rect 288357 274737 288391 274771
rect 304273 270589 304307 270623
rect 504465 278681 504499 278715
rect 288357 270521 288391 270555
rect 153577 270453 153611 270487
rect 128921 263585 128955 263619
rect 128921 260865 128955 260899
rect 257813 270453 257847 270487
rect 257813 263517 257847 263551
rect 288173 270385 288207 270419
rect 153577 260865 153611 260899
rect 504465 269093 504499 269127
rect 288173 260865 288207 260899
rect 126069 260797 126103 260831
rect 126069 251277 126103 251311
rect 209789 260797 209823 260831
rect 257813 260797 257847 260831
rect 257813 253793 257847 253827
rect 304089 260797 304123 260831
rect 209789 251277 209823 251311
rect 504281 260797 504315 260831
rect 504281 253793 504315 253827
rect 304089 251277 304123 251311
rect 304181 251209 304215 251243
rect 304365 251209 304399 251243
rect 257721 251141 257755 251175
rect 257721 241485 257755 241519
rect 288265 251141 288299 251175
rect 504281 251141 504315 251175
rect 288265 241485 288299 241519
rect 304181 244273 304215 244307
rect 304181 241485 304215 241519
rect 504281 241485 504315 241519
rect 304181 241349 304215 241383
rect 129013 236725 129047 236759
rect 129013 231897 129047 231931
rect 288357 235977 288391 236011
rect 288357 231829 288391 231863
rect 304181 231829 304215 231863
rect 504373 231761 504407 231795
rect 153209 224961 153243 224995
rect 153209 222173 153243 222207
rect 504373 222173 504407 222207
rect 153301 212449 153335 212483
rect 126437 205649 126471 205683
rect 126437 205513 126471 205547
rect 153301 202861 153335 202895
rect 304089 205649 304123 205683
rect 304089 202861 304123 202895
rect 504189 205649 504223 205683
rect 504189 202861 504223 202895
rect 199945 202793 199979 202827
rect 239597 202793 239631 202827
rect 258825 202793 258859 202827
rect 258641 202725 258675 202759
rect 239505 202657 239539 202691
rect 239597 202657 239631 202691
rect 253857 202657 253891 202691
rect 200037 202317 200071 202351
rect 211813 202317 211847 202351
rect 199945 202249 199979 202283
rect 199853 202045 199887 202079
rect 219357 202317 219391 202351
rect 211813 201841 211847 201875
rect 215217 202249 215251 202283
rect 219265 202249 219299 202283
rect 215861 201841 215895 201875
rect 216229 201841 216263 201875
rect 216229 201501 216263 201535
rect 216965 201569 216999 201603
rect 219265 201569 219299 201603
rect 215861 201433 215895 201467
rect 215217 201365 215251 201399
rect 229109 202317 229143 202351
rect 219357 201501 219391 201535
rect 223129 201705 223163 201739
rect 223129 201501 223163 201535
rect 238677 202317 238711 202351
rect 229201 202249 229235 202283
rect 238585 202249 238619 202283
rect 229201 201569 229235 201603
rect 233525 201569 233559 201603
rect 233617 201977 233651 202011
rect 233709 201977 233743 202011
rect 236561 201977 236595 202011
rect 237389 201977 237423 202011
rect 238585 201977 238619 202011
rect 236837 201773 236871 201807
rect 237389 201773 237423 201807
rect 233617 201569 233651 201603
rect 229109 201501 229143 201535
rect 239137 201909 239171 201943
rect 239137 201569 239171 201603
rect 238677 201501 238711 201535
rect 248797 202521 248831 202555
rect 253857 202521 253891 202555
rect 255605 202589 255639 202623
rect 244841 202453 244875 202487
rect 258641 202453 258675 202487
rect 255605 202317 255639 202351
rect 258365 202317 258399 202351
rect 248797 202249 248831 202283
rect 258273 202249 258307 202283
rect 257997 202181 258031 202215
rect 244841 201841 244875 201875
rect 258365 201569 258399 201603
rect 239505 201501 239539 201535
rect 315681 202793 315715 202827
rect 302433 202725 302467 202759
rect 302249 202657 302283 202691
rect 258825 201501 258859 201535
rect 262229 202317 262263 202351
rect 264069 202181 264103 202215
rect 264069 201841 264103 201875
rect 262229 201501 262263 201535
rect 304917 202589 304951 202623
rect 302433 202521 302467 202555
rect 302893 202521 302927 202555
rect 302893 202385 302927 202419
rect 302985 202385 303019 202419
rect 302985 202045 303019 202079
rect 311357 202453 311391 202487
rect 308505 202385 308539 202419
rect 306297 201977 306331 202011
rect 311357 202045 311391 202079
rect 308505 201909 308539 201943
rect 306297 201773 306331 201807
rect 304917 201705 304951 201739
rect 375573 202793 375607 202827
rect 318349 202725 318383 202759
rect 347697 202725 347731 202759
rect 347697 202589 347731 202623
rect 351929 202725 351963 202759
rect 375481 202521 375515 202555
rect 375573 202521 375607 202555
rect 374377 202317 374411 202351
rect 375481 202317 375515 202351
rect 416145 202453 416179 202487
rect 351929 202113 351963 202147
rect 374285 202181 374319 202215
rect 374377 202181 374411 202215
rect 318349 201977 318383 202011
rect 315681 201705 315715 201739
rect 416145 201841 416179 201875
rect 417065 202181 417099 202215
rect 374285 201637 374319 201671
rect 417065 201637 417099 201671
rect 302249 201501 302283 201535
rect 216965 201365 216999 201399
rect 131497 198305 131531 198339
rect 131497 195993 131531 196027
rect 131773 196061 131807 196095
rect 131773 195925 131807 195959
rect 132877 196061 132911 196095
rect 132877 195925 132911 195959
rect 131129 186269 131163 186303
rect 131129 183345 131163 183379
rect 128921 180761 128955 180795
rect 128921 171105 128955 171139
rect 131221 157301 131255 157335
rect 57989 154513 58023 154547
rect 99297 154513 99331 154547
rect 57989 154309 58023 154343
rect 67557 154445 67591 154479
rect 99481 154445 99515 154479
rect 118617 154445 118651 154479
rect 80069 154377 80103 154411
rect 80161 154377 80195 154411
rect 118801 154377 118835 154411
rect 67557 154309 67591 154343
rect 32413 153085 32447 153119
rect 108957 153085 108991 153119
rect 109049 153085 109083 153119
rect 22753 153017 22787 153051
rect 17969 152881 18003 152915
rect 17969 152745 18003 152779
rect 27629 153017 27663 153051
rect 27629 152881 27663 152915
rect 86877 153017 86911 153051
rect 32413 152881 32447 152915
rect 77309 152949 77343 152983
rect 77309 152813 77343 152847
rect 86877 152813 86911 152847
rect 22753 152745 22787 152779
rect 131313 153085 131347 153119
rect 131313 151861 131347 151895
rect 131221 147645 131255 147679
rect 67649 144857 67683 144891
rect 79977 144857 80011 144891
rect 38577 144721 38611 144755
rect 41337 144721 41371 144755
rect 41429 144721 41463 144755
rect 57897 144721 57931 144755
rect 60657 144721 60691 144755
rect 60749 144721 60783 144755
rect 29009 144653 29043 144687
rect 29009 144517 29043 144551
rect 38577 144517 38611 144551
rect 48329 144653 48363 144687
rect 48329 144517 48363 144551
rect 96537 144857 96571 144891
rect 99297 144857 99331 144891
rect 80161 144721 80195 144755
rect 86969 144721 87003 144755
rect 67649 144653 67683 144687
rect 86969 144585 87003 144619
rect 99481 144789 99515 144823
rect 109049 144857 109083 144891
rect 118617 144857 118651 144891
rect 109049 144721 109083 144755
rect 118801 144721 118835 144755
rect 96537 144585 96571 144619
rect 57897 144517 57931 144551
rect 132785 143565 132819 143599
rect 132785 142137 132819 142171
rect 128829 142069 128863 142103
rect 128829 133841 128863 133875
rect 134073 122349 134107 122383
rect 134073 120445 134107 120479
rect 138581 120581 138615 120615
rect 138581 120377 138615 120411
rect 143457 120581 143491 120615
rect 143457 120377 143491 120411
rect 143549 120513 143583 120547
rect 161397 120445 161431 120479
rect 143549 120309 143583 120343
rect 151829 120309 151863 120343
rect 151829 120173 151863 120207
rect 171149 120445 171183 120479
rect 171149 120309 171183 120343
rect 180717 120445 180751 120479
rect 180717 120309 180751 120343
rect 182189 120445 182223 120479
rect 182189 120241 182223 120275
rect 161397 120173 161431 120207
rect 145021 120105 145055 120139
rect 145021 118813 145055 118847
rect 123861 118133 123895 118167
rect 115949 117997 115983 118031
rect 89729 117929 89763 117963
rect 89729 117725 89763 117759
rect 108957 117929 108991 117963
rect 108957 117725 108991 117759
rect 115949 117725 115983 117759
rect 123769 117997 123803 118031
rect 123861 117929 123895 117963
rect 137937 117929 137971 117963
rect 123769 117725 123803 117759
rect 135361 117657 135395 117691
rect 130761 117589 130795 117623
rect 130945 117521 130979 117555
rect 135177 117521 135211 117555
rect 137937 117249 137971 117283
rect 138029 117929 138063 117963
rect 138029 117249 138063 117283
rect 128921 106233 128955 106267
rect 128921 99297 128955 99331
rect 210433 118609 210467 118643
rect 220093 118609 220127 118643
rect 210433 118473 210467 118507
rect 210525 118473 210559 118507
rect 210525 118269 210559 118303
rect 243645 118609 243679 118643
rect 220369 118473 220403 118507
rect 220093 118269 220127 118303
rect 220277 118269 220311 118303
rect 220185 118201 220219 118235
rect 147689 117929 147723 117963
rect 164157 117929 164191 117963
rect 219909 117929 219943 117963
rect 147689 117453 147723 117487
rect 150449 117861 150483 117895
rect 150449 117453 150483 117487
rect 154589 117861 154623 117895
rect 154589 117453 154623 117487
rect 220369 117929 220403 117963
rect 238125 118201 238159 118235
rect 200405 117793 200439 117827
rect 226257 117861 226291 117895
rect 220001 117725 220035 117759
rect 220093 117725 220127 117759
rect 200405 117589 200439 117623
rect 164157 117453 164191 117487
rect 226257 117589 226291 117623
rect 229293 117861 229327 117895
rect 220093 117385 220127 117419
rect 229293 117385 229327 117419
rect 229845 117725 229879 117759
rect 253397 118609 253431 118643
rect 243645 117725 243679 117759
rect 249073 118473 249107 118507
rect 253397 118473 253431 118507
rect 431693 118609 431727 118643
rect 237941 117453 237975 117487
rect 240517 117453 240551 117487
rect 240701 117453 240735 117487
rect 229845 117385 229879 117419
rect 384313 118269 384347 118303
rect 359473 118133 359507 118167
rect 324881 118065 324915 118099
rect 384313 117997 384347 118031
rect 359473 117861 359507 117895
rect 416881 117861 416915 117895
rect 324881 117453 324915 117487
rect 325709 117725 325743 117759
rect 249073 117317 249107 117351
rect 391213 117725 391247 117759
rect 413201 117725 413235 117759
rect 398757 117521 398791 117555
rect 398849 117521 398883 117555
rect 413201 117453 413235 117487
rect 416789 117657 416823 117691
rect 391213 117385 391247 117419
rect 396089 117385 396123 117419
rect 416881 117521 416915 117555
rect 420745 117861 420779 117895
rect 422309 117793 422343 117827
rect 422309 117589 422343 117623
rect 423045 117793 423079 117827
rect 427737 117793 427771 117827
rect 431969 117725 432003 117759
rect 423045 117589 423079 117623
rect 424425 117657 424459 117691
rect 427645 117657 427679 117691
rect 420745 117521 420779 117555
rect 424057 117453 424091 117487
rect 430221 117453 430255 117487
rect 416789 117317 416823 117351
rect 396089 117249 396123 117283
rect 430221 117249 430255 117283
rect 433349 117453 433383 117487
rect 433349 117249 433383 117283
rect 325709 114529 325743 114563
rect 403909 115889 403943 115923
rect 174185 114461 174219 114495
rect 157533 106233 157567 106267
rect 230397 114461 230431 114495
rect 229293 113101 229327 113135
rect 174185 104873 174219 104907
rect 179521 106233 179555 106267
rect 157533 99297 157567 99331
rect 221013 106233 221047 106267
rect 215401 104805 215435 104839
rect 179521 99297 179555 99331
rect 186237 103445 186271 103479
rect 145021 96645 145055 96679
rect 173909 97189 173943 97223
rect 138029 96577 138063 96611
rect 173909 95217 173943 95251
rect 138029 89641 138063 89675
rect 140881 95149 140915 95183
rect 140881 86853 140915 86887
rect 150633 95149 150667 95183
rect 162869 95149 162903 95183
rect 229293 103513 229327 103547
rect 248337 114461 248371 114495
rect 420561 115889 420595 115923
rect 420561 108953 420595 108987
rect 431509 115889 431543 115923
rect 431509 108953 431543 108987
rect 403909 106301 403943 106335
rect 248337 104873 248371 104907
rect 301973 106233 302007 106267
rect 230397 103513 230431 103547
rect 276121 104805 276155 104839
rect 233341 103445 233375 103479
rect 223681 102085 223715 102119
rect 221013 96645 221047 96679
rect 222301 100657 222335 100691
rect 215401 95217 215435 95251
rect 216781 96577 216815 96611
rect 186237 93857 186271 93891
rect 216781 89505 216815 89539
rect 162869 86853 162903 86887
rect 150633 85561 150667 85595
rect 128645 85493 128679 85527
rect 147965 85493 147999 85527
rect 128645 75905 128679 75939
rect 140973 84133 141007 84167
rect 214113 85493 214147 85527
rect 147965 75905 147999 75939
rect 192217 84133 192251 84167
rect 140973 74545 141007 74579
rect 207305 80801 207339 80835
rect 207305 77265 207339 77299
rect 240241 100045 240275 100079
rect 240241 95217 240275 95251
rect 248337 100045 248371 100079
rect 248337 95217 248371 95251
rect 276121 95217 276155 95251
rect 279709 103445 279743 103479
rect 233341 93857 233375 93891
rect 271981 95149 272015 95183
rect 223681 92497 223715 92531
rect 222301 82841 222335 82875
rect 227913 92429 227947 92463
rect 301973 99297 302007 99331
rect 322673 106233 322707 106267
rect 394433 106233 394467 106267
rect 322673 99297 322707 99331
rect 325709 104805 325743 104839
rect 279709 93857 279743 93891
rect 290565 96577 290599 96611
rect 394433 99297 394467 99331
rect 415041 104805 415075 104839
rect 325709 95217 325743 95251
rect 383117 96577 383151 96611
rect 290565 89369 290599 89403
rect 383117 86989 383151 87023
rect 388637 96577 388671 96611
rect 388637 86989 388671 87023
rect 403909 96577 403943 96611
rect 426265 104805 426299 104839
rect 415041 95217 415075 95251
rect 420653 96577 420687 96611
rect 403909 86989 403943 87023
rect 426265 95285 426299 95319
rect 431601 104805 431635 104839
rect 420653 86989 420687 87023
rect 426173 86989 426207 87023
rect 431601 86989 431635 87023
rect 271981 85561 272015 85595
rect 290565 86921 290599 86955
rect 227913 82841 227947 82875
rect 230397 84133 230431 84167
rect 216873 80121 216907 80155
rect 216873 79917 216907 79951
rect 223681 80121 223715 80155
rect 214113 75905 214147 75939
rect 192217 74545 192251 74579
rect 223681 74545 223715 74579
rect 229201 80121 229235 80155
rect 229201 74545 229235 74579
rect 248429 84133 248463 84167
rect 232145 80121 232179 80155
rect 232145 79917 232179 79951
rect 230397 74545 230431 74579
rect 244289 75837 244323 75871
rect 245761 75837 245795 75871
rect 279709 84133 279743 84167
rect 248429 74545 248463 74579
rect 271889 75837 271923 75871
rect 245761 70329 245795 70363
rect 244289 70261 244323 70295
rect 216873 67541 216907 67575
rect 128829 66181 128863 66215
rect 162961 66181 162995 66215
rect 144929 64821 144963 64855
rect 128829 56593 128863 56627
rect 140881 57817 140915 57851
rect 125977 51085 126011 51119
rect 144929 55233 144963 55267
rect 157349 64821 157383 64855
rect 162961 56593 162995 56627
rect 214205 66181 214239 66215
rect 216873 61013 216907 61047
rect 238953 67541 238987 67575
rect 271889 66249 271923 66283
rect 290565 79917 290599 79951
rect 322673 86921 322707 86955
rect 394433 86921 394467 86955
rect 322673 77265 322707 77299
rect 325709 85493 325743 85527
rect 301973 77129 302007 77163
rect 426173 85561 426207 85595
rect 394433 77265 394467 77299
rect 426081 84133 426115 84167
rect 325709 75905 325743 75939
rect 341349 77129 341383 77163
rect 301973 67609 302007 67643
rect 341349 67609 341383 67643
rect 383209 77129 383243 77163
rect 383209 67609 383243 67643
rect 388729 77129 388763 77163
rect 388729 67609 388763 67643
rect 404001 77129 404035 77163
rect 426081 69649 426115 69683
rect 431601 75837 431635 75871
rect 404001 67609 404035 67643
rect 279709 66249 279743 66283
rect 431601 66249 431635 66283
rect 325525 66181 325559 66215
rect 238953 57953 238987 57987
rect 290473 64821 290507 64855
rect 214205 56593 214239 56627
rect 280077 57885 280111 57919
rect 157349 55233 157383 55267
rect 179429 56525 179463 56559
rect 140881 48297 140915 48331
rect 157625 51765 157659 51799
rect 125977 46937 126011 46971
rect 133337 46869 133371 46903
rect 133337 37281 133371 37315
rect 150633 46869 150667 46903
rect 192125 56525 192159 56559
rect 179429 46937 179463 46971
rect 186237 55165 186271 55199
rect 157625 38641 157659 38675
rect 162961 46869 162995 46903
rect 150633 37281 150667 37315
rect 192125 46937 192159 46971
rect 207489 56525 207523 56559
rect 186237 45577 186271 45611
rect 192125 45849 192159 45883
rect 183753 45509 183787 45543
rect 162961 37281 162995 37315
rect 174001 40681 174035 40715
rect 140881 28917 140915 28951
rect 125977 27557 126011 27591
rect 133337 27557 133371 27591
rect 162961 27557 162995 27591
rect 140881 19397 140915 19431
rect 161765 22729 161799 22763
rect 133337 19261 133371 19295
rect 140881 19261 140915 19295
rect 125977 9673 126011 9707
rect 179429 37213 179463 37247
rect 179429 27625 179463 27659
rect 190653 45509 190687 45543
rect 192125 41293 192159 41327
rect 183753 27625 183787 27659
rect 186237 40681 186271 40715
rect 190653 40681 190687 40715
rect 290473 55233 290507 55267
rect 301789 57885 301823 57919
rect 280077 51017 280111 51051
rect 290381 51153 290415 51187
rect 271889 48161 271923 48195
rect 207489 38641 207523 38675
rect 214113 46869 214147 46903
rect 214113 37281 214147 37315
rect 215401 46869 215435 46903
rect 215401 37281 215435 37315
rect 248337 46869 248371 46903
rect 301789 48297 301823 48331
rect 322673 57885 322707 57919
rect 415041 66181 415075 66215
rect 325525 56593 325559 56627
rect 383209 57885 383243 57919
rect 322673 48297 322707 48331
rect 341533 51153 341567 51187
rect 290381 47005 290415 47039
rect 290657 46869 290691 46903
rect 271889 41293 271923 41327
rect 276121 46733 276155 46767
rect 248337 37281 248371 37315
rect 271889 38573 271923 38607
rect 244289 37213 244323 37247
rect 192217 31705 192251 31739
rect 244289 31637 244323 31671
rect 245761 37213 245795 37247
rect 245761 31637 245795 31671
rect 325709 46869 325743 46903
rect 290657 38505 290691 38539
rect 322673 38573 322707 38607
rect 276121 29053 276155 29087
rect 271889 28985 271923 29019
rect 383209 48297 383243 48331
rect 388729 57885 388763 57919
rect 388729 48297 388763 48331
rect 404001 57885 404035 57919
rect 415041 56593 415075 56627
rect 404001 48297 404035 48331
rect 341533 45577 341567 45611
rect 425989 46869 426023 46903
rect 414949 45509 414983 45543
rect 341441 45441 341475 45475
rect 341441 38233 341475 38267
rect 383209 38573 383243 38607
rect 325709 29053 325743 29087
rect 322673 28985 322707 29019
rect 383209 28985 383243 29019
rect 404001 38573 404035 38607
rect 425989 37281 426023 37315
rect 414949 35921 414983 35955
rect 431601 37213 431635 37247
rect 431601 31637 431635 31671
rect 404001 28985 404035 29019
rect 186237 27081 186271 27115
rect 190469 27557 190503 27591
rect 192217 27557 192251 27591
rect 207489 28917 207523 28951
rect 174001 26265 174035 26299
rect 183753 26197 183787 26231
rect 162961 17969 162995 18003
rect 179705 19261 179739 19295
rect 161765 11849 161799 11883
rect 168389 12461 168423 12495
rect 140881 9673 140915 9707
rect 168389 9673 168423 9707
rect 190469 17969 190503 18003
rect 192217 26197 192251 26231
rect 183753 16609 183787 16643
rect 279985 28917 280019 28951
rect 207489 19397 207523 19431
rect 214113 27557 214147 27591
rect 192217 16609 192251 16643
rect 207213 19261 207247 19295
rect 179705 9673 179739 9707
rect 207213 9673 207247 9707
rect 214113 9673 214147 9707
rect 215401 27557 215435 27591
rect 276121 27557 276155 27591
rect 222301 24905 222335 24939
rect 222301 23477 222335 23511
rect 230121 24769 230155 24803
rect 215401 9673 215435 9707
rect 227821 20009 227855 20043
rect 125609 8313 125643 8347
rect 123125 7361 123159 7395
rect 123125 7225 123159 7259
rect 125609 6953 125643 6987
rect 227821 6885 227855 6919
rect 238953 22185 238987 22219
rect 238953 19329 238987 19363
rect 238401 19261 238435 19295
rect 325709 27557 325743 27591
rect 279985 19329 280019 19363
rect 301881 26197 301915 26231
rect 276121 17969 276155 18003
rect 290933 19261 290967 19295
rect 238401 9673 238435 9707
rect 274833 15861 274867 15895
rect 274833 9673 274867 9707
rect 290933 9673 290967 9707
rect 420469 27557 420503 27591
rect 415041 26197 415075 26231
rect 383393 25245 383427 25279
rect 383393 19329 383427 19363
rect 420469 17969 420503 18003
rect 431509 26197 431543 26231
rect 415041 16609 415075 16643
rect 431509 16609 431543 16643
rect 325709 9673 325743 9707
rect 383301 12529 383335 12563
rect 383301 9673 383335 9707
rect 301881 8313 301915 8347
rect 414765 8245 414799 8279
rect 415041 8245 415075 8279
rect 412649 7565 412683 7599
rect 412649 7021 412683 7055
rect 230121 6885 230155 6919
rect 55229 4097 55263 4131
rect 55229 3145 55263 3179
rect 64797 4097 64831 4131
rect 64797 3145 64831 3179
rect 74549 4097 74583 4131
rect 74549 3145 74583 3179
rect 84117 4097 84151 4131
rect 84117 3145 84151 3179
rect 93869 4097 93903 4131
rect 93869 2941 93903 2975
rect 103437 4097 103471 4131
rect 103437 2941 103471 2975
rect 113189 4097 113223 4131
rect 113189 2873 113223 2907
rect 123493 4097 123527 4131
rect 123493 2873 123527 2907
rect 133153 4097 133187 4131
rect 133153 2873 133187 2907
rect 142813 4097 142847 4131
rect 148885 4097 148919 4131
rect 504557 4097 504591 4131
rect 149069 4029 149103 4063
rect 218069 4029 218103 4063
rect 355333 4029 355367 4063
rect 355517 4029 355551 4063
rect 217885 3825 217919 3859
rect 355241 3961 355275 3995
rect 229753 3893 229787 3927
rect 218069 3757 218103 3791
rect 225245 3825 225279 3859
rect 217885 3553 217919 3587
rect 217241 3485 217275 3519
rect 210065 3417 210099 3451
rect 194609 3281 194643 3315
rect 210065 3213 210099 3247
rect 225245 3349 225279 3383
rect 228833 3621 228867 3655
rect 326445 3757 326479 3791
rect 229753 3485 229787 3519
rect 234629 3553 234663 3587
rect 228833 3349 228867 3383
rect 234629 3349 234663 3383
rect 217241 3213 217275 3247
rect 194609 3145 194643 3179
rect 142813 2873 142847 2907
rect 340245 3689 340279 3723
rect 340245 3553 340279 3587
rect 398849 3825 398883 3859
rect 398849 3621 398883 3655
rect 407405 3757 407439 3791
rect 355241 3553 355275 3587
rect 407405 3485 407439 3519
rect 417985 3621 418019 3655
rect 427737 3553 427771 3587
rect 417985 3485 418019 3519
rect 418169 3485 418203 3519
rect 442273 3485 442307 3519
rect 418261 2941 418295 2975
rect 422309 2941 422343 2975
rect 427737 2941 427771 2975
rect 432521 3417 432555 3451
rect 422309 2737 422343 2771
rect 437397 3417 437431 3451
rect 437397 2941 437431 2975
rect 504373 3349 504407 3383
rect 482385 3281 482419 3315
rect 485697 3281 485731 3315
rect 480913 3213 480947 3247
rect 442273 2873 442307 2907
rect 463709 3009 463743 3043
rect 463709 2873 463743 2907
rect 473277 3009 473311 3043
rect 480913 3009 480947 3043
rect 481005 3213 481039 3247
rect 485145 3213 485179 3247
rect 481005 2941 481039 2975
rect 481097 2941 481131 2975
rect 482109 2941 482143 2975
rect 485053 2941 485087 2975
rect 485145 2941 485179 2975
rect 473277 2805 473311 2839
rect 489561 3281 489595 3315
rect 489101 3009 489135 3043
rect 489561 3009 489595 3043
rect 489653 3281 489687 3315
rect 496645 3281 496679 3315
rect 504557 3281 504591 3315
rect 504373 3213 504407 3247
rect 496645 3145 496679 3179
rect 485697 2873 485731 2907
rect 480821 2805 480855 2839
rect 483029 2805 483063 2839
rect 485053 2805 485087 2839
rect 432521 2737 432555 2771
rect 483029 2669 483063 2703
rect 326445 561 326479 595
<< metal1 >>
rect 133966 700952 133972 701004
rect 134024 700992 134030 701004
rect 267642 700992 267648 701004
rect 134024 700964 267648 700992
rect 134024 700952 134030 700964
rect 267642 700952 267648 700964
rect 267700 700952 267706 701004
rect 133782 700884 133788 700936
rect 133840 700924 133846 700936
rect 283834 700924 283840 700936
rect 133840 700896 283840 700924
rect 133840 700884 133846 700896
rect 283834 700884 283840 700896
rect 283892 700884 283898 700936
rect 300118 700884 300124 700936
rect 300176 700924 300182 700936
rect 434070 700924 434076 700936
rect 300176 700896 434076 700924
rect 300176 700884 300182 700896
rect 434070 700884 434076 700896
rect 434128 700884 434134 700936
rect 132494 700816 132500 700868
rect 132552 700856 132558 700868
rect 332502 700856 332508 700868
rect 132552 700828 332508 700856
rect 132552 700816 132558 700828
rect 332502 700816 332508 700828
rect 332560 700816 332566 700868
rect 133690 700748 133696 700800
rect 133748 700788 133754 700800
rect 218974 700788 218980 700800
rect 133748 700760 218980 700788
rect 133748 700748 133754 700760
rect 218974 700748 218980 700760
rect 219032 700748 219038 700800
rect 235166 700748 235172 700800
rect 235224 700788 235230 700800
rect 434162 700788 434168 700800
rect 235224 700760 434168 700788
rect 235224 700748 235230 700760
rect 434162 700748 434168 700760
rect 434220 700748 434226 700800
rect 131114 700680 131120 700732
rect 131172 700720 131178 700732
rect 348786 700720 348792 700732
rect 131172 700692 348792 700720
rect 131172 700680 131178 700692
rect 348786 700680 348792 700692
rect 348844 700680 348850 700732
rect 364978 700680 364984 700732
rect 365036 700720 365042 700732
rect 433978 700720 433984 700732
rect 365036 700692 433984 700720
rect 365036 700680 365042 700692
rect 433978 700680 433984 700692
rect 434036 700680 434042 700732
rect 170306 700612 170312 700664
rect 170364 700652 170370 700664
rect 434346 700652 434352 700664
rect 170364 700624 434352 700652
rect 170364 700612 170370 700624
rect 434346 700612 434352 700624
rect 434404 700612 434410 700664
rect 131206 700544 131212 700596
rect 131264 700584 131270 700596
rect 397454 700584 397460 700596
rect 131264 700556 397460 700584
rect 131264 700544 131270 700556
rect 397454 700544 397460 700556
rect 397512 700544 397518 700596
rect 132310 700476 132316 700528
rect 132368 700516 132374 700528
rect 413646 700516 413652 700528
rect 132368 700488 413652 700516
rect 132368 700476 132374 700488
rect 413646 700476 413652 700488
rect 413704 700476 413710 700528
rect 105446 700408 105452 700460
rect 105504 700448 105510 700460
rect 434438 700448 434444 700460
rect 105504 700420 434444 700448
rect 105504 700408 105510 700420
rect 434438 700408 434444 700420
rect 434496 700408 434502 700460
rect 438118 700408 438124 700460
rect 438176 700448 438182 700460
rect 494790 700448 494796 700460
rect 438176 700420 494796 700448
rect 438176 700408 438182 700420
rect 494790 700408 494796 700420
rect 494848 700408 494854 700460
rect 8110 700340 8116 700392
rect 8168 700380 8174 700392
rect 13078 700380 13084 700392
rect 8168 700352 13084 700380
rect 8168 700340 8174 700352
rect 13078 700340 13084 700352
rect 13136 700340 13142 700392
rect 89162 700340 89168 700392
rect 89220 700380 89226 700392
rect 126238 700380 126244 700392
rect 89220 700352 126244 700380
rect 89220 700340 89226 700352
rect 126238 700340 126244 700352
rect 126296 700340 126302 700392
rect 132586 700340 132592 700392
rect 132644 700380 132650 700392
rect 462314 700380 462320 700392
rect 132644 700352 462320 700380
rect 132644 700340 132650 700352
rect 462314 700340 462320 700352
rect 462372 700340 462378 700392
rect 40494 700272 40500 700324
rect 40552 700312 40558 700324
rect 434254 700312 434260 700324
rect 40552 700284 434260 700312
rect 40552 700272 40558 700284
rect 434254 700272 434260 700284
rect 434312 700272 434318 700324
rect 447778 700272 447784 700324
rect 447836 700312 447842 700324
rect 559650 700312 559656 700324
rect 447836 700284 559656 700312
rect 447836 700272 447842 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 133414 700204 133420 700256
rect 133472 700244 133478 700256
rect 202782 700244 202788 700256
rect 133472 700216 202788 700244
rect 133472 700204 133478 700216
rect 202782 700204 202788 700216
rect 202840 700204 202846 700256
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 72418 699660 72424 699712
rect 72476 699700 72482 699712
rect 72970 699700 72976 699712
rect 72476 699672 72976 699700
rect 72476 699660 72482 699672
rect 72970 699660 72976 699672
rect 73028 699660 73034 699712
rect 133322 699660 133328 699712
rect 133380 699700 133386 699712
rect 137830 699700 137836 699712
rect 133380 699672 137836 699700
rect 133380 699660 133386 699672
rect 137830 699660 137836 699672
rect 137888 699660 137894 699712
rect 429838 699660 429844 699712
rect 429896 699700 429902 699712
rect 433886 699700 433892 699712
rect 429896 699672 433892 699700
rect 429896 699660 429902 699672
rect 433886 699660 433892 699672
rect 433944 699660 433950 699712
rect 153562 698232 153568 698284
rect 153620 698272 153626 698284
rect 154206 698272 154212 698284
rect 153620 698244 154212 698272
rect 153620 698232 153626 698244
rect 154206 698232 154212 698244
rect 154264 698232 154270 698284
rect 147582 697076 147588 697128
rect 147640 697116 147646 697128
rect 154482 697116 154488 697128
rect 147640 697088 154488 697116
rect 147640 697076 147646 697088
rect 154482 697076 154488 697088
rect 154540 697076 154546 697128
rect 166902 697076 166908 697128
rect 166960 697116 166966 697128
rect 173802 697116 173808 697128
rect 166960 697088 173808 697116
rect 166960 697076 166966 697088
rect 173802 697076 173808 697088
rect 173860 697076 173866 697128
rect 186222 697076 186228 697128
rect 186280 697116 186286 697128
rect 193122 697116 193128 697128
rect 186280 697088 193128 697116
rect 186280 697076 186286 697088
rect 193122 697076 193128 697088
rect 193180 697076 193186 697128
rect 205542 697076 205548 697128
rect 205600 697116 205606 697128
rect 212442 697116 212448 697128
rect 205600 697088 212448 697116
rect 205600 697076 205606 697088
rect 212442 697076 212448 697088
rect 212500 697076 212506 697128
rect 224862 697076 224868 697128
rect 224920 697116 224926 697128
rect 231762 697116 231768 697128
rect 224920 697088 231768 697116
rect 224920 697076 224926 697088
rect 231762 697076 231768 697088
rect 231820 697076 231826 697128
rect 244182 697076 244188 697128
rect 244240 697116 244246 697128
rect 251082 697116 251088 697128
rect 244240 697088 251088 697116
rect 244240 697076 244246 697088
rect 251082 697076 251088 697088
rect 251140 697076 251146 697128
rect 263502 697076 263508 697128
rect 263560 697116 263566 697128
rect 270402 697116 270408 697128
rect 263560 697088 270408 697116
rect 263560 697076 263566 697088
rect 270402 697076 270408 697088
rect 270460 697076 270466 697128
rect 282822 697076 282828 697128
rect 282880 697116 282886 697128
rect 289722 697116 289728 697128
rect 282880 697088 289728 697116
rect 282880 697076 282886 697088
rect 289722 697076 289728 697088
rect 289780 697076 289786 697128
rect 302142 697076 302148 697128
rect 302200 697116 302206 697128
rect 309042 697116 309048 697128
rect 302200 697088 309048 697116
rect 302200 697076 302206 697088
rect 309042 697076 309048 697088
rect 309100 697076 309106 697128
rect 321462 697076 321468 697128
rect 321520 697116 321526 697128
rect 328362 697116 328368 697128
rect 321520 697088 328368 697116
rect 321520 697076 321526 697088
rect 328362 697076 328368 697088
rect 328420 697076 328426 697128
rect 154574 686264 154580 686316
rect 154632 686304 154638 686316
rect 159450 686304 159456 686316
rect 154632 686276 159456 686304
rect 154632 686264 154638 686276
rect 159450 686264 159456 686276
rect 159508 686264 159514 686316
rect 135254 686128 135260 686180
rect 135312 686168 135318 686180
rect 142890 686168 142896 686180
rect 135312 686140 142896 686168
rect 135312 686128 135318 686140
rect 142890 686128 142896 686140
rect 142948 686128 142954 686180
rect 153286 685924 153292 685976
rect 153344 685964 153350 685976
rect 153654 685964 153660 685976
rect 153344 685936 153660 685964
rect 153344 685924 153350 685936
rect 153654 685924 153660 685936
rect 153712 685924 153718 685976
rect 153286 684428 153292 684480
rect 153344 684468 153350 684480
rect 153565 684471 153623 684477
rect 153565 684468 153577 684471
rect 153344 684440 153577 684468
rect 153344 684428 153350 684440
rect 153565 684437 153577 684440
rect 153611 684437 153623 684471
rect 153565 684431 153623 684437
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 434714 681748 434720 681760
rect 3568 681720 434720 681748
rect 3568 681708 3574 681720
rect 434714 681708 434720 681720
rect 434772 681708 434778 681760
rect 446398 673480 446404 673532
rect 446456 673520 446462 673532
rect 580166 673520 580172 673532
rect 446456 673492 580172 673520
rect 446456 673480 446462 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 19978 667944 19984 667956
rect 3476 667916 19984 667944
rect 3476 667904 3482 667916
rect 19978 667904 19984 667916
rect 20036 667904 20042 667956
rect 153565 666587 153623 666593
rect 153565 666553 153577 666587
rect 153611 666584 153623 666587
rect 153654 666584 153660 666596
rect 153611 666556 153660 666584
rect 153611 666553 153623 666556
rect 153565 666547 153623 666553
rect 153654 666544 153660 666556
rect 153712 666544 153718 666596
rect 153470 656860 153476 656872
rect 153431 656832 153476 656860
rect 153470 656820 153476 656832
rect 153528 656820 153534 656872
rect 154574 650360 154580 650412
rect 154632 650400 154638 650412
rect 159450 650400 159456 650412
rect 154632 650372 159456 650400
rect 154632 650360 154638 650372
rect 159450 650360 159456 650372
rect 159508 650360 159514 650412
rect 135254 650224 135260 650276
rect 135312 650264 135318 650276
rect 142890 650264 142896 650276
rect 135312 650236 142896 650264
rect 135312 650224 135318 650236
rect 142890 650224 142896 650236
rect 142948 650224 142954 650276
rect 153473 647275 153531 647281
rect 153473 647241 153485 647275
rect 153519 647272 153531 647275
rect 153562 647272 153568 647284
rect 153519 647244 153568 647272
rect 153519 647241 153531 647244
rect 153473 647235 153531 647241
rect 153562 647232 153568 647244
rect 153620 647232 153626 647284
rect 153286 637644 153292 637696
rect 153344 637684 153350 637696
rect 153562 637684 153568 637696
rect 153344 637656 153568 637684
rect 153344 637644 153350 637656
rect 153562 637644 153568 637656
rect 153620 637644 153626 637696
rect 153378 630708 153384 630760
rect 153436 630708 153442 630760
rect 153396 630544 153424 630708
rect 153562 630544 153568 630556
rect 153396 630516 153568 630544
rect 153562 630504 153568 630516
rect 153620 630504 153626 630556
rect 445018 626560 445024 626612
rect 445076 626600 445082 626612
rect 580166 626600 580172 626612
rect 445076 626572 580172 626600
rect 445076 626560 445082 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 153562 626492 153568 626544
rect 153620 626532 153626 626544
rect 153746 626532 153752 626544
rect 153620 626504 153752 626532
rect 153620 626492 153626 626504
rect 153746 626492 153752 626504
rect 153804 626492 153810 626544
rect 3418 623772 3424 623824
rect 3476 623812 3482 623824
rect 434806 623812 434812 623824
rect 3476 623784 434812 623812
rect 3476 623772 3482 623784
rect 434806 623772 434812 623784
rect 434864 623772 434870 623824
rect 153562 611192 153568 611244
rect 153620 611232 153626 611244
rect 153746 611232 153752 611244
rect 153620 611204 153752 611232
rect 153620 611192 153626 611204
rect 153746 611192 153752 611204
rect 153804 611192 153810 611244
rect 3418 609968 3424 610020
rect 3476 610008 3482 610020
rect 21358 610008 21364 610020
rect 3476 609980 21364 610008
rect 3476 609968 3482 609980
rect 21358 609968 21364 609980
rect 21416 609968 21422 610020
rect 153378 598952 153384 599004
rect 153436 598992 153442 599004
rect 153562 598992 153568 599004
rect 153436 598964 153568 598992
rect 153436 598952 153442 598964
rect 153562 598952 153568 598964
rect 153620 598952 153626 599004
rect 4062 594804 4068 594856
rect 4120 594844 4126 594856
rect 4890 594844 4896 594856
rect 4120 594816 4896 594844
rect 4120 594804 4126 594816
rect 4890 594804 4896 594816
rect 4948 594804 4954 594856
rect 153286 591948 153292 592000
rect 153344 591988 153350 592000
rect 153562 591988 153568 592000
rect 153344 591960 153568 591988
rect 153344 591948 153350 591960
rect 153562 591948 153568 591960
rect 153620 591948 153626 592000
rect 175918 583652 175924 583704
rect 175976 583692 175982 583704
rect 302786 583692 302792 583704
rect 175976 583664 302792 583692
rect 175976 583652 175982 583664
rect 302786 583652 302792 583664
rect 302844 583652 302850 583704
rect 270402 583584 270408 583636
rect 270460 583624 270466 583636
rect 307018 583624 307024 583636
rect 270460 583596 307024 583624
rect 270460 583584 270466 583596
rect 307018 583584 307024 583596
rect 307076 583584 307082 583636
rect 286318 583516 286324 583568
rect 286376 583556 286382 583568
rect 319714 583556 319720 583568
rect 286376 583528 319720 583556
rect 286376 583516 286382 583528
rect 319714 583516 319720 583528
rect 319772 583516 319778 583568
rect 129274 583448 129280 583500
rect 129332 583488 129338 583500
rect 347498 583488 347504 583500
rect 129332 583460 347504 583488
rect 129332 583448 129338 583460
rect 347498 583448 347504 583460
rect 347556 583448 347562 583500
rect 126330 583380 126336 583432
rect 126388 583420 126394 583432
rect 324130 583420 324136 583432
rect 126388 583392 324136 583420
rect 126388 583380 126394 583392
rect 324130 583380 324136 583392
rect 324188 583380 324194 583432
rect 85390 583312 85396 583364
rect 85448 583352 85454 583364
rect 334618 583352 334624 583364
rect 85448 583324 334624 583352
rect 85448 583312 85454 583324
rect 334618 583312 334624 583324
rect 334676 583312 334682 583364
rect 85574 583244 85580 583296
rect 85632 583284 85638 583296
rect 345290 583284 345296 583296
rect 85632 583256 345296 583284
rect 85632 583244 85638 583256
rect 345290 583244 345296 583256
rect 345348 583244 345354 583296
rect 291838 583176 291844 583228
rect 291896 583216 291902 583228
rect 328362 583216 328368 583228
rect 291896 583188 328368 583216
rect 291896 583176 291902 583188
rect 328362 583176 328368 583188
rect 328420 583176 328426 583228
rect 298922 583108 298928 583160
rect 298980 583148 298986 583160
rect 341058 583148 341064 583160
rect 298980 583120 341064 583148
rect 298980 583108 298986 583120
rect 341058 583108 341064 583120
rect 341116 583108 341122 583160
rect 294598 583040 294604 583092
rect 294656 583080 294662 583092
rect 338850 583080 338856 583092
rect 294656 583052 338856 583080
rect 294656 583040 294662 583052
rect 338850 583040 338856 583052
rect 338908 583040 338914 583092
rect 281350 582972 281356 583024
rect 281408 583012 281414 583024
rect 326154 583012 326160 583024
rect 281408 582984 326160 583012
rect 281408 582972 281414 582984
rect 326154 582972 326160 582984
rect 326212 582972 326218 583024
rect 299014 582904 299020 582956
rect 299072 582944 299078 582956
rect 353754 582944 353760 582956
rect 299072 582916 353760 582944
rect 299072 582904 299078 582916
rect 353754 582904 353760 582916
rect 353812 582904 353818 582956
rect 298646 582836 298652 582888
rect 298704 582876 298710 582888
rect 355962 582876 355968 582888
rect 298704 582848 355968 582876
rect 298704 582836 298710 582848
rect 355962 582836 355968 582848
rect 356020 582836 356026 582888
rect 291102 582768 291108 582820
rect 291160 582808 291166 582820
rect 351730 582808 351736 582820
rect 291160 582780 351736 582808
rect 291160 582768 291166 582780
rect 351730 582768 351736 582780
rect 351788 582768 351794 582820
rect 298738 582700 298744 582752
rect 298796 582740 298802 582752
rect 360194 582740 360200 582752
rect 298796 582712 360200 582740
rect 298796 582700 298802 582712
rect 360194 582700 360200 582712
rect 360252 582700 360258 582752
rect 300486 582632 300492 582684
rect 300544 582672 300550 582684
rect 362402 582672 362408 582684
rect 300544 582644 362408 582672
rect 300544 582632 300550 582644
rect 362402 582632 362408 582644
rect 362460 582632 362466 582684
rect 366634 582632 366640 582684
rect 366692 582672 366698 582684
rect 378870 582672 378876 582684
rect 366692 582644 378876 582672
rect 366692 582632 366698 582644
rect 378870 582632 378876 582644
rect 378928 582632 378934 582684
rect 298830 582564 298836 582616
rect 298888 582604 298894 582616
rect 332594 582604 332600 582616
rect 298888 582576 332600 582604
rect 298888 582564 298894 582576
rect 332594 582564 332600 582576
rect 332652 582564 332658 582616
rect 357986 582564 357992 582616
rect 358044 582604 358050 582616
rect 378410 582604 378416 582616
rect 358044 582576 378416 582604
rect 358044 582564 358050 582576
rect 378410 582564 378416 582576
rect 378468 582564 378474 582616
rect 298462 582496 298468 582548
rect 298520 582536 298526 582548
rect 321922 582536 321928 582548
rect 298520 582508 321928 582536
rect 298520 582496 298526 582508
rect 321922 582496 321928 582508
rect 321980 582496 321986 582548
rect 370866 582496 370872 582548
rect 370924 582536 370930 582548
rect 378686 582536 378692 582548
rect 370924 582508 378692 582536
rect 370924 582496 370930 582508
rect 378686 582496 378692 582508
rect 378744 582496 378750 582548
rect 287698 582428 287704 582480
rect 287756 582468 287762 582480
rect 313458 582468 313464 582480
rect 287756 582440 313464 582468
rect 287756 582428 287762 582440
rect 313458 582428 313464 582440
rect 313516 582428 313522 582480
rect 298554 582360 298560 582412
rect 298612 582400 298618 582412
rect 309226 582400 309232 582412
rect 298612 582372 309232 582400
rect 298612 582360 298618 582372
rect 309226 582360 309232 582372
rect 309284 582360 309290 582412
rect 372890 582360 372896 582412
rect 372948 582400 372954 582412
rect 378594 582400 378600 582412
rect 372948 582372 378600 582400
rect 372948 582360 372954 582372
rect 378594 582360 378600 582372
rect 378652 582360 378658 582412
rect 299382 579640 299388 579692
rect 299440 579680 299446 579692
rect 304810 579680 304816 579692
rect 299440 579652 304816 579680
rect 299440 579640 299446 579652
rect 304810 579640 304816 579652
rect 304868 579640 304874 579692
rect 442258 579640 442264 579692
rect 442316 579680 442322 579692
rect 580166 579680 580172 579692
rect 442316 579652 580172 579680
rect 442316 579640 442322 579652
rect 580166 579640 580172 579652
rect 580224 579640 580230 579692
rect 153378 579612 153384 579624
rect 153339 579584 153384 579612
rect 153378 579572 153384 579584
rect 153436 579572 153442 579624
rect 299474 579300 299480 579352
rect 299532 579340 299538 579352
rect 300670 579340 300676 579352
rect 299532 579312 300676 579340
rect 299532 579300 299538 579312
rect 300670 579300 300676 579312
rect 300728 579300 300734 579352
rect 310974 579340 310980 579352
rect 310935 579312 310980 579340
rect 310974 579300 310980 579312
rect 311032 579300 311038 579352
rect 315206 579340 315212 579352
rect 315167 579312 315212 579340
rect 315206 579300 315212 579312
rect 315264 579300 315270 579352
rect 317414 579340 317420 579352
rect 317375 579312 317420 579340
rect 317414 579300 317420 579312
rect 317472 579300 317478 579352
rect 330202 579300 330208 579352
rect 330260 579300 330266 579352
rect 336642 579340 336648 579352
rect 336603 579312 336648 579340
rect 336642 579300 336648 579312
rect 336700 579300 336706 579352
rect 342990 579340 342996 579352
rect 342951 579312 342996 579340
rect 342990 579300 342996 579312
rect 343048 579300 343054 579352
rect 364242 579340 364248 579352
rect 364203 579312 364248 579340
rect 364242 579300 364248 579312
rect 364300 579300 364306 579352
rect 375374 579300 375380 579352
rect 375432 579340 375438 579352
rect 378502 579340 378508 579352
rect 375432 579312 378508 579340
rect 375432 579300 375438 579312
rect 378502 579300 378508 579312
rect 378560 579300 378566 579352
rect 183557 578935 183615 578941
rect 183557 578901 183569 578935
rect 183603 578932 183615 578935
rect 193125 578935 193183 578941
rect 193125 578932 193137 578935
rect 183603 578904 193137 578932
rect 183603 578901 183615 578904
rect 183557 578895 183615 578901
rect 193125 578901 193137 578904
rect 193171 578901 193183 578935
rect 193125 578895 193183 578901
rect 202877 578935 202935 578941
rect 202877 578901 202889 578935
rect 202923 578932 202935 578935
rect 212445 578935 212503 578941
rect 212445 578932 212457 578935
rect 202923 578904 212457 578932
rect 202923 578901 202935 578904
rect 202877 578895 202935 578901
rect 212445 578901 212457 578904
rect 212491 578901 212503 578935
rect 212445 578895 212503 578901
rect 222197 578935 222255 578941
rect 222197 578901 222209 578935
rect 222243 578932 222255 578935
rect 231765 578935 231823 578941
rect 231765 578932 231777 578935
rect 222243 578904 231777 578932
rect 222243 578901 222255 578904
rect 222197 578895 222255 578901
rect 231765 578901 231777 578904
rect 231811 578901 231823 578935
rect 231765 578895 231823 578901
rect 241517 578935 241575 578941
rect 241517 578901 241529 578935
rect 241563 578932 241575 578935
rect 251085 578935 251143 578941
rect 251085 578932 251097 578935
rect 241563 578904 251097 578932
rect 241563 578901 241575 578904
rect 241517 578895 241575 578901
rect 251085 578901 251097 578904
rect 251131 578901 251143 578935
rect 251085 578895 251143 578901
rect 270497 578935 270555 578941
rect 270497 578901 270509 578935
rect 270543 578932 270555 578935
rect 282825 578935 282883 578941
rect 282825 578932 282837 578935
rect 270543 578904 282837 578932
rect 270543 578901 270555 578904
rect 270497 578895 270555 578901
rect 282825 578901 282837 578904
rect 282871 578901 282883 578935
rect 282825 578895 282883 578901
rect 282917 578935 282975 578941
rect 282917 578901 282929 578935
rect 282963 578932 282975 578935
rect 292485 578935 292543 578941
rect 292485 578932 292497 578935
rect 282963 578904 292497 578932
rect 282963 578901 282975 578904
rect 282917 578895 282975 578901
rect 292485 578901 292497 578904
rect 292531 578901 292543 578935
rect 292485 578895 292543 578901
rect 318797 578935 318855 578941
rect 318797 578901 318809 578935
rect 318843 578932 318855 578935
rect 323581 578935 323639 578941
rect 323581 578932 323593 578935
rect 318843 578904 323593 578932
rect 318843 578901 318855 578904
rect 318797 578895 318855 578901
rect 323581 578901 323593 578904
rect 323627 578901 323639 578935
rect 323581 578895 323639 578901
rect 154577 578867 154635 578873
rect 154577 578833 154589 578867
rect 154623 578864 154635 578867
rect 164145 578867 164203 578873
rect 164145 578864 164157 578867
rect 154623 578836 164157 578864
rect 154623 578833 154635 578836
rect 154577 578827 154635 578833
rect 164145 578833 164157 578836
rect 164191 578833 164203 578867
rect 270405 578867 270463 578873
rect 270405 578864 270417 578867
rect 164145 578827 164203 578833
rect 263428 578836 270417 578864
rect 128998 578756 129004 578808
rect 129056 578796 129062 578808
rect 142801 578799 142859 578805
rect 142801 578796 142813 578799
rect 129056 578768 142813 578796
rect 129056 578756 129062 578768
rect 142801 578765 142813 578768
rect 142847 578765 142859 578799
rect 176565 578799 176623 578805
rect 176565 578796 176577 578799
rect 142801 578759 142859 578765
rect 166920 578768 176577 578796
rect 130378 578688 130384 578740
rect 130436 578728 130442 578740
rect 154577 578731 154635 578737
rect 154577 578728 154589 578731
rect 130436 578700 154589 578728
rect 130436 578688 130442 578700
rect 154577 578697 154589 578700
rect 154623 578697 154635 578731
rect 154577 578691 154635 578697
rect 164145 578731 164203 578737
rect 164145 578697 164157 578731
rect 164191 578728 164203 578731
rect 166920 578728 166948 578768
rect 176565 578765 176577 578768
rect 176611 578765 176623 578799
rect 176565 578759 176623 578765
rect 176657 578799 176715 578805
rect 176657 578765 176669 578799
rect 176703 578796 176715 578799
rect 193125 578799 193183 578805
rect 176703 578768 178632 578796
rect 176703 578765 176715 578768
rect 176657 578759 176715 578765
rect 164191 578700 166948 578728
rect 178604 578728 178632 578768
rect 193125 578765 193137 578799
rect 193171 578796 193183 578799
rect 195885 578799 195943 578805
rect 195885 578796 195897 578799
rect 193171 578768 195897 578796
rect 193171 578765 193183 578768
rect 193125 578759 193183 578765
rect 195885 578765 195897 578768
rect 195931 578765 195943 578799
rect 195885 578759 195943 578765
rect 212445 578799 212503 578805
rect 212445 578765 212457 578799
rect 212491 578796 212503 578799
rect 215205 578799 215263 578805
rect 215205 578796 215217 578799
rect 212491 578768 215217 578796
rect 212491 578765 212503 578768
rect 212445 578759 212503 578765
rect 215205 578765 215217 578768
rect 215251 578765 215263 578799
rect 215205 578759 215263 578765
rect 231765 578799 231823 578805
rect 231765 578765 231777 578799
rect 231811 578796 231823 578799
rect 234525 578799 234583 578805
rect 234525 578796 234537 578799
rect 231811 578768 234537 578796
rect 231811 578765 231823 578768
rect 231765 578759 231823 578765
rect 234525 578765 234537 578768
rect 234571 578765 234583 578799
rect 234525 578759 234583 578765
rect 251085 578799 251143 578805
rect 251085 578765 251097 578799
rect 251131 578796 251143 578799
rect 253845 578799 253903 578805
rect 253845 578796 253857 578799
rect 251131 578768 253857 578796
rect 251131 578765 251143 578768
rect 251085 578759 251143 578765
rect 253845 578765 253857 578768
rect 253891 578765 253903 578799
rect 253845 578759 253903 578765
rect 183557 578731 183615 578737
rect 183557 578728 183569 578731
rect 178604 578700 183569 578728
rect 164191 578697 164203 578700
rect 164145 578691 164203 578697
rect 183557 578697 183569 578700
rect 183603 578697 183615 578731
rect 183557 578691 183615 578697
rect 196069 578731 196127 578737
rect 196069 578697 196081 578731
rect 196115 578728 196127 578731
rect 202877 578731 202935 578737
rect 202877 578728 202889 578731
rect 196115 578700 202889 578728
rect 196115 578697 196127 578700
rect 196069 578691 196127 578697
rect 202877 578697 202889 578700
rect 202923 578697 202935 578731
rect 202877 578691 202935 578697
rect 215389 578731 215447 578737
rect 215389 578697 215401 578731
rect 215435 578728 215447 578731
rect 222197 578731 222255 578737
rect 222197 578728 222209 578731
rect 215435 578700 222209 578728
rect 215435 578697 215447 578700
rect 215389 578691 215447 578697
rect 222197 578697 222209 578700
rect 222243 578697 222255 578731
rect 222197 578691 222255 578697
rect 234709 578731 234767 578737
rect 234709 578697 234721 578731
rect 234755 578728 234767 578731
rect 241517 578731 241575 578737
rect 241517 578728 241529 578731
rect 234755 578700 241529 578728
rect 234755 578697 234767 578700
rect 234709 578691 234767 578697
rect 241517 578697 241529 578700
rect 241563 578697 241575 578731
rect 241517 578691 241575 578697
rect 254029 578731 254087 578737
rect 254029 578697 254041 578731
rect 254075 578728 254087 578731
rect 263428 578728 263456 578836
rect 270405 578833 270417 578836
rect 270451 578833 270463 578867
rect 270405 578827 270463 578833
rect 268381 578799 268439 578805
rect 268381 578765 268393 578799
rect 268427 578796 268439 578799
rect 278041 578799 278099 578805
rect 278041 578796 278053 578799
rect 268427 578768 278053 578796
rect 268427 578765 268439 578768
rect 268381 578759 268439 578765
rect 278041 578765 278053 578768
rect 278087 578765 278099 578799
rect 278041 578759 278099 578765
rect 284113 578799 284171 578805
rect 284113 578765 284125 578799
rect 284159 578796 284171 578799
rect 294417 578799 294475 578805
rect 294417 578796 294429 578799
rect 284159 578768 294429 578796
rect 284159 578765 284171 578768
rect 284113 578759 284171 578765
rect 294417 578765 294429 578768
rect 294463 578765 294475 578799
rect 294417 578759 294475 578765
rect 311989 578799 312047 578805
rect 311989 578765 312001 578799
rect 312035 578796 312047 578799
rect 318797 578799 318855 578805
rect 318797 578796 318809 578799
rect 312035 578768 318809 578796
rect 312035 578765 312047 578768
rect 311989 578759 312047 578765
rect 318797 578765 318809 578768
rect 318843 578765 318855 578799
rect 318797 578759 318855 578765
rect 323581 578799 323639 578805
rect 323581 578765 323593 578799
rect 323627 578796 323639 578799
rect 330220 578796 330248 579300
rect 323627 578768 330248 578796
rect 323627 578765 323639 578768
rect 323581 578759 323639 578765
rect 254075 578700 263456 578728
rect 306377 578731 306435 578737
rect 254075 578697 254087 578700
rect 254029 578691 254087 578697
rect 306377 578697 306389 578731
rect 306423 578728 306435 578731
rect 311805 578731 311863 578737
rect 311805 578728 311817 578731
rect 306423 578700 311817 578728
rect 306423 578697 306435 578700
rect 306377 578691 306435 578697
rect 311805 578697 311817 578700
rect 311851 578697 311863 578731
rect 311805 578691 311863 578697
rect 270405 578663 270463 578669
rect 270405 578629 270417 578663
rect 270451 578660 270463 578663
rect 270497 578663 270555 578669
rect 270497 578660 270509 578663
rect 270451 578632 270509 578660
rect 270451 578629 270463 578632
rect 270405 578623 270463 578629
rect 270497 578629 270509 578632
rect 270543 578629 270555 578663
rect 270497 578623 270555 578629
rect 292485 578663 292543 578669
rect 292485 578629 292497 578663
rect 292531 578660 292543 578663
rect 310977 578663 311035 578669
rect 310977 578660 310989 578663
rect 292531 578632 310989 578660
rect 292531 578629 292543 578632
rect 292485 578623 292543 578629
rect 310977 578629 310989 578632
rect 311023 578629 311035 578663
rect 310977 578623 311035 578629
rect 122742 578552 122748 578604
rect 122800 578592 122806 578604
rect 315209 578595 315267 578601
rect 315209 578592 315221 578595
rect 122800 578564 315221 578592
rect 122800 578552 122806 578564
rect 315209 578561 315221 578564
rect 315255 578561 315267 578595
rect 315209 578555 315267 578561
rect 142801 578527 142859 578533
rect 142801 578493 142813 578527
rect 142847 578524 142859 578527
rect 268381 578527 268439 578533
rect 268381 578524 268393 578527
rect 142847 578496 268393 578524
rect 142847 578493 142859 578496
rect 142801 578487 142859 578493
rect 268381 578493 268393 578496
rect 268427 578493 268439 578527
rect 268381 578487 268439 578493
rect 278041 578527 278099 578533
rect 278041 578493 278053 578527
rect 278087 578524 278099 578527
rect 284113 578527 284171 578533
rect 284113 578524 284125 578527
rect 278087 578496 284125 578524
rect 278087 578493 278099 578496
rect 278041 578487 278099 578493
rect 284113 578493 284125 578496
rect 284159 578493 284171 578527
rect 284113 578487 284171 578493
rect 294417 578527 294475 578533
rect 294417 578493 294429 578527
rect 294463 578524 294475 578527
rect 306377 578527 306435 578533
rect 306377 578524 306389 578527
rect 294463 578496 306389 578524
rect 294463 578493 294475 578496
rect 294417 578487 294475 578493
rect 306377 578493 306389 578496
rect 306423 578493 306435 578527
rect 306377 578487 306435 578493
rect 115382 578416 115388 578468
rect 115440 578456 115446 578468
rect 317417 578459 317475 578465
rect 317417 578456 317429 578459
rect 115440 578428 317429 578456
rect 115440 578416 115446 578428
rect 317417 578425 317429 578428
rect 317463 578425 317475 578459
rect 317417 578419 317475 578425
rect 119338 578348 119344 578400
rect 119396 578388 119402 578400
rect 336645 578391 336703 578397
rect 336645 578388 336657 578391
rect 119396 578360 336657 578388
rect 119396 578348 119402 578360
rect 336645 578357 336657 578360
rect 336691 578357 336703 578391
rect 336645 578351 336703 578357
rect 115198 578280 115204 578332
rect 115256 578320 115262 578332
rect 342993 578323 343051 578329
rect 342993 578320 343005 578323
rect 115256 578292 343005 578320
rect 115256 578280 115262 578292
rect 342993 578289 343005 578292
rect 343039 578289 343051 578323
rect 342993 578283 343051 578289
rect 129182 578212 129188 578264
rect 129240 578252 129246 578264
rect 364245 578255 364303 578261
rect 364245 578252 364257 578255
rect 129240 578224 364257 578252
rect 129240 578212 129246 578224
rect 364245 578221 364257 578224
rect 364291 578221 364303 578255
rect 364245 578215 364303 578221
rect 110322 575492 110328 575544
rect 110380 575532 110386 575544
rect 296714 575532 296720 575544
rect 110380 575504 296720 575532
rect 110380 575492 110386 575504
rect 296714 575492 296720 575504
rect 296772 575492 296778 575544
rect 153381 569959 153439 569965
rect 153381 569925 153393 569959
rect 153427 569956 153439 569959
rect 153470 569956 153476 569968
rect 153427 569928 153476 569956
rect 153427 569925 153439 569928
rect 153381 569919 153439 569925
rect 153470 569916 153476 569928
rect 153528 569916 153534 569968
rect 272518 569916 272524 569968
rect 272576 569956 272582 569968
rect 298002 569956 298008 569968
rect 272576 569928 298008 569956
rect 272576 569916 272582 569928
rect 298002 569916 298008 569928
rect 298060 569916 298066 569968
rect 153289 563159 153347 563165
rect 153289 563125 153301 563159
rect 153335 563156 153347 563159
rect 153470 563156 153476 563168
rect 153335 563128 153476 563156
rect 153335 563125 153347 563128
rect 153289 563119 153347 563125
rect 153470 563116 153476 563128
rect 153528 563116 153534 563168
rect 129550 563048 129556 563100
rect 129608 563088 129614 563100
rect 296898 563088 296904 563100
rect 129608 563060 296904 563088
rect 129608 563048 129614 563060
rect 296898 563048 296904 563060
rect 296956 563048 296962 563100
rect 153286 563020 153292 563032
rect 153247 562992 153292 563020
rect 153286 562980 153292 562992
rect 153344 562980 153350 563032
rect 200117 562139 200175 562145
rect 200117 562105 200129 562139
rect 200163 562136 200175 562139
rect 208765 562139 208823 562145
rect 208765 562136 208777 562139
rect 200163 562108 208777 562136
rect 200163 562105 200175 562108
rect 200117 562099 200175 562105
rect 208765 562105 208777 562108
rect 208811 562105 208823 562139
rect 208765 562099 208823 562105
rect 195882 561960 195888 562012
rect 195940 562000 195946 562012
rect 200117 562003 200175 562009
rect 200117 562000 200129 562003
rect 195940 561972 200129 562000
rect 195940 561960 195946 561972
rect 200117 561969 200129 561972
rect 200163 561969 200175 562003
rect 200117 561963 200175 561969
rect 197078 561892 197084 561944
rect 197136 561932 197142 561944
rect 208670 561932 208676 561944
rect 197136 561904 208676 561932
rect 197136 561892 197142 561904
rect 208670 561892 208676 561904
rect 208728 561892 208734 561944
rect 208765 561935 208823 561941
rect 208765 561901 208777 561935
rect 208811 561932 208823 561935
rect 217870 561932 217876 561944
rect 208811 561904 217876 561932
rect 208811 561901 208823 561904
rect 208765 561895 208823 561901
rect 217870 561892 217876 561904
rect 217928 561892 217934 561944
rect 196986 561824 196992 561876
rect 197044 561864 197050 561876
rect 205542 561864 205548 561876
rect 197044 561836 205548 561864
rect 197044 561824 197050 561836
rect 205542 561824 205548 561836
rect 205600 561824 205606 561876
rect 197262 561756 197268 561808
rect 197320 561796 197326 561808
rect 214742 561796 214748 561808
rect 197320 561768 214748 561796
rect 197320 561756 197326 561768
rect 214742 561756 214748 561768
rect 214800 561756 214806 561808
rect 153286 560232 153292 560244
rect 153247 560204 153292 560232
rect 153286 560192 153292 560204
rect 153344 560192 153350 560244
rect 197170 560192 197176 560244
rect 197228 560232 197234 560244
rect 202046 560232 202052 560244
rect 197228 560204 202052 560232
rect 197228 560192 197234 560204
rect 202046 560192 202052 560204
rect 202104 560192 202110 560244
rect 420178 556248 420184 556300
rect 420236 556288 420242 556300
rect 511258 556288 511264 556300
rect 420236 556260 511264 556288
rect 420236 556248 420242 556260
rect 511258 556248 511264 556260
rect 511316 556248 511322 556300
rect 273162 556180 273168 556232
rect 273220 556220 273226 556232
rect 297082 556220 297088 556232
rect 273220 556192 297088 556220
rect 273220 556180 273226 556192
rect 297082 556180 297088 556192
rect 297140 556180 297146 556232
rect 378778 556180 378784 556232
rect 378836 556220 378842 556232
rect 484394 556220 484400 556232
rect 378836 556192 484400 556220
rect 378836 556180 378842 556192
rect 484394 556180 484400 556192
rect 484452 556180 484458 556232
rect 109402 554752 109408 554804
rect 109460 554792 109466 554804
rect 110322 554792 110328 554804
rect 109460 554764 110328 554792
rect 109460 554752 109466 554764
rect 110322 554752 110328 554764
rect 110380 554792 110386 554804
rect 115934 554792 115940 554804
rect 110380 554764 115940 554792
rect 110380 554752 110386 554764
rect 115934 554752 115940 554764
rect 115992 554752 115998 554804
rect 92106 553936 92112 553988
rect 92164 553976 92170 553988
rect 115290 553976 115296 553988
rect 92164 553948 115296 553976
rect 92164 553936 92170 553948
rect 115290 553936 115296 553948
rect 115348 553936 115354 553988
rect 89162 553868 89168 553920
rect 89220 553908 89226 553920
rect 162118 553908 162124 553920
rect 89220 553880 162124 553908
rect 89220 553868 89226 553880
rect 162118 553868 162124 553880
rect 162176 553868 162182 553920
rect 115106 553800 115112 553852
rect 115164 553840 115170 553852
rect 128354 553840 128360 553852
rect 115164 553812 128360 553840
rect 115164 553800 115170 553812
rect 128354 553800 128360 553812
rect 128412 553840 128418 553852
rect 129274 553840 129280 553852
rect 128412 553812 129280 553840
rect 128412 553800 128418 553812
rect 129274 553800 129280 553812
rect 129332 553800 129338 553852
rect 95050 553732 95056 553784
rect 95108 553772 95114 553784
rect 120718 553772 120724 553784
rect 95108 553744 120724 553772
rect 95108 553732 95114 553744
rect 120718 553732 120724 553744
rect 120776 553732 120782 553784
rect 100754 553664 100760 553716
rect 100812 553704 100818 553716
rect 129090 553704 129096 553716
rect 100812 553676 129096 553704
rect 100812 553664 100818 553676
rect 129090 553664 129096 553676
rect 129148 553664 129154 553716
rect 106458 553596 106464 553648
rect 106516 553636 106522 553648
rect 140038 553636 140044 553648
rect 106516 553608 140044 553636
rect 106516 553596 106522 553608
rect 140038 553596 140044 553608
rect 140096 553596 140102 553648
rect 103698 553528 103704 553580
rect 103756 553568 103762 553580
rect 151078 553568 151084 553580
rect 103756 553540 151084 553568
rect 103756 553528 103762 553540
rect 151078 553528 151084 553540
rect 151136 553528 151142 553580
rect 97810 553460 97816 553512
rect 97868 553500 97874 553512
rect 157978 553500 157984 553512
rect 97868 553472 157984 553500
rect 97868 553460 97874 553472
rect 157978 553460 157984 553472
rect 158036 553460 158042 553512
rect 112346 553392 112352 553444
rect 112404 553432 112410 553444
rect 116026 553432 116032 553444
rect 112404 553404 116032 553432
rect 112404 553392 112410 553404
rect 116026 553392 116032 553404
rect 116084 553392 116090 553444
rect 3142 552032 3148 552084
rect 3200 552072 3206 552084
rect 28258 552072 28264 552084
rect 3200 552044 28264 552072
rect 3200 552032 3206 552044
rect 28258 552032 28264 552044
rect 28316 552032 28322 552084
rect 153289 550647 153347 550653
rect 153289 550613 153301 550647
rect 153335 550644 153347 550647
rect 153470 550644 153476 550656
rect 153335 550616 153476 550644
rect 153335 550613 153347 550616
rect 153289 550607 153347 550613
rect 153470 550604 153476 550616
rect 153528 550604 153534 550656
rect 85482 549856 85488 549908
rect 85540 549896 85546 549908
rect 86402 549896 86408 549908
rect 85540 549868 86408 549896
rect 85540 549856 85546 549868
rect 86402 549856 86408 549868
rect 86460 549896 86466 549908
rect 115382 549896 115388 549908
rect 86460 549868 115388 549896
rect 86460 549856 86466 549868
rect 115382 549856 115388 549868
rect 115440 549856 115446 549908
rect 153286 543600 153292 543652
rect 153344 543640 153350 543652
rect 153470 543640 153476 543652
rect 153344 543612 153476 543640
rect 153344 543600 153350 543612
rect 153470 543600 153476 543612
rect 153528 543600 153534 543652
rect 286870 538228 286876 538280
rect 286928 538268 286934 538280
rect 297726 538268 297732 538280
rect 286928 538240 297732 538268
rect 286928 538228 286934 538240
rect 297726 538228 297732 538240
rect 297784 538228 297790 538280
rect 117314 536800 117320 536852
rect 117372 536840 117378 536852
rect 146938 536840 146944 536852
rect 117372 536812 146944 536840
rect 117372 536800 117378 536812
rect 146938 536800 146944 536812
rect 146996 536800 147002 536852
rect 118234 534012 118240 534064
rect 118292 534052 118298 534064
rect 118510 534052 118516 534064
rect 118292 534024 118516 534052
rect 118292 534012 118298 534024
rect 118510 534012 118516 534024
rect 118568 534012 118574 534064
rect 153286 534012 153292 534064
rect 153344 534052 153350 534064
rect 153470 534052 153476 534064
rect 153344 534024 153476 534052
rect 153344 534012 153350 534024
rect 153470 534012 153476 534024
rect 153528 534012 153534 534064
rect 295978 532856 295984 532908
rect 296036 532896 296042 532908
rect 297450 532896 297456 532908
rect 296036 532868 297456 532896
rect 296036 532856 296042 532868
rect 297450 532856 297456 532868
rect 297508 532856 297514 532908
rect 117314 532720 117320 532772
rect 117372 532760 117378 532772
rect 160738 532760 160744 532772
rect 117372 532732 160744 532760
rect 117372 532720 117378 532732
rect 160738 532720 160744 532732
rect 160796 532720 160802 532772
rect 514018 532720 514024 532772
rect 514076 532760 514082 532772
rect 580166 532760 580172 532772
rect 514076 532732 580172 532760
rect 514076 532720 514082 532732
rect 580166 532720 580172 532732
rect 580224 532720 580230 532772
rect 117958 529864 117964 529916
rect 118016 529904 118022 529916
rect 119338 529904 119344 529916
rect 118016 529876 119344 529904
rect 118016 529864 118022 529876
rect 119338 529864 119344 529876
rect 119396 529864 119402 529916
rect 117314 525036 117320 525088
rect 117372 525076 117378 525088
rect 129182 525076 129188 525088
rect 117372 525048 129188 525076
rect 117372 525036 117378 525048
rect 129182 525036 129188 525048
rect 129240 525036 129246 525088
rect 118510 524532 118516 524544
rect 118436 524504 118516 524532
rect 70302 524424 70308 524476
rect 70360 524464 70366 524476
rect 82814 524464 82820 524476
rect 70360 524436 82820 524464
rect 70360 524424 70366 524436
rect 82814 524424 82820 524436
rect 82872 524424 82878 524476
rect 118436 524408 118464 524504
rect 118510 524492 118516 524504
rect 118568 524492 118574 524544
rect 118418 524356 118424 524408
rect 118476 524356 118482 524408
rect 128906 521636 128912 521688
rect 128964 521676 128970 521688
rect 129182 521676 129188 521688
rect 128964 521648 129188 521676
rect 128964 521636 128970 521648
rect 129182 521636 129188 521648
rect 129240 521636 129246 521688
rect 153562 521636 153568 521688
rect 153620 521676 153626 521688
rect 153746 521676 153752 521688
rect 153620 521648 153752 521676
rect 153620 521636 153626 521648
rect 153746 521636 153752 521648
rect 153804 521636 153810 521688
rect 280062 521636 280068 521688
rect 280120 521676 280126 521688
rect 297082 521676 297088 521688
rect 280120 521648 297088 521676
rect 280120 521636 280126 521648
rect 297082 521636 297088 521648
rect 297140 521636 297146 521688
rect 295334 521568 295340 521620
rect 295392 521608 295398 521620
rect 295978 521608 295984 521620
rect 295392 521580 295984 521608
rect 295392 521568 295398 521580
rect 295978 521568 295984 521580
rect 296036 521568 296042 521620
rect 85298 521228 85304 521280
rect 85356 521268 85362 521280
rect 295334 521268 295340 521280
rect 85356 521240 295340 521268
rect 85356 521228 85362 521240
rect 295334 521228 295340 521240
rect 295392 521228 295398 521280
rect 199378 521092 199384 521144
rect 199436 521132 199442 521144
rect 222378 521132 222384 521144
rect 199436 521104 222384 521132
rect 199436 521092 199442 521104
rect 222378 521092 222384 521104
rect 222436 521092 222442 521144
rect 199470 521024 199476 521076
rect 199528 521064 199534 521076
rect 222562 521064 222568 521076
rect 199528 521036 222568 521064
rect 199528 521024 199534 521036
rect 222562 521024 222568 521036
rect 222620 521024 222626 521076
rect 198274 520956 198280 521008
rect 198332 520996 198338 521008
rect 222654 520996 222660 521008
rect 198332 520968 222660 520996
rect 198332 520956 198338 520968
rect 222654 520956 222660 520968
rect 222712 520956 222718 521008
rect 117314 520888 117320 520940
rect 117372 520928 117378 520940
rect 128446 520928 128452 520940
rect 117372 520900 128452 520928
rect 117372 520888 117378 520900
rect 128446 520888 128452 520900
rect 128504 520928 128510 520940
rect 128998 520928 129004 520940
rect 128504 520900 129004 520928
rect 128504 520888 128510 520900
rect 128998 520888 129004 520900
rect 129056 520888 129062 520940
rect 198182 520888 198188 520940
rect 198240 520928 198246 520940
rect 222470 520928 222476 520940
rect 198240 520900 222476 520928
rect 198240 520888 198246 520900
rect 222470 520888 222476 520900
rect 222528 520888 222534 520940
rect 96525 518959 96583 518965
rect 96525 518956 96537 518959
rect 87984 518928 96537 518956
rect 86586 518712 86592 518764
rect 86644 518752 86650 518764
rect 87984 518752 88012 518928
rect 96525 518925 96537 518928
rect 96571 518925 96583 518959
rect 96525 518919 96583 518925
rect 115937 518959 115995 518965
rect 115937 518925 115949 518959
rect 115983 518956 115995 518959
rect 122742 518956 122748 518968
rect 115983 518928 122748 518956
rect 115983 518925 115995 518928
rect 115937 518919 115995 518925
rect 122742 518916 122748 518928
rect 122800 518956 122806 518968
rect 125505 518959 125563 518965
rect 125505 518956 125517 518959
rect 122800 518928 125517 518956
rect 122800 518916 122806 518928
rect 125505 518925 125517 518928
rect 125551 518925 125563 518959
rect 125505 518919 125563 518925
rect 279418 518916 279424 518968
rect 279476 518956 279482 518968
rect 297726 518956 297732 518968
rect 279476 518928 297732 518956
rect 279476 518916 279482 518928
rect 297726 518916 297732 518928
rect 297784 518916 297790 518968
rect 89346 518848 89352 518900
rect 89404 518888 89410 518900
rect 129826 518888 129832 518900
rect 89404 518860 129832 518888
rect 89404 518848 89410 518860
rect 129826 518848 129832 518860
rect 129884 518888 129890 518900
rect 130378 518888 130384 518900
rect 129884 518860 130384 518888
rect 129884 518848 129890 518860
rect 130378 518848 130384 518860
rect 130436 518848 130442 518900
rect 109586 518780 109592 518832
rect 109644 518820 109650 518832
rect 113818 518820 113824 518832
rect 109644 518792 113824 518820
rect 109644 518780 109650 518792
rect 113818 518780 113824 518792
rect 113876 518820 113882 518832
rect 115198 518820 115204 518832
rect 113876 518792 115204 518820
rect 113876 518780 113882 518792
rect 115198 518780 115204 518792
rect 115256 518780 115262 518832
rect 125505 518823 125563 518829
rect 125505 518789 125517 518823
rect 125551 518820 125563 518823
rect 127710 518820 127716 518832
rect 125551 518792 127716 518820
rect 125551 518789 125563 518792
rect 125505 518783 125563 518789
rect 127710 518780 127716 518792
rect 127768 518780 127774 518832
rect 86644 518724 88012 518752
rect 96525 518755 96583 518761
rect 86644 518712 86650 518724
rect 96525 518721 96537 518755
rect 96571 518752 96583 518755
rect 96571 518724 99328 518752
rect 96571 518721 96583 518724
rect 96525 518715 96583 518721
rect 99300 518684 99328 518724
rect 115937 518687 115995 518693
rect 115937 518684 115949 518687
rect 99300 518656 115949 518684
rect 115937 518653 115949 518656
rect 115983 518653 115995 518687
rect 115937 518647 115995 518653
rect 97994 518372 98000 518424
rect 98052 518412 98058 518424
rect 144178 518412 144184 518424
rect 98052 518384 144184 518412
rect 98052 518372 98058 518384
rect 144178 518372 144184 518384
rect 144236 518372 144242 518424
rect 106642 518304 106648 518356
rect 106700 518344 106706 518356
rect 153838 518344 153844 518356
rect 106700 518316 153844 518344
rect 106700 518304 106706 518316
rect 153838 518304 153844 518316
rect 153896 518304 153902 518356
rect 100938 518236 100944 518288
rect 100996 518276 101002 518288
rect 159358 518276 159364 518288
rect 100996 518248 159364 518276
rect 100996 518236 101002 518248
rect 159358 518236 159364 518248
rect 159416 518236 159422 518288
rect 198090 518236 198096 518288
rect 198148 518276 198154 518288
rect 218974 518276 218980 518288
rect 198148 518248 218980 518276
rect 198148 518236 198154 518248
rect 218974 518236 218980 518248
rect 219032 518236 219038 518288
rect 92290 518168 92296 518220
rect 92348 518208 92354 518220
rect 126974 518208 126980 518220
rect 92348 518180 126980 518208
rect 92348 518168 92354 518180
rect 126974 518168 126980 518180
rect 127032 518208 127038 518220
rect 297450 518208 297456 518220
rect 127032 518180 297456 518208
rect 127032 518168 127038 518180
rect 297450 518168 297456 518180
rect 297508 518168 297514 518220
rect 205634 517488 205640 517540
rect 205692 517528 205698 517540
rect 206646 517528 206652 517540
rect 205692 517500 206652 517528
rect 205692 517488 205698 517500
rect 206646 517488 206652 517500
rect 206704 517488 206710 517540
rect 284938 516128 284944 516180
rect 284996 516168 285002 516180
rect 297726 516168 297732 516180
rect 284996 516140 297732 516168
rect 284996 516128 285002 516140
rect 297726 516128 297732 516140
rect 297784 516128 297790 516180
rect 118234 511980 118240 512032
rect 118292 512020 118298 512032
rect 118510 512020 118516 512032
rect 118292 511992 118516 512020
rect 118292 511980 118298 511992
rect 118510 511980 118516 511992
rect 118568 511980 118574 512032
rect 293862 509260 293868 509312
rect 293920 509300 293926 509312
rect 297634 509300 297640 509312
rect 293920 509272 297640 509300
rect 293920 509260 293926 509272
rect 297634 509260 297640 509272
rect 297692 509260 297698 509312
rect 192478 506472 192484 506524
rect 192536 506512 192542 506524
rect 297634 506512 297640 506524
rect 192536 506484 297640 506512
rect 192536 506472 192542 506484
rect 297634 506472 297640 506484
rect 297692 506472 297698 506524
rect 153378 505152 153384 505164
rect 153339 505124 153384 505152
rect 153378 505112 153384 505124
rect 153436 505112 153442 505164
rect 380710 503112 380716 503124
rect 380671 503084 380716 503112
rect 380710 503072 380716 503084
rect 380768 503072 380774 503124
rect 118326 502324 118332 502376
rect 118384 502364 118390 502376
rect 118510 502364 118516 502376
rect 118384 502336 118516 502364
rect 118384 502324 118390 502336
rect 118510 502324 118516 502336
rect 118568 502324 118574 502376
rect 128538 502324 128544 502376
rect 128596 502364 128602 502376
rect 128814 502364 128820 502376
rect 128596 502336 128820 502364
rect 128596 502324 128602 502336
rect 128814 502324 128820 502336
rect 128872 502324 128878 502376
rect 153378 502364 153384 502376
rect 153339 502336 153384 502364
rect 153378 502324 153384 502336
rect 153436 502324 153442 502376
rect 96522 500896 96528 500948
rect 96580 500936 96586 500948
rect 380434 500936 380440 500948
rect 96580 500908 380440 500936
rect 96580 500896 96586 500908
rect 380434 500896 380440 500908
rect 380492 500896 380498 500948
rect 380713 500939 380771 500945
rect 380713 500905 380725 500939
rect 380759 500905 380771 500939
rect 380713 500899 380771 500905
rect 103514 500828 103520 500880
rect 103572 500868 103578 500880
rect 104802 500868 104808 500880
rect 103572 500840 104808 500868
rect 103572 500828 103578 500840
rect 104802 500828 104808 500840
rect 104860 500868 104866 500880
rect 380728 500868 380756 500899
rect 104860 500840 380756 500868
rect 104860 500828 104866 500840
rect 380434 500760 380440 500812
rect 380492 500800 380498 500812
rect 380710 500800 380716 500812
rect 380492 500772 380716 500800
rect 380492 500760 380498 500772
rect 380710 500760 380716 500772
rect 380768 500760 380774 500812
rect 70210 500216 70216 500268
rect 70268 500256 70274 500268
rect 95234 500256 95240 500268
rect 70268 500228 95240 500256
rect 70268 500216 70274 500228
rect 95234 500216 95240 500228
rect 95292 500256 95298 500268
rect 96522 500256 96528 500268
rect 95292 500228 96528 500256
rect 95292 500216 95298 500228
rect 96522 500216 96528 500228
rect 96580 500216 96586 500268
rect 300486 499128 300492 499180
rect 300544 499168 300550 499180
rect 311894 499168 311900 499180
rect 300544 499140 311900 499168
rect 300544 499128 300550 499140
rect 311894 499128 311900 499140
rect 311952 499128 311958 499180
rect 298922 499060 298928 499112
rect 298980 499100 298986 499112
rect 310606 499100 310612 499112
rect 298980 499072 310612 499100
rect 298980 499060 298986 499072
rect 310606 499060 310612 499072
rect 310664 499060 310670 499112
rect 324222 499060 324228 499112
rect 324280 499100 324286 499112
rect 378410 499100 378416 499112
rect 324280 499072 378416 499100
rect 324280 499060 324286 499072
rect 378410 499060 378416 499072
rect 378468 499060 378474 499112
rect 299014 498992 299020 499044
rect 299072 499032 299078 499044
rect 314838 499032 314844 499044
rect 299072 499004 314844 499032
rect 299072 498992 299078 499004
rect 314838 498992 314844 499004
rect 314896 498992 314902 499044
rect 321462 498992 321468 499044
rect 321520 499032 321526 499044
rect 378502 499032 378508 499044
rect 321520 499004 378508 499032
rect 321520 498992 321526 499004
rect 378502 498992 378508 499004
rect 378560 498992 378566 499044
rect 298646 498924 298652 498976
rect 298704 498964 298710 498976
rect 316034 498964 316040 498976
rect 298704 498936 316040 498964
rect 298704 498924 298710 498936
rect 316034 498924 316040 498936
rect 316092 498924 316098 498976
rect 317322 498924 317328 498976
rect 317380 498964 317386 498976
rect 378870 498964 378876 498976
rect 317380 498936 378876 498964
rect 317380 498924 317386 498936
rect 378870 498924 378876 498936
rect 378928 498924 378934 498976
rect 298830 498856 298836 498908
rect 298888 498896 298894 498908
rect 309134 498896 309140 498908
rect 298888 498868 309140 498896
rect 298888 498856 298894 498868
rect 309134 498856 309140 498868
rect 309192 498856 309198 498908
rect 310422 498856 310428 498908
rect 310480 498896 310486 498908
rect 378686 498896 378692 498908
rect 310480 498868 378692 498896
rect 310480 498856 310486 498868
rect 378686 498856 378692 498868
rect 378744 498856 378750 498908
rect 298462 498788 298468 498840
rect 298520 498828 298526 498840
rect 306466 498828 306472 498840
rect 298520 498800 306472 498828
rect 298520 498788 298526 498800
rect 306466 498788 306472 498800
rect 306524 498788 306530 498840
rect 309042 498788 309048 498840
rect 309100 498828 309106 498840
rect 378594 498828 378600 498840
rect 309100 498800 378600 498828
rect 309100 498788 309106 498800
rect 378594 498788 378600 498800
rect 378652 498788 378658 498840
rect 298554 498244 298560 498296
rect 298612 498284 298618 498296
rect 302418 498284 302424 498296
rect 298612 498256 302424 498284
rect 298612 498244 298618 498256
rect 302418 498244 302424 498256
rect 302476 498244 302482 498296
rect 132126 498176 132132 498228
rect 132184 498216 132190 498228
rect 580166 498216 580172 498228
rect 132184 498188 580172 498216
rect 132184 498176 132190 498188
rect 580166 498176 580172 498188
rect 580224 498176 580230 498228
rect 129090 498108 129096 498160
rect 129148 498148 129154 498160
rect 364242 498148 364248 498160
rect 129148 498120 364248 498148
rect 129148 498108 129154 498120
rect 364242 498108 364248 498120
rect 364300 498108 364306 498160
rect 116026 498040 116032 498092
rect 116084 498080 116090 498092
rect 347314 498080 347320 498092
rect 116084 498052 347320 498080
rect 116084 498040 116090 498052
rect 347314 498040 347320 498052
rect 347372 498040 347378 498092
rect 120718 497972 120724 498024
rect 120776 498012 120782 498024
rect 121362 498012 121368 498024
rect 120776 497984 121368 498012
rect 120776 497972 120782 497984
rect 121362 497972 121368 497984
rect 121420 498012 121426 498024
rect 338850 498012 338856 498024
rect 121420 497984 338856 498012
rect 121420 497972 121426 497984
rect 338850 497972 338856 497984
rect 338908 497972 338914 498024
rect 111702 497904 111708 497956
rect 111760 497944 111766 497956
rect 115290 497944 115296 497956
rect 111760 497916 115296 497944
rect 111760 497904 111766 497916
rect 115290 497904 115296 497916
rect 115348 497944 115354 497956
rect 313274 497944 313280 497956
rect 115348 497916 313280 497944
rect 115348 497904 115354 497916
rect 313274 497904 313280 497916
rect 313332 497904 313338 497956
rect 320082 497904 320088 497956
rect 320140 497944 320146 497956
rect 357986 497944 357992 497956
rect 320140 497916 357992 497944
rect 320140 497904 320146 497916
rect 357986 497904 357992 497916
rect 358044 497904 358050 497956
rect 144178 497836 144184 497888
rect 144236 497876 144242 497888
rect 334434 497876 334440 497888
rect 144236 497848 334440 497876
rect 144236 497836 144242 497848
rect 334434 497836 334440 497848
rect 334492 497836 334498 497888
rect 338758 497836 338764 497888
rect 338816 497876 338822 497888
rect 362218 497876 362224 497888
rect 338816 497848 362224 497876
rect 338816 497836 338822 497848
rect 362218 497836 362224 497848
rect 362276 497836 362282 497888
rect 284110 497768 284116 497820
rect 284168 497808 284174 497820
rect 368474 497808 368480 497820
rect 284168 497780 368480 497808
rect 284168 497768 284174 497780
rect 368474 497768 368480 497780
rect 368532 497768 368538 497820
rect 291010 497700 291016 497752
rect 291068 497740 291074 497752
rect 377122 497740 377128 497752
rect 291068 497712 377128 497740
rect 291068 497700 291074 497712
rect 377122 497700 377128 497712
rect 377180 497700 377186 497752
rect 284202 497632 284208 497684
rect 284260 497672 284266 497684
rect 374914 497672 374920 497684
rect 284260 497644 374920 497672
rect 284260 497632 284266 497644
rect 374914 497632 374920 497644
rect 374972 497632 374978 497684
rect 108942 497564 108948 497616
rect 109000 497604 109006 497616
rect 116026 497604 116032 497616
rect 109000 497576 116032 497604
rect 109000 497564 109006 497576
rect 116026 497564 116032 497576
rect 116084 497564 116090 497616
rect 118050 497564 118056 497616
rect 118108 497604 118114 497616
rect 302602 497604 302608 497616
rect 118108 497576 302608 497604
rect 118108 497564 118114 497576
rect 302602 497564 302608 497576
rect 302660 497564 302666 497616
rect 304534 497564 304540 497616
rect 304592 497604 304598 497616
rect 366450 497604 366456 497616
rect 304592 497576 366456 497604
rect 304592 497564 304598 497576
rect 366450 497564 366456 497576
rect 366508 497564 366514 497616
rect 83918 497496 83924 497548
rect 83976 497536 83982 497548
rect 127066 497536 127072 497548
rect 83976 497508 127072 497536
rect 83976 497496 83982 497508
rect 127066 497496 127072 497508
rect 127124 497536 127130 497548
rect 360010 497536 360016 497548
rect 127124 497508 360016 497536
rect 127124 497496 127130 497508
rect 360010 497496 360016 497508
rect 360068 497496 360074 497548
rect 111794 497428 111800 497480
rect 111852 497468 111858 497480
rect 125870 497468 125876 497480
rect 111852 497440 125876 497468
rect 111852 497428 111858 497440
rect 125870 497428 125876 497440
rect 125928 497468 125934 497480
rect 372706 497468 372712 497480
rect 125928 497440 372712 497468
rect 125928 497428 125934 497440
rect 372706 497428 372712 497440
rect 372764 497428 372770 497480
rect 285582 497360 285588 497412
rect 285640 497400 285646 497412
rect 345106 497400 345112 497412
rect 285640 497372 345112 497400
rect 285640 497360 285646 497372
rect 345106 497360 345112 497372
rect 345164 497360 345170 497412
rect 292298 497292 292304 497344
rect 292356 497332 292362 497344
rect 351546 497332 351552 497344
rect 292356 497304 351552 497332
rect 292356 497292 292362 497304
rect 351546 497292 351552 497304
rect 351604 497292 351610 497344
rect 277302 497224 277308 497276
rect 277360 497264 277366 497276
rect 317506 497264 317512 497276
rect 277360 497236 317512 497264
rect 277360 497224 277366 497236
rect 317506 497224 317512 497236
rect 317564 497224 317570 497276
rect 337378 497224 337384 497276
rect 337436 497264 337442 497276
rect 355778 497264 355784 497276
rect 337436 497236 355784 497264
rect 337436 497224 337442 497236
rect 355778 497224 355784 497236
rect 355836 497224 355842 497276
rect 276658 497156 276664 497208
rect 276716 497196 276722 497208
rect 311066 497196 311072 497208
rect 276716 497168 311072 497196
rect 276716 497156 276722 497168
rect 311066 497156 311072 497168
rect 311124 497156 311130 497208
rect 315942 497156 315948 497208
rect 316000 497196 316006 497208
rect 349338 497196 349344 497208
rect 316000 497168 349344 497196
rect 316000 497156 316006 497168
rect 349338 497156 349344 497168
rect 349396 497156 349402 497208
rect 288345 497131 288403 497137
rect 288345 497097 288357 497131
rect 288391 497128 288403 497131
rect 321738 497128 321744 497140
rect 288391 497100 321744 497128
rect 288391 497097 288403 497100
rect 288345 497091 288403 497097
rect 321738 497088 321744 497100
rect 321796 497088 321802 497140
rect 301498 497020 301504 497072
rect 301556 497060 301562 497072
rect 325970 497060 325976 497072
rect 301556 497032 325976 497060
rect 301556 497020 301562 497032
rect 325970 497020 325976 497032
rect 326028 497020 326034 497072
rect 286410 496952 286416 497004
rect 286468 496992 286474 497004
rect 306834 496992 306840 497004
rect 286468 496964 306840 496992
rect 286468 496952 286474 496964
rect 306834 496952 306840 496964
rect 306892 496952 306898 497004
rect 308950 496952 308956 497004
rect 309008 496992 309014 497004
rect 321738 496992 321744 497004
rect 309008 496964 321744 496992
rect 309008 496952 309014 496964
rect 321738 496952 321744 496964
rect 321796 496952 321802 497004
rect 305638 496884 305644 496936
rect 305696 496924 305702 496936
rect 323946 496924 323952 496936
rect 305696 496896 323952 496924
rect 305696 496884 305702 496896
rect 323946 496884 323952 496896
rect 324004 496884 324010 496936
rect 302142 496816 302148 496868
rect 302200 496856 302206 496868
rect 302602 496856 302608 496868
rect 302200 496828 302608 496856
rect 302200 496816 302206 496828
rect 302602 496816 302608 496828
rect 302660 496816 302666 496868
rect 308398 496816 308404 496868
rect 308456 496856 308462 496868
rect 315298 496856 315304 496868
rect 308456 496828 315304 496856
rect 308456 496816 308462 496828
rect 315298 496816 315304 496828
rect 315356 496816 315362 496868
rect 330478 496816 330484 496868
rect 330536 496856 330542 496868
rect 336642 496856 336648 496868
rect 330536 496828 336648 496856
rect 330536 496816 330542 496828
rect 336642 496816 336648 496828
rect 336700 496816 336706 496868
rect 340138 496816 340144 496868
rect 340196 496856 340202 496868
rect 343082 496856 343088 496868
rect 340196 496828 343088 496856
rect 340196 496816 340202 496828
rect 343082 496816 343088 496828
rect 343140 496816 343146 496868
rect 3326 495456 3332 495508
rect 3384 495496 3390 495508
rect 31018 495496 31024 495508
rect 3384 495468 31024 495496
rect 3384 495456 3390 495468
rect 31018 495456 31024 495468
rect 31076 495456 31082 495508
rect 153378 495388 153384 495440
rect 153436 495428 153442 495440
rect 153562 495428 153568 495440
rect 153436 495400 153568 495428
rect 153436 495388 153442 495400
rect 153562 495388 153568 495400
rect 153620 495388 153626 495440
rect 288342 492708 288348 492720
rect 288303 492680 288348 492708
rect 288342 492668 288348 492680
rect 288400 492668 288406 492720
rect 118326 492600 118332 492652
rect 118384 492640 118390 492652
rect 118510 492640 118516 492652
rect 118384 492612 118516 492640
rect 118384 492600 118390 492612
rect 118510 492600 118516 492612
rect 118568 492600 118574 492652
rect 128538 492600 128544 492652
rect 128596 492640 128602 492652
rect 128722 492640 128728 492652
rect 128596 492612 128728 492640
rect 128596 492600 128602 492612
rect 128722 492600 128728 492612
rect 128780 492600 128786 492652
rect 153286 492600 153292 492652
rect 153344 492640 153350 492652
rect 153562 492640 153568 492652
rect 153344 492612 153568 492640
rect 153344 492600 153350 492612
rect 153562 492600 153568 492612
rect 153620 492600 153626 492652
rect 288342 485868 288348 485920
rect 288400 485868 288406 485920
rect 288250 485664 288256 485716
rect 288308 485704 288314 485716
rect 288360 485704 288388 485868
rect 299934 485800 299940 485852
rect 299992 485840 299998 485852
rect 300578 485840 300584 485852
rect 299992 485812 300584 485840
rect 299992 485800 299998 485812
rect 300578 485800 300584 485812
rect 300636 485800 300642 485852
rect 304166 485800 304172 485852
rect 304224 485800 304230 485852
rect 438210 485800 438216 485852
rect 438268 485840 438274 485852
rect 580166 485840 580172 485852
rect 438268 485812 580172 485840
rect 438268 485800 438274 485812
rect 580166 485800 580172 485812
rect 580224 485800 580230 485852
rect 288308 485676 288388 485704
rect 304184 485704 304212 485800
rect 304258 485704 304264 485716
rect 304184 485676 304264 485704
rect 288308 485664 288314 485676
rect 304258 485664 304264 485676
rect 304316 485664 304322 485716
rect 288250 482984 288256 482996
rect 288211 482956 288256 482984
rect 288250 482944 288256 482956
rect 288308 482944 288314 482996
rect 304258 482944 304264 482996
rect 304316 482984 304322 482996
rect 304442 482984 304448 482996
rect 304316 482956 304448 482984
rect 304316 482944 304322 482956
rect 304442 482944 304448 482956
rect 304500 482944 304506 482996
rect 4062 480632 4068 480684
rect 4120 480672 4126 480684
rect 4982 480672 4988 480684
rect 4120 480644 4988 480672
rect 4120 480632 4126 480644
rect 4982 480632 4988 480644
rect 5040 480632 5046 480684
rect 153286 476076 153292 476128
rect 153344 476116 153350 476128
rect 153470 476116 153476 476128
rect 153344 476088 153476 476116
rect 153344 476076 153350 476088
rect 153470 476076 153476 476088
rect 153528 476076 153534 476128
rect 299750 476076 299756 476128
rect 299808 476116 299814 476128
rect 299934 476116 299940 476128
rect 299808 476088 299940 476116
rect 299808 476076 299814 476088
rect 299934 476076 299940 476088
rect 299992 476076 299998 476128
rect 288250 476048 288256 476060
rect 288211 476020 288256 476048
rect 288250 476008 288256 476020
rect 288308 476008 288314 476060
rect 299842 473328 299848 473340
rect 299803 473300 299848 473328
rect 299842 473288 299848 473300
rect 299900 473288 299906 473340
rect 304258 473288 304264 473340
rect 304316 473328 304322 473340
rect 304350 473328 304356 473340
rect 304316 473300 304356 473328
rect 304316 473288 304322 473300
rect 304350 473288 304356 473300
rect 304408 473288 304414 473340
rect 118418 466528 118424 466540
rect 118344 466500 118424 466528
rect 118344 466404 118372 466500
rect 118418 466488 118424 466500
rect 118476 466488 118482 466540
rect 288253 466531 288311 466537
rect 288253 466497 288265 466531
rect 288299 466528 288311 466531
rect 288342 466528 288348 466540
rect 288299 466500 288348 466528
rect 288299 466497 288311 466500
rect 288253 466491 288311 466497
rect 288342 466488 288348 466500
rect 288400 466488 288406 466540
rect 153378 466420 153384 466472
rect 153436 466420 153442 466472
rect 118326 466352 118332 466404
rect 118384 466352 118390 466404
rect 153396 466392 153424 466420
rect 153470 466392 153476 466404
rect 153396 466364 153476 466392
rect 153470 466352 153476 466364
rect 153528 466352 153534 466404
rect 299842 466392 299848 466404
rect 299803 466364 299848 466392
rect 299842 466352 299848 466364
rect 299900 466352 299906 466404
rect 288250 463808 288256 463820
rect 288211 463780 288256 463808
rect 288250 463768 288256 463780
rect 288308 463768 288314 463820
rect 118050 463632 118056 463684
rect 118108 463672 118114 463684
rect 118326 463672 118332 463684
rect 118108 463644 118332 463672
rect 118108 463632 118114 463644
rect 118326 463632 118332 463644
rect 118384 463632 118390 463684
rect 153470 463672 153476 463684
rect 153431 463644 153476 463672
rect 153470 463632 153476 463644
rect 153528 463632 153534 463684
rect 288250 463672 288256 463684
rect 288211 463644 288256 463672
rect 288250 463632 288256 463644
rect 288308 463632 288314 463684
rect 133138 462340 133144 462392
rect 133196 462380 133202 462392
rect 579798 462380 579804 462392
rect 133196 462352 579804 462380
rect 133196 462340 133202 462352
rect 579798 462340 579804 462352
rect 579856 462340 579862 462392
rect 304258 456832 304264 456884
rect 304316 456832 304322 456884
rect 299750 456764 299756 456816
rect 299808 456804 299814 456816
rect 299934 456804 299940 456816
rect 299808 456776 299940 456804
rect 299808 456764 299814 456776
rect 299934 456764 299940 456776
rect 299992 456764 299998 456816
rect 304276 456748 304304 456832
rect 153470 456736 153476 456748
rect 153431 456708 153476 456736
rect 153470 456696 153476 456708
rect 153528 456696 153534 456748
rect 288250 456736 288256 456748
rect 288211 456708 288256 456736
rect 288250 456696 288256 456708
rect 288308 456696 288314 456748
rect 304258 456696 304264 456748
rect 304316 456696 304322 456748
rect 299842 454016 299848 454028
rect 299803 453988 299848 454016
rect 299842 453976 299848 453988
rect 299900 453976 299906 454028
rect 304258 453976 304264 454028
rect 304316 454016 304322 454028
rect 304350 454016 304356 454028
rect 304316 453988 304356 454016
rect 304316 453976 304322 453988
rect 304350 453976 304356 453988
rect 304408 453976 304414 454028
rect 304169 452591 304227 452597
rect 304169 452557 304181 452591
rect 304215 452588 304227 452591
rect 304350 452588 304356 452600
rect 304215 452560 304356 452588
rect 304215 452557 304227 452560
rect 304169 452551 304227 452557
rect 304350 452548 304356 452560
rect 304408 452548 304414 452600
rect 3050 451324 3056 451376
rect 3108 451364 3114 451376
rect 267274 451364 267280 451376
rect 3108 451336 267280 451364
rect 3108 451324 3114 451336
rect 267274 451324 267280 451336
rect 267332 451324 267338 451376
rect 133230 451256 133236 451308
rect 133288 451296 133294 451308
rect 580166 451296 580172 451308
rect 133288 451268 580172 451296
rect 133288 451256 133294 451268
rect 580166 451256 580172 451268
rect 580224 451256 580230 451308
rect 288342 447216 288348 447228
rect 288303 447188 288348 447216
rect 288342 447176 288348 447188
rect 288400 447176 288406 447228
rect 118234 447108 118240 447160
rect 118292 447108 118298 447160
rect 153378 447108 153384 447160
rect 153436 447148 153442 447160
rect 153562 447148 153568 447160
rect 153436 447120 153568 447148
rect 153436 447108 153442 447120
rect 153562 447108 153568 447120
rect 153620 447108 153626 447160
rect 118252 447080 118280 447108
rect 118326 447080 118332 447092
rect 118252 447052 118332 447080
rect 118326 447040 118332 447052
rect 118384 447040 118390 447092
rect 299842 447080 299848 447092
rect 299803 447052 299848 447080
rect 299842 447040 299848 447052
rect 299900 447040 299906 447092
rect 288342 444428 288348 444440
rect 288303 444400 288348 444428
rect 288342 444388 288348 444400
rect 288400 444388 288406 444440
rect 118050 444320 118056 444372
rect 118108 444360 118114 444372
rect 118326 444360 118332 444372
rect 118108 444332 118332 444360
rect 118108 444320 118114 444332
rect 118326 444320 118332 444332
rect 118384 444320 118390 444372
rect 153378 444360 153384 444372
rect 153339 444332 153384 444360
rect 153378 444320 153384 444332
rect 153436 444320 153442 444372
rect 288250 444360 288256 444372
rect 288211 444332 288256 444360
rect 288250 444320 288256 444332
rect 288308 444320 288314 444372
rect 436738 438880 436744 438932
rect 436796 438920 436802 438932
rect 580166 438920 580172 438932
rect 436796 438892 580172 438920
rect 436796 438880 436802 438892
rect 580166 438880 580172 438892
rect 580224 438880 580230 438932
rect 299750 437452 299756 437504
rect 299808 437492 299814 437504
rect 299934 437492 299940 437504
rect 299808 437464 299940 437492
rect 299808 437452 299814 437464
rect 299934 437452 299940 437464
rect 299992 437452 299998 437504
rect 153378 437424 153384 437436
rect 153339 437396 153384 437424
rect 153378 437384 153384 437396
rect 153436 437384 153442 437436
rect 288250 437424 288256 437436
rect 288211 437396 288256 437424
rect 288250 437384 288256 437396
rect 288308 437384 288314 437436
rect 304166 434772 304172 434784
rect 304127 434744 304172 434772
rect 304166 434732 304172 434744
rect 304224 434732 304230 434784
rect 299842 434704 299848 434716
rect 299803 434676 299848 434704
rect 299842 434664 299848 434676
rect 299900 434664 299906 434716
rect 288342 427904 288348 427916
rect 288303 427876 288348 427904
rect 288342 427864 288348 427876
rect 288400 427864 288406 427916
rect 118234 427796 118240 427848
rect 118292 427796 118298 427848
rect 118252 427768 118280 427796
rect 118326 427768 118332 427780
rect 118252 427740 118332 427768
rect 118326 427728 118332 427740
rect 118384 427728 118390 427780
rect 299842 427768 299848 427780
rect 299803 427740 299848 427768
rect 299842 427728 299848 427740
rect 299900 427728 299906 427780
rect 288342 425116 288348 425128
rect 288303 425088 288348 425116
rect 288342 425076 288348 425088
rect 288400 425076 288406 425128
rect 288066 425008 288072 425060
rect 288124 425048 288130 425060
rect 288250 425048 288256 425060
rect 288124 425020 288256 425048
rect 288124 425008 288130 425020
rect 288250 425008 288256 425020
rect 288308 425008 288314 425060
rect 4062 423648 4068 423700
rect 4120 423688 4126 423700
rect 5074 423688 5080 423700
rect 4120 423660 5080 423688
rect 4120 423648 4126 423660
rect 5074 423648 5080 423660
rect 5132 423648 5138 423700
rect 153286 418248 153292 418260
rect 153212 418220 153292 418248
rect 153212 418124 153240 418220
rect 153286 418208 153292 418220
rect 153344 418208 153350 418260
rect 304258 418248 304264 418260
rect 304184 418220 304264 418248
rect 299750 418140 299756 418192
rect 299808 418180 299814 418192
rect 299934 418180 299940 418192
rect 299808 418152 299940 418180
rect 299808 418140 299814 418152
rect 299934 418140 299940 418152
rect 299992 418140 299998 418192
rect 304184 418124 304212 418220
rect 304258 418208 304264 418220
rect 304316 418208 304322 418260
rect 153194 418072 153200 418124
rect 153252 418072 153258 418124
rect 304166 418072 304172 418124
rect 304224 418072 304230 418124
rect 132954 415420 132960 415472
rect 133012 415460 133018 415472
rect 579798 415460 579804 415472
rect 133012 415432 579804 415460
rect 133012 415420 133018 415432
rect 579798 415420 579804 415432
rect 579856 415420 579862 415472
rect 118418 415392 118424 415404
rect 118379 415364 118424 415392
rect 118418 415352 118424 415364
rect 118476 415352 118482 415404
rect 128541 415395 128599 415401
rect 128541 415361 128553 415395
rect 128587 415392 128599 415395
rect 128630 415392 128636 415404
rect 128587 415364 128636 415392
rect 128587 415361 128599 415364
rect 128541 415355 128599 415361
rect 128630 415352 128636 415364
rect 128688 415352 128694 415404
rect 299842 415392 299848 415404
rect 299803 415364 299848 415392
rect 299842 415352 299848 415364
rect 299900 415352 299906 415404
rect 248966 410796 248972 410848
rect 249024 410836 249030 410848
rect 266538 410836 266544 410848
rect 249024 410808 266544 410836
rect 249024 410796 249030 410808
rect 266538 410796 266544 410808
rect 266596 410796 266602 410848
rect 246022 410728 246028 410780
rect 246080 410768 246086 410780
rect 267734 410768 267740 410780
rect 246080 410740 267740 410768
rect 246080 410728 246086 410740
rect 267734 410728 267740 410740
rect 267792 410728 267798 410780
rect 234614 410660 234620 410712
rect 234672 410700 234678 410712
rect 266630 410700 266636 410712
rect 234672 410672 266636 410700
rect 234672 410660 234678 410672
rect 266630 410660 266636 410672
rect 266688 410660 266694 410712
rect 228910 410592 228916 410644
rect 228968 410632 228974 410644
rect 266998 410632 267004 410644
rect 228968 410604 267004 410632
rect 228968 410592 228974 410604
rect 266998 410592 267004 410604
rect 267056 410592 267062 410644
rect 223390 410524 223396 410576
rect 223448 410564 223454 410576
rect 266906 410564 266912 410576
rect 223448 410536 266912 410564
rect 223448 410524 223454 410536
rect 266906 410524 266912 410536
rect 266964 410524 266970 410576
rect 211982 410456 211988 410508
rect 212040 410496 212046 410508
rect 267090 410496 267096 410508
rect 212040 410468 267096 410496
rect 212040 410456 212046 410468
rect 267090 410456 267096 410468
rect 267148 410456 267154 410508
rect 206278 410388 206284 410440
rect 206336 410428 206342 410440
rect 266354 410428 266360 410440
rect 206336 410400 266360 410428
rect 206336 410388 206342 410400
rect 266354 410388 266360 410400
rect 266412 410388 266418 410440
rect 243262 410320 243268 410372
rect 243320 410360 243326 410372
rect 266814 410360 266820 410372
rect 243320 410332 266820 410360
rect 243320 410320 243326 410332
rect 266814 410320 266820 410332
rect 266872 410320 266878 410372
rect 240318 410252 240324 410304
rect 240376 410292 240382 410304
rect 266722 410292 266728 410304
rect 240376 410264 266728 410292
rect 240376 410252 240382 410264
rect 266722 410252 266728 410264
rect 266780 410252 266786 410304
rect 237558 410184 237564 410236
rect 237616 410224 237622 410236
rect 267642 410224 267648 410236
rect 237616 410196 267648 410224
rect 237616 410184 237622 410196
rect 267642 410184 267648 410196
rect 267700 410184 267706 410236
rect 196894 410116 196900 410168
rect 196952 410156 196958 410168
rect 200574 410156 200580 410168
rect 196952 410128 200580 410156
rect 196952 410116 196958 410128
rect 200574 410116 200580 410128
rect 200632 410116 200638 410168
rect 257430 410116 257436 410168
rect 257488 410156 257494 410168
rect 268746 410156 268752 410168
rect 257488 410128 268752 410156
rect 257488 410116 257494 410128
rect 268746 410116 268752 410128
rect 268804 410116 268810 410168
rect 199746 410048 199752 410100
rect 199804 410088 199810 410100
rect 217686 410088 217692 410100
rect 199804 410060 217692 410088
rect 199804 410048 199810 410060
rect 217686 410048 217692 410060
rect 217744 410048 217750 410100
rect 254670 410048 254676 410100
rect 254728 410088 254734 410100
rect 268838 410088 268844 410100
rect 254728 410060 268844 410088
rect 254728 410048 254734 410060
rect 268838 410048 268844 410060
rect 268896 410048 268902 410100
rect 199930 409980 199936 410032
rect 199988 410020 199994 410032
rect 220446 410020 220452 410032
rect 199988 409992 220452 410020
rect 199988 409980 199994 409992
rect 220446 409980 220452 409992
rect 220504 409980 220510 410032
rect 251726 409980 251732 410032
rect 251784 410020 251790 410032
rect 266446 410020 266452 410032
rect 251784 409992 266452 410020
rect 251784 409980 251790 409992
rect 266446 409980 266452 409992
rect 266504 409980 266510 410032
rect 200022 409912 200028 409964
rect 200080 409952 200086 409964
rect 214742 409952 214748 409964
rect 200080 409924 214748 409952
rect 200080 409912 200086 409924
rect 214742 409912 214748 409924
rect 214800 409912 214806 409964
rect 260374 409912 260380 409964
rect 260432 409952 260438 409964
rect 267550 409952 267556 409964
rect 260432 409924 267556 409952
rect 260432 409912 260438 409924
rect 267550 409912 267556 409924
rect 267608 409912 267614 409964
rect 199838 409844 199844 409896
rect 199896 409884 199902 409896
rect 209038 409884 209044 409896
rect 199896 409856 209044 409884
rect 199896 409844 199902 409856
rect 209038 409844 209044 409856
rect 209096 409844 209102 409896
rect 265894 409844 265900 409896
rect 265952 409884 265958 409896
rect 268930 409884 268936 409896
rect 265952 409856 268936 409884
rect 265952 409844 265958 409856
rect 268930 409844 268936 409856
rect 268988 409844 268994 409896
rect 199562 409640 199568 409692
rect 199620 409680 199626 409692
rect 202874 409680 202880 409692
rect 199620 409652 202880 409680
rect 199620 409640 199626 409652
rect 202874 409640 202880 409652
rect 202932 409640 202938 409692
rect 199654 409572 199660 409624
rect 199712 409612 199718 409624
rect 205634 409612 205640 409624
rect 199712 409584 205640 409612
rect 199712 409572 199718 409584
rect 205634 409572 205640 409584
rect 205692 409572 205698 409624
rect 196802 409504 196808 409556
rect 196860 409544 196866 409556
rect 209774 409544 209780 409556
rect 196860 409516 209780 409544
rect 196860 409504 196866 409516
rect 209774 409504 209780 409516
rect 209832 409504 209838 409556
rect 195698 409436 195704 409488
rect 195756 409476 195762 409488
rect 212534 409476 212540 409488
rect 195756 409448 212540 409476
rect 195756 409436 195762 409448
rect 212534 409436 212540 409448
rect 212592 409436 212598 409488
rect 195790 409368 195796 409420
rect 195848 409408 195854 409420
rect 215294 409408 215300 409420
rect 195848 409380 215300 409408
rect 195848 409368 195854 409380
rect 215294 409368 215300 409380
rect 215352 409368 215358 409420
rect 196710 409300 196716 409352
rect 196768 409340 196774 409352
rect 222746 409340 222752 409352
rect 196768 409312 222752 409340
rect 196768 409300 196774 409312
rect 222746 409300 222752 409312
rect 222804 409300 222810 409352
rect 196618 409232 196624 409284
rect 196676 409272 196682 409284
rect 222838 409272 222844 409284
rect 196676 409244 222844 409272
rect 196676 409232 196682 409244
rect 222838 409232 222844 409244
rect 222896 409232 222902 409284
rect 195606 409164 195612 409216
rect 195664 409204 195670 409216
rect 222194 409204 222200 409216
rect 195664 409176 222200 409204
rect 195664 409164 195670 409176
rect 222194 409164 222200 409176
rect 222252 409164 222258 409216
rect 195514 409096 195520 409148
rect 195572 409136 195578 409148
rect 222286 409136 222292 409148
rect 195572 409108 222292 409136
rect 195572 409096 195578 409108
rect 222286 409096 222292 409108
rect 222344 409096 222350 409148
rect 153194 408484 153200 408536
rect 153252 408484 153258 408536
rect 153212 408456 153240 408484
rect 153378 408456 153384 408468
rect 153212 408428 153384 408456
rect 153378 408416 153384 408428
rect 153436 408416 153442 408468
rect 287974 408348 287980 408400
rect 288032 408388 288038 408400
rect 288342 408388 288348 408400
rect 288032 408360 288348 408388
rect 288032 408348 288038 408360
rect 288342 408348 288348 408360
rect 288400 408348 288406 408400
rect 132865 407915 132923 407921
rect 132865 407881 132877 407915
rect 132911 407912 132923 407915
rect 380618 407912 380624 407924
rect 132911 407884 380624 407912
rect 132911 407881 132923 407884
rect 132865 407875 132923 407881
rect 380618 407872 380624 407884
rect 380676 407872 380682 407924
rect 70118 407804 70124 407856
rect 70176 407844 70182 407856
rect 104802 407844 104808 407856
rect 70176 407816 104808 407844
rect 70176 407804 70182 407816
rect 104802 407804 104808 407816
rect 104860 407844 104866 407856
rect 416958 407844 416964 407856
rect 104860 407816 416964 407844
rect 104860 407804 104866 407816
rect 416958 407804 416964 407816
rect 417016 407804 417022 407856
rect 71590 407736 71596 407788
rect 71648 407776 71654 407788
rect 85574 407776 85580 407788
rect 71648 407748 85580 407776
rect 71648 407736 71654 407748
rect 85574 407736 85580 407748
rect 85632 407776 85638 407788
rect 402974 407776 402980 407788
rect 85632 407748 402980 407776
rect 85632 407736 85638 407748
rect 402974 407736 402980 407748
rect 403032 407736 403038 407788
rect 197998 407192 198004 407244
rect 198056 407232 198062 407244
rect 411254 407232 411260 407244
rect 198056 407204 411260 407232
rect 198056 407192 198062 407204
rect 411254 407192 411260 407204
rect 411312 407192 411318 407244
rect 130378 407124 130384 407176
rect 130436 407164 130442 407176
rect 416866 407164 416872 407176
rect 130436 407136 416872 407164
rect 130436 407124 130442 407136
rect 416866 407124 416872 407136
rect 416924 407124 416930 407176
rect 222197 406895 222255 406901
rect 222197 406861 222209 406895
rect 222243 406892 222255 406895
rect 231765 406895 231823 406901
rect 231765 406892 231777 406895
rect 222243 406864 231777 406892
rect 222243 406861 222255 406864
rect 222197 406855 222255 406861
rect 231765 406861 231777 406864
rect 231811 406861 231823 406895
rect 231765 406855 231823 406861
rect 241517 406895 241575 406901
rect 241517 406861 241529 406895
rect 241563 406892 241575 406895
rect 251085 406895 251143 406901
rect 251085 406892 251097 406895
rect 241563 406864 251097 406892
rect 241563 406861 241575 406864
rect 241517 406855 241575 406861
rect 251085 406861 251097 406864
rect 251131 406861 251143 406895
rect 251085 406855 251143 406861
rect 202877 406759 202935 406765
rect 202877 406725 202889 406759
rect 202923 406756 202935 406759
rect 212445 406759 212503 406765
rect 212445 406756 212457 406759
rect 202923 406728 212457 406756
rect 202923 406725 202935 406728
rect 202877 406719 202935 406725
rect 212445 406725 212457 406728
rect 212491 406725 212503 406759
rect 212445 406719 212503 406725
rect 215389 406759 215447 406765
rect 215389 406725 215401 406759
rect 215435 406756 215447 406759
rect 222197 406759 222255 406765
rect 222197 406756 222209 406759
rect 215435 406728 222209 406756
rect 215435 406725 215447 406728
rect 215389 406719 215447 406725
rect 222197 406725 222209 406728
rect 222243 406725 222255 406759
rect 241517 406759 241575 406765
rect 241517 406756 241529 406759
rect 222197 406719 222255 406725
rect 236564 406728 241529 406756
rect 231765 406691 231823 406697
rect 231765 406657 231777 406691
rect 231811 406688 231823 406691
rect 234525 406691 234583 406697
rect 234525 406688 234537 406691
rect 231811 406660 234537 406688
rect 231811 406657 231823 406660
rect 231765 406651 231823 406657
rect 234525 406657 234537 406660
rect 234571 406657 234583 406691
rect 234525 406651 234583 406657
rect 234617 406691 234675 406697
rect 234617 406657 234629 406691
rect 234663 406688 234675 406691
rect 236564 406688 236592 406728
rect 241517 406725 241529 406728
rect 241563 406725 241575 406759
rect 260837 406759 260895 406765
rect 260837 406756 260849 406759
rect 241517 406719 241575 406725
rect 255884 406728 260849 406756
rect 234663 406660 236592 406688
rect 251085 406691 251143 406697
rect 234663 406657 234675 406660
rect 234617 406651 234675 406657
rect 251085 406657 251097 406691
rect 251131 406688 251143 406691
rect 253845 406691 253903 406697
rect 253845 406688 253857 406691
rect 251131 406660 253857 406688
rect 251131 406657 251143 406660
rect 251085 406651 251143 406657
rect 253845 406657 253857 406660
rect 253891 406657 253903 406691
rect 253845 406651 253903 406657
rect 253937 406691 253995 406697
rect 253937 406657 253949 406691
rect 253983 406688 253995 406691
rect 255884 406688 255912 406728
rect 260837 406725 260849 406728
rect 260883 406725 260895 406759
rect 260837 406719 260895 406725
rect 289817 406759 289875 406765
rect 289817 406725 289829 406759
rect 289863 406756 289875 406759
rect 295334 406756 295340 406768
rect 289863 406728 295340 406756
rect 289863 406725 289875 406728
rect 289817 406719 289875 406725
rect 295334 406716 295340 406728
rect 295392 406716 295398 406768
rect 253983 406660 255912 406688
rect 253983 406657 253995 406660
rect 253937 406651 253995 406657
rect 212445 406623 212503 406629
rect 212445 406589 212457 406623
rect 212491 406620 212503 406623
rect 215205 406623 215263 406629
rect 215205 406620 215217 406623
rect 212491 406592 215217 406620
rect 212491 406589 212503 406592
rect 212445 406583 212503 406589
rect 215205 406589 215217 406592
rect 215251 406589 215263 406623
rect 289817 406623 289875 406629
rect 289817 406620 289829 406623
rect 215205 406583 215263 406589
rect 282840 406592 289829 406620
rect 197722 406512 197728 406564
rect 197780 406552 197786 406564
rect 202877 406555 202935 406561
rect 202877 406552 202889 406555
rect 197780 406524 202889 406552
rect 197780 406512 197786 406524
rect 202877 406521 202889 406524
rect 202923 406521 202935 406555
rect 202877 406515 202935 406521
rect 260837 406555 260895 406561
rect 260837 406521 260849 406555
rect 260883 406552 260895 406555
rect 266081 406555 266139 406561
rect 266081 406552 266093 406555
rect 260883 406524 266093 406552
rect 260883 406521 260895 406524
rect 260837 406515 260895 406521
rect 266081 406521 266093 406524
rect 266127 406521 266139 406555
rect 266081 406515 266139 406521
rect 282840 406484 282868 406592
rect 289817 406589 289829 406592
rect 289863 406589 289875 406623
rect 289817 406583 289875 406589
rect 273272 406456 282868 406484
rect 266081 406419 266139 406425
rect 266081 406385 266093 406419
rect 266127 406416 266139 406419
rect 273272 406416 273300 406456
rect 266127 406388 273300 406416
rect 266127 406385 266139 406388
rect 266081 406379 266139 406385
rect 295334 405832 295340 405884
rect 295392 405872 295398 405884
rect 295978 405872 295984 405884
rect 295392 405844 295984 405872
rect 295392 405832 295398 405844
rect 295978 405832 295984 405844
rect 296036 405832 296042 405884
rect 118421 405739 118479 405745
rect 118421 405705 118433 405739
rect 118467 405736 118479 405739
rect 118510 405736 118516 405748
rect 118467 405708 118516 405736
rect 118467 405705 118479 405708
rect 118421 405699 118479 405705
rect 118510 405696 118516 405708
rect 118568 405696 118574 405748
rect 128538 405736 128544 405748
rect 128499 405708 128544 405736
rect 128538 405696 128544 405708
rect 128596 405696 128602 405748
rect 132862 405736 132868 405748
rect 132823 405708 132868 405736
rect 132862 405696 132868 405708
rect 132920 405696 132926 405748
rect 299845 405739 299903 405745
rect 299845 405705 299857 405739
rect 299891 405736 299903 405739
rect 299934 405736 299940 405748
rect 299891 405708 299940 405736
rect 299891 405705 299903 405708
rect 299845 405699 299903 405705
rect 299934 405696 299940 405708
rect 299992 405696 299998 405748
rect 128538 404308 128544 404320
rect 128499 404280 128544 404308
rect 128538 404268 128544 404280
rect 128596 404268 128602 404320
rect 153378 398936 153384 398948
rect 153339 398908 153384 398936
rect 153378 398896 153384 398908
rect 153436 398896 153442 398948
rect 304258 398896 304264 398948
rect 304316 398896 304322 398948
rect 71682 398828 71688 398880
rect 71740 398868 71746 398880
rect 85482 398868 85488 398880
rect 71740 398840 85488 398868
rect 71740 398828 71746 398840
rect 85482 398828 85488 398840
rect 85540 398828 85546 398880
rect 120902 398828 120908 398880
rect 120960 398868 120966 398880
rect 121362 398868 121368 398880
rect 120960 398840 121368 398868
rect 120960 398828 120966 398840
rect 121362 398828 121368 398840
rect 121420 398868 121426 398880
rect 125686 398868 125692 398880
rect 121420 398840 125692 398868
rect 121420 398828 121426 398840
rect 125686 398828 125692 398840
rect 125744 398828 125750 398880
rect 304276 398812 304304 398896
rect 117314 398760 117320 398812
rect 117372 398800 117378 398812
rect 118602 398800 118608 398812
rect 117372 398772 118608 398800
rect 117372 398760 117378 398772
rect 118602 398760 118608 398772
rect 118660 398800 118666 398812
rect 129734 398800 129740 398812
rect 118660 398772 129740 398800
rect 118660 398760 118666 398772
rect 129734 398760 129740 398772
rect 129792 398760 129798 398812
rect 132678 398760 132684 398812
rect 132736 398800 132742 398812
rect 132862 398800 132868 398812
rect 132736 398772 132868 398800
rect 132736 398760 132742 398772
rect 132862 398760 132868 398772
rect 132920 398760 132926 398812
rect 304258 398760 304264 398812
rect 304316 398760 304322 398812
rect 85482 398692 85488 398744
rect 85540 398732 85546 398744
rect 90266 398732 90272 398744
rect 85540 398704 90272 398732
rect 85540 398692 85546 398704
rect 90266 398692 90272 398704
rect 90324 398692 90330 398744
rect 129734 398284 129740 398336
rect 129792 398324 129798 398336
rect 130378 398324 130384 398336
rect 129792 398296 130384 398324
rect 129792 398284 129798 398296
rect 130378 398284 130384 398296
rect 130436 398284 130442 398336
rect 100662 398216 100668 398268
rect 100720 398256 100726 398268
rect 113818 398256 113824 398268
rect 100720 398228 113824 398256
rect 100720 398216 100726 398228
rect 113818 398216 113824 398228
rect 113876 398256 113882 398268
rect 129458 398256 129464 398268
rect 113876 398228 129464 398256
rect 113876 398216 113882 398228
rect 129458 398216 129464 398228
rect 129516 398216 129522 398268
rect 85942 398148 85948 398200
rect 86000 398188 86006 398200
rect 117314 398188 117320 398200
rect 86000 398160 117320 398188
rect 86000 398148 86006 398160
rect 117314 398148 117320 398160
rect 117372 398148 117378 398200
rect 75822 398080 75828 398132
rect 75880 398120 75886 398132
rect 115934 398120 115940 398132
rect 75880 398092 115940 398120
rect 75880 398080 75886 398092
rect 115934 398080 115940 398092
rect 115992 398120 115998 398132
rect 127158 398120 127164 398132
rect 115992 398092 127164 398120
rect 115992 398080 115998 398092
rect 127158 398080 127164 398092
rect 127216 398080 127222 398132
rect 133046 398080 133052 398132
rect 133104 398120 133110 398132
rect 175918 398120 175924 398132
rect 133104 398092 175924 398120
rect 133104 398080 133110 398092
rect 175918 398080 175924 398092
rect 175976 398080 175982 398132
rect 80790 397808 80796 397860
rect 80848 397848 80854 397860
rect 126146 397848 126152 397860
rect 80848 397820 126152 397848
rect 80848 397808 80854 397820
rect 126146 397808 126152 397820
rect 126204 397848 126210 397860
rect 126330 397848 126336 397860
rect 126204 397820 126336 397848
rect 126204 397808 126210 397820
rect 126330 397808 126336 397820
rect 126388 397808 126394 397860
rect 115842 397740 115848 397792
rect 115900 397780 115906 397792
rect 126422 397780 126428 397792
rect 115900 397752 126428 397780
rect 115900 397740 115906 397752
rect 126422 397740 126428 397752
rect 126480 397740 126486 397792
rect 110966 397672 110972 397724
rect 111024 397712 111030 397724
rect 111702 397712 111708 397724
rect 111024 397684 111708 397712
rect 111024 397672 111030 397684
rect 111702 397672 111708 397684
rect 111760 397712 111766 397724
rect 127250 397712 127256 397724
rect 111760 397684 127256 397712
rect 111760 397672 111766 397684
rect 127250 397672 127256 397684
rect 127308 397672 127314 397724
rect 105998 397604 106004 397656
rect 106056 397644 106062 397656
rect 127618 397644 127624 397656
rect 106056 397616 127624 397644
rect 106056 397604 106062 397616
rect 127618 397604 127624 397616
rect 127676 397604 127682 397656
rect 95878 397536 95884 397588
rect 95936 397576 95942 397588
rect 133046 397576 133052 397588
rect 95936 397548 133052 397576
rect 95936 397536 95942 397548
rect 133046 397536 133052 397548
rect 133104 397536 133110 397588
rect 125594 397468 125600 397520
rect 125652 397508 125658 397520
rect 144178 397508 144184 397520
rect 125652 397480 144184 397508
rect 125652 397468 125658 397480
rect 144178 397468 144184 397480
rect 144236 397468 144242 397520
rect 129458 397400 129464 397452
rect 129516 397440 129522 397452
rect 197998 397440 198004 397452
rect 129516 397412 198004 397440
rect 129516 397400 129522 397412
rect 197998 397400 198004 397412
rect 198056 397400 198062 397452
rect 69934 396720 69940 396772
rect 69992 396760 69998 396772
rect 117958 396760 117964 396772
rect 69992 396732 117964 396760
rect 69992 396720 69998 396732
rect 117958 396720 117964 396732
rect 118016 396760 118022 396772
rect 126514 396760 126520 396772
rect 118016 396732 126520 396760
rect 118016 396720 118022 396732
rect 126514 396720 126520 396732
rect 126572 396720 126578 396772
rect 153378 396080 153384 396092
rect 153339 396052 153384 396080
rect 153378 396040 153384 396052
rect 153436 396040 153442 396092
rect 299842 396040 299848 396092
rect 299900 396080 299906 396092
rect 299934 396080 299940 396092
rect 299900 396052 299940 396080
rect 299900 396040 299906 396052
rect 299934 396040 299940 396052
rect 299992 396040 299998 396092
rect 153289 395947 153347 395953
rect 153289 395913 153301 395947
rect 153335 395944 153347 395947
rect 153378 395944 153384 395956
rect 153335 395916 153384 395944
rect 153335 395913 153347 395916
rect 153289 395907 153347 395913
rect 153378 395904 153384 395916
rect 153436 395904 153442 395956
rect 84010 395836 84016 395888
rect 84068 395876 84074 395888
rect 84105 395879 84163 395885
rect 84105 395876 84117 395879
rect 84068 395848 84117 395876
rect 84068 395836 84074 395848
rect 84105 395845 84117 395848
rect 84151 395845 84163 395879
rect 84105 395839 84163 395845
rect 84013 395743 84071 395749
rect 84013 395709 84025 395743
rect 84059 395740 84071 395743
rect 84102 395740 84108 395752
rect 84059 395712 84108 395740
rect 84059 395709 84071 395712
rect 84013 395703 84071 395709
rect 84102 395700 84108 395712
rect 84160 395700 84166 395752
rect 70026 395632 70032 395684
rect 70084 395672 70090 395684
rect 108942 395672 108948 395684
rect 70084 395644 108948 395672
rect 70084 395632 70090 395644
rect 108942 395632 108948 395644
rect 109000 395672 109006 395684
rect 125778 395672 125784 395684
rect 109000 395644 125784 395672
rect 109000 395632 109006 395644
rect 125778 395632 125784 395644
rect 125836 395632 125842 395684
rect 84013 395607 84071 395613
rect 84013 395573 84025 395607
rect 84059 395573 84071 395607
rect 84013 395567 84071 395573
rect 84105 395607 84163 395613
rect 84105 395573 84117 395607
rect 84151 395604 84163 395607
rect 168650 395604 168656 395616
rect 84151 395576 168656 395604
rect 84151 395573 84163 395576
rect 84105 395567 84163 395573
rect 84028 395536 84056 395567
rect 168650 395564 168656 395576
rect 168708 395564 168714 395616
rect 179506 395536 179512 395548
rect 84028 395508 179512 395536
rect 179506 395496 179512 395508
rect 179564 395496 179570 395548
rect 128541 394723 128599 394729
rect 128541 394689 128553 394723
rect 128587 394720 128599 394723
rect 128630 394720 128636 394732
rect 128587 394692 128636 394720
rect 128587 394689 128599 394692
rect 128541 394683 128599 394689
rect 128630 394680 128636 394692
rect 128688 394680 128694 394732
rect 402974 393252 402980 393304
rect 403032 393292 403038 393304
rect 403894 393292 403900 393304
rect 403032 393264 403900 393292
rect 403032 393252 403038 393264
rect 403894 393252 403900 393264
rect 403952 393252 403958 393304
rect 288158 391892 288164 391944
rect 288216 391932 288222 391944
rect 288342 391932 288348 391944
rect 288216 391904 288348 391932
rect 288216 391892 288222 391904
rect 288342 391892 288348 391904
rect 288400 391892 288406 391944
rect 69658 390532 69664 390584
rect 69716 390572 69722 390584
rect 71590 390572 71596 390584
rect 69716 390544 71596 390572
rect 69716 390532 69722 390544
rect 71590 390532 71596 390544
rect 71648 390532 71654 390584
rect 416590 389376 416596 389428
rect 416648 389416 416654 389428
rect 464246 389416 464252 389428
rect 416648 389388 464252 389416
rect 416648 389376 416654 389388
rect 464246 389376 464252 389388
rect 464304 389376 464310 389428
rect 414658 389308 414664 389360
rect 414716 389348 414722 389360
rect 475838 389348 475844 389360
rect 414716 389320 475844 389348
rect 414716 389308 414722 389320
rect 475838 389308 475844 389320
rect 475896 389308 475902 389360
rect 132862 389240 132868 389292
rect 132920 389240 132926 389292
rect 418062 389240 418068 389292
rect 418120 389280 418126 389292
rect 487430 389280 487436 389292
rect 418120 389252 487436 389280
rect 418120 389240 418126 389252
rect 487430 389240 487436 389252
rect 487488 389240 487494 389292
rect 132880 389156 132908 389240
rect 304258 389172 304264 389224
rect 304316 389172 304322 389224
rect 416682 389172 416688 389224
rect 416740 389212 416746 389224
rect 499022 389212 499028 389224
rect 416740 389184 499028 389212
rect 416740 389172 416746 389184
rect 499022 389172 499028 389184
rect 499080 389172 499086 389224
rect 132862 389104 132868 389156
rect 132920 389104 132926 389156
rect 153286 389144 153292 389156
rect 153247 389116 153292 389144
rect 153286 389104 153292 389116
rect 153344 389104 153350 389156
rect 304166 389104 304172 389156
rect 304224 389144 304230 389156
rect 304276 389144 304304 389172
rect 304224 389116 304304 389144
rect 304224 389104 304230 389116
rect 128722 388424 128728 388476
rect 128780 388464 128786 388476
rect 128817 388467 128875 388473
rect 128817 388464 128829 388467
rect 128780 388436 128829 388464
rect 128780 388424 128786 388436
rect 128817 388433 128829 388436
rect 128863 388433 128875 388467
rect 128817 388427 128875 388433
rect 375282 387064 375288 387116
rect 375340 387104 375346 387116
rect 478874 387104 478880 387116
rect 375340 387076 478880 387104
rect 375340 387064 375346 387076
rect 478874 387064 478880 387076
rect 478932 387064 478938 387116
rect 304258 386356 304264 386368
rect 304219 386328 304264 386356
rect 304258 386316 304264 386328
rect 304316 386316 304322 386368
rect 344922 385772 344928 385824
rect 344980 385812 344986 385824
rect 408862 385812 408868 385824
rect 344980 385784 408868 385812
rect 344980 385772 344986 385784
rect 408862 385772 408868 385784
rect 408920 385772 408926 385824
rect 295978 385704 295984 385756
rect 296036 385744 296042 385756
rect 388254 385744 388260 385756
rect 296036 385716 388260 385744
rect 296036 385704 296042 385716
rect 388254 385704 388260 385716
rect 388312 385704 388318 385756
rect 267274 385636 267280 385688
rect 267332 385676 267338 385688
rect 436094 385676 436100 385688
rect 267332 385648 436100 385676
rect 267332 385636 267338 385648
rect 436094 385636 436100 385648
rect 436152 385636 436158 385688
rect 369118 385568 369124 385620
rect 369176 385608 369182 385620
rect 392854 385608 392860 385620
rect 369176 385580 392860 385608
rect 369176 385568 369182 385580
rect 392854 385568 392860 385580
rect 392912 385568 392918 385620
rect 349062 385500 349068 385552
rect 349120 385540 349126 385552
rect 385862 385540 385868 385552
rect 349120 385512 385868 385540
rect 349120 385500 349126 385512
rect 385862 385500 385868 385512
rect 385920 385500 385926 385552
rect 355870 385432 355876 385484
rect 355928 385472 355934 385484
rect 399662 385472 399668 385484
rect 355928 385444 399668 385472
rect 355928 385432 355934 385444
rect 399662 385432 399668 385444
rect 399720 385432 399726 385484
rect 357342 385364 357348 385416
rect 357400 385404 357406 385416
rect 406654 385404 406660 385416
rect 357400 385376 406660 385404
rect 357400 385364 357406 385376
rect 406654 385364 406660 385376
rect 406712 385364 406718 385416
rect 353202 385296 353208 385348
rect 353260 385336 353266 385348
rect 402054 385336 402060 385348
rect 353260 385308 402060 385336
rect 353260 385296 353266 385308
rect 402054 385296 402060 385308
rect 402112 385296 402118 385348
rect 347682 385228 347688 385280
rect 347740 385268 347746 385280
rect 397454 385268 397460 385280
rect 347740 385240 397460 385268
rect 347740 385228 347746 385240
rect 397454 385228 397460 385240
rect 397512 385228 397518 385280
rect 343542 385160 343548 385212
rect 343600 385200 343606 385212
rect 395062 385200 395068 385212
rect 343600 385172 395068 385200
rect 343600 385160 343606 385172
rect 395062 385160 395068 385172
rect 395120 385160 395126 385212
rect 355962 385092 355968 385144
rect 356020 385132 356026 385144
rect 413462 385132 413468 385144
rect 356020 385104 413468 385132
rect 356020 385092 356026 385104
rect 413462 385092 413468 385104
rect 413520 385092 413526 385144
rect 367002 385024 367008 385076
rect 367060 385064 367066 385076
rect 390462 385064 390468 385076
rect 367060 385036 390468 385064
rect 367060 385024 367066 385036
rect 390462 385024 390468 385036
rect 390520 385024 390526 385076
rect 126514 384276 126520 384328
rect 126572 384316 126578 384328
rect 140774 384316 140780 384328
rect 126572 384288 140780 384316
rect 126572 384276 126578 384288
rect 140774 384276 140780 384288
rect 140832 384276 140838 384328
rect 126146 383664 126152 383716
rect 126204 383704 126210 383716
rect 126330 383704 126336 383716
rect 126204 383676 126336 383704
rect 126204 383664 126210 383676
rect 126330 383664 126336 383676
rect 126388 383664 126394 383716
rect 301590 381488 301596 381540
rect 301648 381528 301654 381540
rect 302142 381528 302148 381540
rect 301648 381500 302148 381528
rect 301648 381488 301654 381500
rect 302142 381488 302148 381500
rect 302200 381528 302206 381540
rect 380894 381528 380900 381540
rect 302200 381500 380900 381528
rect 302200 381488 302206 381500
rect 380894 381488 380900 381500
rect 380952 381488 380958 381540
rect 153286 379448 153292 379500
rect 153344 379488 153350 379500
rect 153470 379488 153476 379500
rect 153344 379460 153476 379488
rect 153344 379448 153350 379460
rect 153470 379448 153476 379460
rect 153528 379448 153534 379500
rect 304258 379352 304264 379364
rect 304219 379324 304264 379352
rect 304258 379312 304264 379324
rect 304316 379312 304322 379364
rect 132770 376796 132776 376848
rect 132828 376836 132834 376848
rect 132862 376836 132868 376848
rect 132828 376808 132868 376836
rect 132828 376796 132834 376808
rect 132862 376796 132868 376808
rect 132920 376796 132926 376848
rect 128817 376771 128875 376777
rect 128817 376737 128829 376771
rect 128863 376768 128875 376771
rect 128906 376768 128912 376780
rect 128863 376740 128912 376768
rect 128863 376737 128875 376740
rect 128817 376731 128875 376737
rect 128906 376728 128912 376740
rect 128964 376728 128970 376780
rect 299842 376728 299848 376780
rect 299900 376768 299906 376780
rect 299934 376768 299940 376780
rect 299900 376740 299940 376768
rect 299900 376728 299906 376740
rect 299934 376728 299940 376740
rect 299992 376728 299998 376780
rect 351822 376728 351828 376780
rect 351880 376768 351886 376780
rect 380894 376768 380900 376780
rect 351880 376740 380900 376768
rect 351880 376728 351886 376740
rect 380894 376728 380900 376740
rect 380952 376728 380958 376780
rect 132678 375340 132684 375352
rect 132639 375312 132684 375340
rect 132678 375300 132684 375312
rect 132736 375300 132742 375352
rect 126330 374116 126336 374128
rect 126164 374088 126336 374116
rect 126164 374060 126192 374088
rect 126330 374076 126336 374088
rect 126388 374076 126394 374128
rect 126146 374008 126152 374060
rect 126204 374008 126210 374060
rect 364242 374008 364248 374060
rect 364300 374048 364306 374060
rect 380894 374048 380900 374060
rect 364300 374020 380900 374048
rect 364300 374008 364306 374020
rect 380894 374008 380900 374020
rect 380952 374008 380958 374060
rect 416038 374008 416044 374060
rect 416096 374048 416102 374060
rect 456794 374048 456800 374060
rect 416096 374020 456800 374048
rect 416096 374008 416102 374020
rect 456794 374008 456800 374020
rect 456852 374008 456858 374060
rect 288342 372580 288348 372632
rect 288400 372620 288406 372632
rect 288526 372620 288532 372632
rect 288400 372592 288532 372620
rect 288400 372580 288406 372592
rect 288526 372580 288532 372592
rect 288584 372580 288590 372632
rect 288342 369900 288348 369912
rect 288303 369872 288348 369900
rect 288342 369860 288348 369872
rect 288400 369860 288406 369912
rect 304258 369900 304264 369912
rect 304184 369872 304264 369900
rect 304184 369844 304212 369872
rect 304258 369860 304264 369872
rect 304316 369860 304322 369912
rect 347590 369860 347596 369912
rect 347648 369900 347654 369912
rect 380894 369900 380900 369912
rect 347648 369872 380900 369900
rect 347648 369860 347654 369872
rect 380894 369860 380900 369872
rect 380952 369860 380958 369912
rect 304166 369792 304172 369844
rect 304224 369792 304230 369844
rect 133046 367004 133052 367056
rect 133104 367004 133110 367056
rect 133138 367004 133144 367056
rect 133196 367044 133202 367056
rect 153473 367047 153531 367053
rect 133196 367016 133241 367044
rect 133196 367004 133202 367016
rect 153473 367013 153485 367047
rect 153519 367044 153531 367047
rect 153562 367044 153568 367056
rect 153519 367016 153568 367044
rect 153519 367013 153531 367016
rect 153473 367007 153531 367013
rect 153562 367004 153568 367016
rect 153620 367004 153626 367056
rect 132681 366979 132739 366985
rect 132681 366945 132693 366979
rect 132727 366976 132739 366979
rect 132770 366976 132776 366988
rect 132727 366948 132776 366976
rect 132727 366945 132739 366948
rect 132681 366939 132739 366945
rect 132770 366936 132776 366948
rect 132828 366936 132834 366988
rect 132954 366868 132960 366920
rect 133012 366868 133018 366920
rect 132972 366784 133000 366868
rect 133064 366852 133092 367004
rect 133046 366800 133052 366852
rect 133104 366800 133110 366852
rect 132954 366732 132960 366784
rect 133012 366732 133018 366784
rect 2774 365712 2780 365764
rect 2832 365752 2838 365764
rect 5166 365752 5172 365764
rect 2832 365724 5172 365752
rect 2832 365712 2838 365724
rect 5166 365712 5172 365724
rect 5224 365712 5230 365764
rect 129366 365644 129372 365696
rect 129424 365684 129430 365696
rect 197722 365684 197728 365696
rect 129424 365656 197728 365684
rect 129424 365644 129430 365656
rect 197722 365644 197728 365656
rect 197780 365644 197786 365696
rect 126146 364352 126152 364404
rect 126204 364392 126210 364404
rect 126330 364392 126336 364404
rect 126204 364364 126336 364392
rect 126204 364352 126210 364364
rect 126330 364352 126336 364364
rect 126388 364352 126394 364404
rect 288342 362964 288348 362976
rect 288303 362936 288348 362964
rect 288342 362924 288348 362936
rect 288400 362924 288406 362976
rect 333882 362924 333888 362976
rect 333940 362964 333946 362976
rect 380894 362964 380900 362976
rect 333940 362936 380900 362964
rect 333940 362924 333946 362936
rect 380894 362924 380900 362936
rect 380952 362924 380958 362976
rect 132770 360204 132776 360256
rect 132828 360204 132834 360256
rect 288342 360244 288348 360256
rect 288303 360216 288348 360244
rect 288342 360204 288348 360216
rect 288400 360204 288406 360256
rect 304166 360204 304172 360256
rect 304224 360204 304230 360256
rect 132788 360120 132816 360204
rect 304184 360176 304212 360204
rect 304258 360176 304264 360188
rect 304184 360148 304264 360176
rect 304258 360136 304264 360148
rect 304316 360136 304322 360188
rect 132770 360068 132776 360120
rect 132828 360068 132834 360120
rect 133138 358680 133144 358692
rect 133099 358652 133144 358680
rect 133138 358640 133144 358652
rect 133196 358640 133202 358692
rect 153470 357456 153476 357468
rect 153431 357428 153476 357456
rect 153470 357416 153476 357428
rect 153528 357416 153534 357468
rect 144178 357348 144184 357400
rect 144236 357388 144242 357400
rect 145558 357388 145564 357400
rect 144236 357360 145564 357388
rect 144236 357348 144242 357360
rect 145558 357348 145564 357360
rect 145616 357348 145622 357400
rect 304258 357252 304264 357264
rect 304219 357224 304264 357252
rect 304258 357212 304264 357224
rect 304316 357212 304322 357264
rect 126330 354804 126336 354816
rect 126164 354776 126336 354804
rect 126164 354748 126192 354776
rect 126330 354764 126336 354776
rect 126388 354764 126394 354816
rect 126146 354696 126152 354748
rect 126204 354696 126210 354748
rect 288342 353308 288348 353320
rect 288303 353280 288348 353308
rect 288342 353268 288348 353280
rect 288400 353268 288406 353320
rect 354582 353268 354588 353320
rect 354640 353308 354646 353320
rect 380894 353308 380900 353320
rect 354640 353280 380900 353308
rect 354640 353268 354646 353280
rect 380894 353268 380900 353280
rect 380952 353268 380958 353320
rect 128998 351160 129004 351212
rect 129056 351200 129062 351212
rect 129826 351200 129832 351212
rect 129056 351172 129832 351200
rect 129056 351160 129062 351172
rect 129826 351160 129832 351172
rect 129884 351200 129890 351212
rect 130378 351200 130384 351212
rect 129884 351172 130384 351200
rect 129884 351160 129890 351172
rect 130378 351160 130384 351172
rect 130436 351160 130442 351212
rect 153470 350588 153476 350600
rect 153396 350560 153476 350588
rect 153396 350532 153424 350560
rect 153470 350548 153476 350560
rect 153528 350548 153534 350600
rect 153378 350480 153384 350532
rect 153436 350480 153442 350532
rect 299842 350480 299848 350532
rect 299900 350480 299906 350532
rect 299860 350452 299888 350480
rect 299934 350452 299940 350464
rect 299860 350424 299940 350452
rect 299934 350412 299940 350424
rect 299992 350412 299998 350464
rect 304258 347868 304264 347880
rect 304219 347840 304264 347868
rect 304258 347828 304264 347840
rect 304316 347828 304322 347880
rect 132678 347760 132684 347812
rect 132736 347800 132742 347812
rect 132862 347800 132868 347812
rect 132736 347772 132868 347800
rect 132736 347760 132742 347772
rect 132862 347760 132868 347772
rect 132920 347760 132926 347812
rect 381538 347692 381544 347744
rect 381596 347732 381602 347744
rect 386782 347732 386788 347744
rect 381596 347704 386788 347732
rect 381596 347692 381602 347704
rect 386782 347692 386788 347704
rect 386840 347692 386846 347744
rect 360102 347624 360108 347676
rect 360160 347664 360166 347676
rect 391382 347664 391388 347676
rect 360160 347636 391388 347664
rect 360160 347624 360166 347636
rect 391382 347624 391388 347636
rect 391440 347624 391446 347676
rect 362862 347556 362868 347608
rect 362920 347596 362926 347608
rect 398190 347596 398196 347608
rect 362920 347568 398196 347596
rect 362920 347556 362926 347568
rect 398190 347556 398196 347568
rect 398248 347556 398254 347608
rect 358722 347488 358728 347540
rect 358780 347528 358786 347540
rect 393590 347528 393596 347540
rect 358780 347500 393596 347528
rect 358780 347488 358786 347500
rect 393590 347488 393596 347500
rect 393648 347488 393654 347540
rect 362770 347420 362776 347472
rect 362828 347460 362834 347472
rect 402790 347460 402796 347472
rect 362828 347432 402796 347460
rect 362828 347420 362834 347432
rect 402790 347420 402796 347432
rect 402848 347420 402854 347472
rect 350442 347352 350448 347404
rect 350500 347392 350506 347404
rect 395982 347392 395988 347404
rect 350500 347364 395988 347392
rect 350500 347352 350506 347364
rect 395982 347352 395988 347364
rect 396040 347352 396046 347404
rect 342162 347284 342168 347336
rect 342220 347324 342226 347336
rect 388990 347324 388996 347336
rect 342220 347296 388996 347324
rect 342220 347284 342226 347296
rect 388990 347284 388996 347296
rect 389048 347284 389054 347336
rect 361482 347216 361488 347268
rect 361540 347256 361546 347268
rect 407390 347256 407396 347268
rect 361540 347228 407396 347256
rect 361540 347216 361546 347228
rect 407390 347216 407396 347228
rect 407448 347216 407454 347268
rect 354490 347148 354496 347200
rect 354548 347188 354554 347200
rect 400582 347188 400588 347200
rect 354548 347160 400588 347188
rect 354548 347148 354554 347160
rect 400582 347148 400588 347160
rect 400640 347148 400646 347200
rect 361390 347080 361396 347132
rect 361448 347120 361454 347132
rect 414382 347120 414388 347132
rect 361448 347092 414388 347120
rect 361448 347080 361454 347092
rect 414382 347080 414388 347092
rect 414440 347080 414446 347132
rect 333790 347012 333796 347064
rect 333848 347052 333854 347064
rect 411990 347052 411996 347064
rect 333848 347024 411996 347052
rect 333848 347012 333854 347024
rect 411990 347012 411996 347024
rect 412048 347012 412054 347064
rect 126146 345040 126152 345092
rect 126204 345080 126210 345092
rect 126330 345080 126336 345092
rect 126204 345052 126336 345080
rect 126204 345040 126210 345052
rect 126330 345040 126336 345052
rect 126388 345040 126394 345092
rect 504818 345040 504824 345092
rect 504876 345080 504882 345092
rect 579982 345080 579988 345092
rect 504876 345052 579988 345080
rect 504876 345040 504882 345052
rect 579982 345040 579988 345052
rect 580040 345040 580046 345092
rect 288161 344607 288219 344613
rect 288161 344573 288173 344607
rect 288207 344604 288219 344607
rect 288342 344604 288348 344616
rect 288207 344576 288348 344604
rect 288207 344573 288219 344576
rect 288161 344567 288219 344573
rect 288342 344564 288348 344576
rect 288400 344564 288406 344616
rect 128998 342864 129004 342916
rect 129056 342904 129062 342916
rect 130654 342904 130660 342916
rect 129056 342876 130660 342904
rect 129056 342864 129062 342876
rect 130654 342864 130660 342876
rect 130712 342904 130718 342916
rect 192478 342904 192484 342916
rect 130712 342876 192484 342904
rect 130712 342864 130718 342876
rect 192478 342864 192484 342876
rect 192536 342864 192542 342916
rect 199286 342864 199292 342916
rect 199344 342904 199350 342916
rect 200206 342904 200212 342916
rect 199344 342876 200212 342904
rect 199344 342864 199350 342876
rect 200206 342864 200212 342876
rect 200264 342864 200270 342916
rect 130286 342048 130292 342100
rect 130344 342088 130350 342100
rect 132678 342088 132684 342100
rect 130344 342060 132684 342088
rect 130344 342048 130350 342060
rect 132678 342048 132684 342060
rect 132736 342088 132742 342100
rect 132865 342091 132923 342097
rect 132865 342088 132877 342091
rect 132736 342060 132877 342088
rect 132736 342048 132742 342060
rect 132865 342057 132877 342060
rect 132911 342057 132923 342091
rect 132865 342051 132923 342057
rect 132494 341980 132500 342032
rect 132552 341980 132558 342032
rect 503806 341980 503812 342032
rect 503864 342020 503870 342032
rect 504174 342020 504180 342032
rect 503864 341992 504180 342020
rect 503864 341980 503870 341992
rect 504174 341980 504180 341992
rect 504232 341980 504238 342032
rect 132512 341896 132540 341980
rect 132494 341844 132500 341896
rect 132552 341844 132558 341896
rect 131942 341640 131948 341692
rect 132000 341680 132006 341692
rect 580626 341680 580632 341692
rect 132000 341652 580632 341680
rect 132000 341640 132006 341652
rect 580626 341640 580632 341652
rect 580684 341640 580690 341692
rect 132034 341572 132040 341624
rect 132092 341612 132098 341624
rect 580810 341612 580816 341624
rect 132092 341584 580816 341612
rect 132092 341572 132098 341584
rect 580810 341572 580816 341584
rect 580868 341572 580874 341624
rect 131666 341504 131672 341556
rect 131724 341544 131730 341556
rect 580718 341544 580724 341556
rect 131724 341516 580724 341544
rect 131724 341504 131730 341516
rect 580718 341504 580724 341516
rect 580776 341504 580782 341556
rect 153378 341000 153384 341012
rect 153339 340972 153384 341000
rect 153378 340960 153384 340972
rect 153436 340960 153442 341012
rect 127250 340824 127256 340876
rect 127308 340864 127314 340876
rect 408494 340864 408500 340876
rect 127308 340836 408500 340864
rect 127308 340824 127314 340836
rect 408494 340824 408500 340836
rect 408552 340824 408558 340876
rect 504726 340864 504732 340876
rect 504100 340836 504732 340864
rect 127158 340756 127164 340808
rect 127216 340796 127222 340808
rect 404354 340796 404360 340808
rect 127216 340768 404360 340796
rect 127216 340756 127222 340768
rect 404354 340756 404360 340768
rect 404412 340756 404418 340808
rect 503898 340756 503904 340808
rect 503956 340796 503962 340808
rect 504100 340796 504128 340836
rect 504726 340824 504732 340836
rect 504784 340824 504790 340876
rect 503956 340768 504128 340796
rect 503956 340756 503962 340768
rect 127710 340688 127716 340740
rect 127768 340728 127774 340740
rect 381722 340728 381728 340740
rect 127768 340700 381728 340728
rect 127768 340688 127774 340700
rect 381722 340688 381728 340700
rect 381780 340688 381786 340740
rect 130378 340620 130384 340672
rect 130436 340660 130442 340672
rect 381630 340660 381636 340672
rect 130436 340632 381636 340660
rect 130436 340620 130442 340632
rect 381630 340620 381636 340632
rect 381688 340620 381694 340672
rect 132862 340592 132868 340604
rect 132823 340564 132868 340592
rect 132862 340552 132868 340564
rect 132920 340552 132926 340604
rect 140774 340552 140780 340604
rect 140832 340592 140838 340604
rect 383654 340592 383660 340604
rect 140832 340564 383660 340592
rect 140832 340552 140838 340564
rect 383654 340552 383660 340564
rect 383712 340552 383718 340604
rect 145558 340484 145564 340536
rect 145616 340524 145622 340536
rect 381814 340524 381820 340536
rect 145616 340496 381820 340524
rect 145616 340484 145622 340496
rect 381814 340484 381820 340496
rect 381872 340484 381878 340536
rect 153378 340456 153384 340468
rect 153339 340428 153384 340456
rect 153378 340416 153384 340428
rect 153436 340416 153442 340468
rect 111702 340212 111708 340264
rect 111760 340252 111766 340264
rect 127250 340252 127256 340264
rect 111760 340224 127256 340252
rect 111760 340212 111766 340224
rect 127250 340212 127256 340224
rect 127308 340212 127314 340264
rect 110322 340144 110328 340196
rect 110380 340184 110386 340196
rect 127158 340184 127164 340196
rect 110380 340156 127164 340184
rect 110380 340144 110386 340156
rect 127158 340144 127164 340156
rect 127216 340144 127222 340196
rect 130746 340144 130752 340196
rect 130804 340184 130810 340196
rect 140774 340184 140780 340196
rect 130804 340156 140780 340184
rect 130804 340144 130810 340156
rect 140774 340144 140780 340156
rect 140832 340144 140838 340196
rect 130378 339668 130384 339720
rect 130436 339708 130442 339720
rect 130838 339708 130844 339720
rect 130436 339680 130844 339708
rect 130436 339668 130442 339680
rect 130838 339668 130844 339680
rect 130896 339668 130902 339720
rect 262122 339124 262128 339176
rect 262180 339164 262186 339176
rect 268930 339164 268936 339176
rect 262180 339136 268936 339164
rect 262180 339124 262186 339136
rect 268930 339124 268936 339136
rect 268988 339124 268994 339176
rect 198090 338988 198096 339040
rect 198148 339028 198154 339040
rect 209958 339028 209964 339040
rect 198148 339000 209964 339028
rect 198148 338988 198154 339000
rect 209958 338988 209964 339000
rect 210016 338988 210022 339040
rect 199470 338920 199476 338972
rect 199528 338960 199534 338972
rect 214098 338960 214104 338972
rect 199528 338932 214104 338960
rect 199528 338920 199534 338932
rect 214098 338920 214104 338932
rect 214156 338920 214162 338972
rect 257706 338920 257712 338972
rect 257764 338960 257770 338972
rect 267550 338960 267556 338972
rect 257764 338932 267556 338960
rect 257764 338920 257770 338932
rect 267550 338920 267556 338932
rect 267608 338920 267614 338972
rect 199378 338852 199384 338904
rect 199436 338892 199442 338904
rect 215294 338892 215300 338904
rect 199436 338864 215300 338892
rect 199436 338852 199442 338864
rect 215294 338852 215300 338864
rect 215352 338852 215358 338904
rect 253658 338852 253664 338904
rect 253716 338892 253722 338904
rect 268838 338892 268844 338904
rect 253716 338864 268844 338892
rect 253716 338852 253722 338864
rect 268838 338852 268844 338864
rect 268896 338852 268902 338904
rect 198274 338784 198280 338836
rect 198332 338824 198338 338836
rect 220814 338824 220820 338836
rect 198332 338796 220820 338824
rect 198332 338784 198338 338796
rect 220814 338784 220820 338796
rect 220872 338784 220878 338836
rect 244182 338784 244188 338836
rect 244240 338824 244246 338836
rect 268746 338824 268752 338836
rect 244240 338796 268752 338824
rect 244240 338784 244246 338796
rect 268746 338784 268752 338796
rect 268804 338784 268810 338836
rect 198182 338716 198188 338768
rect 198240 338756 198246 338768
rect 222194 338756 222200 338768
rect 198240 338728 222200 338756
rect 198240 338716 198246 338728
rect 222194 338716 222200 338728
rect 222252 338716 222258 338768
rect 237282 338716 237288 338768
rect 237340 338756 237346 338768
rect 267642 338756 267648 338768
rect 237340 338728 267648 338756
rect 237340 338716 237346 338728
rect 267642 338716 267648 338728
rect 267700 338716 267706 338768
rect 128906 338104 128912 338156
rect 128964 338144 128970 338156
rect 128998 338144 129004 338156
rect 128964 338116 129004 338144
rect 128964 338104 128970 338116
rect 128998 338104 129004 338116
rect 129056 338104 129062 338156
rect 288161 338147 288219 338153
rect 288161 338113 288173 338147
rect 288207 338144 288219 338147
rect 288342 338144 288348 338156
rect 288207 338116 288348 338144
rect 288207 338113 288219 338116
rect 288161 338107 288219 338113
rect 288342 338104 288348 338116
rect 288400 338104 288406 338156
rect 107562 338036 107568 338088
rect 107620 338076 107626 338088
rect 301590 338076 301596 338088
rect 107620 338048 301596 338076
rect 107620 338036 107626 338048
rect 301590 338036 301596 338048
rect 301648 338036 301654 338088
rect 97902 337968 97908 338020
rect 97960 338008 97966 338020
rect 126974 338008 126980 338020
rect 97960 337980 126980 338008
rect 97960 337968 97966 337980
rect 126974 337968 126980 337980
rect 127032 337968 127038 338020
rect 132954 337968 132960 338020
rect 133012 337968 133018 338020
rect 133046 337968 133052 338020
rect 133104 337968 133110 338020
rect 133138 337968 133144 338020
rect 133196 338008 133202 338020
rect 133196 337980 133241 338008
rect 133196 337968 133202 337980
rect 220446 337968 220452 338020
rect 220504 338008 220510 338020
rect 238110 338008 238116 338020
rect 220504 337980 238116 338008
rect 220504 337968 220510 337980
rect 238110 337968 238116 337980
rect 238168 337968 238174 338020
rect 241333 338011 241391 338017
rect 241333 337977 241345 338011
rect 241379 338008 241391 338011
rect 244918 338008 244924 338020
rect 241379 337980 244924 338008
rect 241379 337977 241391 337980
rect 241333 337971 241391 337977
rect 244918 337968 244924 337980
rect 244976 337968 244982 338020
rect 112806 337900 112812 337952
rect 112864 337940 112870 337952
rect 113082 337940 113088 337952
rect 112864 337912 113088 337940
rect 112864 337900 112870 337912
rect 113082 337900 113088 337912
rect 113140 337940 113146 337952
rect 127066 337940 127072 337952
rect 113140 337912 127072 337940
rect 113140 337900 113146 337912
rect 127066 337900 127072 337912
rect 127124 337900 127130 337952
rect 132972 337884 133000 337968
rect 133064 337884 133092 337968
rect 209038 337900 209044 337952
rect 209096 337940 209102 337952
rect 220078 337940 220084 337952
rect 209096 337912 220084 337940
rect 209096 337900 209102 337912
rect 220078 337900 220084 337912
rect 220136 337900 220142 337952
rect 226150 337900 226156 337952
rect 226208 337940 226214 337952
rect 248690 337940 248696 337952
rect 226208 337912 248696 337940
rect 226208 337900 226214 337912
rect 248690 337900 248696 337912
rect 248748 337900 248754 337952
rect 250990 337900 250996 337952
rect 251048 337940 251054 337952
rect 260190 337940 260196 337952
rect 251048 337912 260196 337940
rect 251048 337900 251054 337912
rect 260190 337900 260196 337912
rect 260248 337900 260254 337952
rect 122742 337832 122748 337884
rect 122800 337872 122806 337884
rect 127710 337872 127716 337884
rect 122800 337844 127716 337872
rect 122800 337832 122806 337844
rect 127710 337832 127716 337844
rect 127768 337832 127774 337884
rect 132954 337832 132960 337884
rect 133012 337832 133018 337884
rect 133046 337832 133052 337884
rect 133104 337832 133110 337884
rect 203334 337832 203340 337884
rect 203392 337872 203398 337884
rect 215938 337872 215944 337884
rect 203392 337844 215944 337872
rect 203392 337832 203398 337844
rect 215938 337832 215944 337844
rect 215996 337832 216002 337884
rect 217502 337832 217508 337884
rect 217560 337872 217566 337884
rect 241333 337875 241391 337881
rect 241333 337872 241345 337875
rect 217560 337844 241345 337872
rect 217560 337832 217566 337844
rect 241333 337841 241345 337844
rect 241379 337841 241391 337875
rect 241333 337835 241391 337841
rect 241422 337832 241428 337884
rect 241480 337872 241486 337884
rect 246022 337872 246028 337884
rect 241480 337844 246028 337872
rect 241480 337832 241486 337844
rect 246022 337832 246028 337844
rect 246080 337832 246086 337884
rect 253750 337832 253756 337884
rect 253808 337872 253814 337884
rect 263134 337872 263140 337884
rect 253808 337844 263140 337872
rect 253808 337832 253814 337844
rect 263134 337832 263140 337844
rect 263192 337832 263198 337884
rect 200574 337764 200580 337816
rect 200632 337804 200638 337816
rect 233513 337807 233571 337813
rect 233513 337804 233525 337807
rect 200632 337776 233525 337804
rect 200632 337764 200638 337776
rect 233513 337773 233525 337776
rect 233559 337773 233571 337807
rect 233513 337767 233571 337773
rect 234614 337764 234620 337816
rect 234672 337804 234678 337816
rect 237742 337804 237748 337816
rect 234672 337776 237748 337804
rect 234672 337764 234678 337776
rect 237742 337764 237748 337776
rect 237800 337764 237806 337816
rect 240042 337764 240048 337816
rect 240100 337804 240106 337816
rect 243078 337804 243084 337816
rect 240100 337776 243084 337804
rect 240100 337764 240106 337776
rect 243078 337764 243084 337776
rect 243136 337764 243142 337816
rect 247678 337764 247684 337816
rect 247736 337804 247742 337816
rect 257430 337804 257436 337816
rect 247736 337776 257436 337804
rect 247736 337764 247742 337776
rect 257430 337764 257436 337776
rect 257488 337764 257494 337816
rect 92750 337696 92756 337748
rect 92808 337736 92814 337748
rect 93762 337736 93768 337748
rect 92808 337708 93768 337736
rect 92808 337696 92814 337708
rect 93762 337696 93768 337708
rect 93820 337696 93826 337748
rect 102870 337696 102876 337748
rect 102928 337736 102934 337748
rect 103422 337736 103428 337748
rect 102928 337708 103428 337736
rect 102928 337696 102934 337708
rect 103422 337696 103428 337708
rect 103480 337696 103486 337748
rect 214742 337696 214748 337748
rect 214800 337736 214806 337748
rect 258718 337736 258724 337748
rect 214800 337708 258724 337736
rect 214800 337696 214806 337708
rect 258718 337696 258724 337708
rect 258776 337696 258782 337748
rect 206094 337628 206100 337680
rect 206152 337668 206158 337680
rect 251637 337671 251695 337677
rect 251637 337668 251649 337671
rect 206152 337640 251649 337668
rect 206152 337628 206158 337640
rect 251637 337637 251649 337640
rect 251683 337637 251695 337671
rect 251637 337631 251695 337637
rect 251726 337628 251732 337680
rect 251784 337668 251790 337680
rect 252462 337668 252468 337680
rect 251784 337640 252468 337668
rect 251784 337628 251790 337640
rect 252462 337628 252468 337640
rect 252520 337628 252526 337680
rect 72878 337560 72884 337612
rect 72936 337600 72942 337612
rect 134058 337600 134064 337612
rect 72936 337572 134064 337600
rect 72936 337560 72942 337572
rect 134058 337560 134064 337572
rect 134116 337600 134122 337612
rect 299934 337600 299940 337612
rect 134116 337572 299940 337600
rect 134116 337560 134122 337572
rect 299934 337560 299940 337572
rect 299992 337560 299998 337612
rect 401502 337560 401508 337612
rect 401560 337600 401566 337612
rect 460566 337600 460572 337612
rect 401560 337572 460572 337600
rect 401560 337560 401566 337572
rect 460566 337560 460572 337572
rect 460624 337560 460630 337612
rect 117958 337492 117964 337544
rect 118016 337532 118022 337544
rect 124122 337532 124128 337544
rect 118016 337504 124128 337532
rect 118016 337492 118022 337504
rect 124122 337492 124128 337504
rect 124180 337532 124186 337544
rect 297358 337532 297364 337544
rect 124180 337504 297364 337532
rect 124180 337492 124186 337504
rect 297358 337492 297364 337504
rect 297416 337492 297422 337544
rect 411162 337492 411168 337544
rect 411220 337532 411226 337544
rect 472158 337532 472164 337544
rect 411220 337504 472164 337532
rect 411220 337492 411226 337504
rect 472158 337492 472164 337504
rect 472216 337492 472222 337544
rect 77846 337424 77852 337476
rect 77904 337464 77910 337476
rect 99282 337464 99288 337476
rect 77904 337436 99288 337464
rect 77904 337424 77910 337436
rect 99282 337424 99288 337436
rect 99340 337464 99346 337476
rect 329834 337464 329840 337476
rect 99340 337436 329840 337464
rect 99340 337424 99346 337436
rect 329834 337424 329840 337436
rect 329892 337424 329898 337476
rect 408402 337424 408408 337476
rect 408460 337464 408466 337476
rect 483750 337464 483756 337476
rect 408460 337436 483756 337464
rect 408460 337424 408466 337436
rect 483750 337424 483756 337436
rect 483808 337424 483814 337476
rect 87782 337356 87788 337408
rect 87840 337396 87846 337408
rect 128262 337396 128268 337408
rect 87840 337368 128268 337396
rect 87840 337356 87846 337368
rect 128262 337356 128268 337368
rect 128320 337396 128326 337408
rect 380526 337396 380532 337408
rect 128320 337368 380532 337396
rect 128320 337356 128326 337368
rect 380526 337356 380532 337368
rect 380584 337356 380590 337408
rect 413922 337356 413928 337408
rect 413980 337396 413986 337408
rect 495342 337396 495348 337408
rect 413980 337368 495348 337396
rect 413980 337356 413986 337368
rect 495342 337356 495348 337368
rect 495400 337356 495406 337408
rect 231854 337288 231860 337340
rect 231912 337328 231918 337340
rect 248782 337328 248788 337340
rect 231912 337300 248788 337328
rect 231912 337288 231918 337300
rect 248782 337288 248788 337300
rect 248840 337288 248846 337340
rect 251637 337331 251695 337337
rect 251637 337297 251649 337331
rect 251683 337328 251695 337331
rect 255314 337328 255320 337340
rect 251683 337300 255320 337328
rect 251683 337297 251695 337300
rect 251637 337291 251695 337297
rect 255314 337288 255320 337300
rect 255372 337288 255378 337340
rect 228910 337220 228916 337272
rect 228968 337260 228974 337272
rect 232498 337260 232504 337272
rect 228968 337232 232504 337260
rect 228968 337220 228974 337232
rect 232498 337220 232504 337232
rect 232556 337220 232562 337272
rect 237558 337220 237564 337272
rect 237616 337260 237622 337272
rect 243078 337260 243084 337272
rect 237616 337232 243084 337260
rect 237616 337220 237622 337232
rect 243078 337220 243084 337232
rect 243136 337220 243142 337272
rect 233513 337195 233571 337201
rect 233513 337161 233525 337195
rect 233559 337192 233571 337195
rect 238018 337192 238024 337204
rect 233559 337164 238024 337192
rect 233559 337161 233571 337164
rect 233513 337155 233571 337161
rect 238018 337152 238024 337164
rect 238076 337152 238082 337204
rect 223206 336812 223212 336864
rect 223264 336852 223270 336864
rect 229738 336852 229744 336864
rect 223264 336824 229744 336852
rect 223264 336812 223270 336824
rect 229738 336812 229744 336824
rect 229796 336812 229802 336864
rect 244090 336812 244096 336864
rect 244148 336852 244154 336864
rect 248598 336852 248604 336864
rect 244148 336824 248604 336852
rect 244148 336812 244154 336824
rect 248598 336812 248604 336824
rect 248656 336812 248662 336864
rect 254486 336812 254492 336864
rect 254544 336852 254550 336864
rect 258258 336852 258264 336864
rect 254544 336824 258264 336852
rect 254544 336812 254550 336824
rect 258258 336812 258264 336824
rect 258316 336812 258322 336864
rect 2958 336744 2964 336796
rect 3016 336784 3022 336796
rect 434898 336784 434904 336796
rect 3016 336756 434904 336784
rect 3016 336744 3022 336756
rect 434898 336744 434904 336756
rect 434956 336744 434962 336796
rect 82722 336676 82728 336728
rect 82780 336716 82786 336728
rect 125870 336716 125876 336728
rect 82780 336688 125876 336716
rect 82780 336676 82786 336688
rect 125870 336676 125876 336688
rect 125928 336676 125934 336728
rect 257706 336676 257712 336728
rect 257764 336716 257770 336728
rect 257798 336716 257804 336728
rect 257764 336688 257804 336716
rect 257764 336676 257770 336688
rect 257798 336676 257804 336688
rect 257856 336676 257862 336728
rect 126146 335316 126152 335368
rect 126204 335356 126210 335368
rect 126330 335356 126336 335368
rect 126204 335328 126336 335356
rect 126204 335316 126210 335328
rect 126330 335316 126336 335328
rect 126388 335316 126394 335368
rect 257709 335291 257767 335297
rect 257709 335257 257721 335291
rect 257755 335288 257767 335291
rect 257798 335288 257804 335300
rect 257755 335260 257804 335288
rect 257755 335257 257767 335260
rect 257709 335251 257767 335257
rect 257798 335248 257804 335260
rect 257856 335248 257862 335300
rect 133138 333316 133144 333328
rect 133099 333288 133144 333316
rect 133138 333276 133144 333288
rect 133196 333276 133202 333328
rect 288342 332024 288348 332036
rect 288303 331996 288348 332024
rect 288342 331984 288348 331996
rect 288400 331984 288406 332036
rect 213917 331347 213975 331353
rect 213917 331313 213929 331347
rect 213963 331344 213975 331347
rect 214006 331344 214012 331356
rect 213963 331316 214012 331344
rect 213963 331313 213975 331316
rect 213917 331307 213975 331313
rect 214006 331304 214012 331316
rect 214064 331304 214070 331356
rect 503717 331279 503775 331285
rect 503717 331245 503729 331279
rect 503763 331276 503775 331279
rect 503806 331276 503812 331288
rect 503763 331248 503812 331276
rect 503763 331245 503775 331248
rect 503717 331239 503775 331245
rect 503806 331236 503812 331248
rect 503864 331236 503870 331288
rect 503622 331168 503628 331220
rect 503680 331208 503686 331220
rect 503990 331208 503996 331220
rect 503680 331180 503996 331208
rect 503680 331168 503686 331180
rect 503990 331168 503996 331180
rect 504048 331168 504054 331220
rect 503714 328556 503720 328568
rect 503675 328528 503720 328556
rect 503714 328516 503720 328528
rect 503772 328516 503778 328568
rect 209774 328448 209780 328500
rect 209832 328488 209838 328500
rect 209958 328488 209964 328500
rect 209832 328460 209964 328488
rect 209832 328448 209838 328460
rect 209958 328448 209964 328460
rect 210016 328448 210022 328500
rect 213914 328488 213920 328500
rect 213875 328460 213920 328488
rect 213914 328448 213920 328460
rect 213972 328448 213978 328500
rect 288158 328448 288164 328500
rect 288216 328488 288222 328500
rect 288345 328491 288403 328497
rect 288345 328488 288357 328491
rect 288216 328460 288357 328488
rect 288216 328448 288222 328460
rect 288345 328457 288357 328460
rect 288391 328457 288403 328491
rect 288345 328451 288403 328457
rect 128998 328420 129004 328432
rect 128959 328392 129004 328420
rect 128998 328380 129004 328392
rect 129056 328380 129062 328432
rect 504266 328380 504272 328432
rect 504324 328420 504330 328432
rect 504358 328420 504364 328432
rect 504324 328392 504364 328420
rect 504324 328380 504330 328392
rect 504358 328380 504364 328392
rect 504416 328380 504422 328432
rect 288158 328352 288164 328364
rect 288119 328324 288164 328352
rect 288158 328312 288164 328324
rect 288216 328312 288222 328364
rect 504266 327060 504272 327072
rect 504227 327032 504272 327060
rect 504266 327020 504272 327032
rect 504324 327020 504330 327072
rect 126146 325660 126152 325712
rect 126204 325700 126210 325712
rect 126330 325700 126336 325712
rect 126204 325672 126336 325700
rect 126204 325660 126210 325672
rect 126330 325660 126336 325672
rect 126388 325660 126394 325712
rect 503898 321716 503904 321768
rect 503956 321756 503962 321768
rect 503956 321728 504001 321756
rect 503956 321716 503962 321728
rect 503714 321688 503720 321700
rect 503675 321660 503720 321688
rect 503714 321648 503720 321660
rect 503772 321648 503778 321700
rect 503990 321688 503996 321700
rect 503951 321660 503996 321688
rect 503990 321648 503996 321660
rect 504048 321648 504054 321700
rect 132770 321580 132776 321632
rect 132828 321620 132834 321632
rect 579614 321620 579620 321632
rect 132828 321592 579620 321620
rect 132828 321580 132834 321592
rect 579614 321580 579620 321592
rect 579672 321580 579678 321632
rect 503898 321552 503904 321564
rect 503859 321524 503904 321552
rect 503898 321512 503904 321524
rect 503956 321512 503962 321564
rect 128814 318860 128820 318912
rect 128872 318900 128878 318912
rect 129001 318903 129059 318909
rect 129001 318900 129013 318903
rect 128872 318872 129013 318900
rect 128872 318860 128878 318872
rect 129001 318869 129013 318872
rect 129047 318869 129059 318903
rect 129001 318863 129059 318869
rect 153378 318792 153384 318844
rect 153436 318832 153442 318844
rect 153470 318832 153476 318844
rect 153436 318804 153476 318832
rect 153436 318792 153442 318804
rect 153470 318792 153476 318804
rect 153528 318792 153534 318844
rect 288161 318835 288219 318841
rect 288161 318801 288173 318835
rect 288207 318832 288219 318835
rect 288342 318832 288348 318844
rect 288207 318804 288348 318832
rect 288207 318801 288219 318804
rect 288161 318795 288219 318801
rect 288342 318792 288348 318804
rect 288400 318792 288406 318844
rect 503990 318832 503996 318844
rect 503951 318804 503996 318832
rect 503990 318792 503996 318804
rect 504048 318792 504054 318844
rect 209774 318764 209780 318776
rect 209735 318736 209780 318764
rect 209774 318724 209780 318736
rect 209832 318724 209838 318776
rect 304258 318764 304264 318776
rect 304219 318736 304264 318764
rect 304258 318724 304264 318736
rect 304316 318724 304322 318776
rect 257706 317472 257712 317484
rect 257667 317444 257712 317472
rect 257706 317432 257712 317444
rect 257764 317432 257770 317484
rect 503714 317472 503720 317484
rect 503675 317444 503720 317472
rect 503714 317432 503720 317444
rect 503772 317432 503778 317484
rect 504269 317475 504327 317481
rect 504269 317441 504281 317475
rect 504315 317472 504327 317475
rect 504358 317472 504364 317484
rect 504315 317444 504364 317472
rect 504315 317441 504327 317444
rect 504269 317435 504327 317441
rect 504358 317432 504364 317444
rect 504416 317432 504422 317484
rect 128633 317407 128691 317413
rect 128633 317373 128645 317407
rect 128679 317404 128691 317407
rect 128906 317404 128912 317416
rect 128679 317376 128912 317404
rect 128679 317373 128691 317376
rect 128633 317367 128691 317373
rect 128906 317364 128912 317376
rect 128964 317364 128970 317416
rect 126146 316004 126152 316056
rect 126204 316044 126210 316056
rect 126330 316044 126336 316056
rect 126204 316016 126336 316044
rect 126204 316004 126210 316016
rect 126330 316004 126336 316016
rect 126388 316004 126394 316056
rect 288342 313392 288348 313404
rect 288303 313364 288348 313392
rect 288342 313352 288348 313364
rect 288400 313352 288406 313404
rect 504358 312644 504364 312656
rect 504319 312616 504364 312644
rect 504358 312604 504364 312616
rect 504416 312604 504422 312656
rect 153378 311924 153384 311976
rect 153436 311964 153442 311976
rect 153470 311964 153476 311976
rect 153436 311936 153476 311964
rect 153436 311924 153442 311936
rect 153470 311924 153476 311936
rect 153528 311924 153534 311976
rect 503622 311856 503628 311908
rect 503680 311896 503686 311908
rect 503990 311896 503996 311908
rect 503680 311868 503996 311896
rect 503680 311856 503686 311868
rect 503990 311856 503996 311868
rect 504048 311856 504054 311908
rect 503622 311720 503628 311772
rect 503680 311760 503686 311772
rect 503990 311760 503996 311772
rect 503680 311732 503996 311760
rect 503680 311720 503686 311732
rect 503990 311720 503996 311732
rect 504048 311720 504054 311772
rect 131850 310496 131856 310548
rect 131908 310536 131914 310548
rect 579706 310536 579712 310548
rect 131908 310508 579712 310536
rect 131908 310496 131914 310508
rect 579706 310496 579712 310508
rect 579764 310496 579770 310548
rect 304258 309244 304264 309256
rect 304219 309216 304264 309244
rect 304258 309204 304264 309216
rect 304316 309204 304322 309256
rect 209774 309176 209780 309188
rect 209735 309148 209780 309176
rect 209774 309136 209780 309148
rect 209832 309136 209838 309188
rect 288342 309176 288348 309188
rect 288303 309148 288348 309176
rect 288342 309136 288348 309148
rect 288400 309136 288406 309188
rect 304258 309108 304264 309120
rect 304219 309080 304264 309108
rect 304258 309068 304264 309080
rect 304316 309068 304322 309120
rect 132678 308252 132684 308304
rect 132736 308292 132742 308304
rect 132862 308292 132868 308304
rect 132736 308264 132868 308292
rect 132736 308252 132742 308264
rect 132862 308252 132868 308264
rect 132920 308252 132926 308304
rect 4062 307776 4068 307828
rect 4120 307816 4126 307828
rect 5258 307816 5264 307828
rect 4120 307788 5264 307816
rect 4120 307776 4126 307788
rect 5258 307776 5264 307788
rect 5316 307776 5322 307828
rect 128630 307816 128636 307828
rect 128591 307788 128636 307816
rect 128630 307776 128636 307788
rect 128688 307776 128694 307828
rect 257798 307748 257804 307760
rect 257759 307720 257804 307748
rect 257798 307708 257804 307720
rect 257856 307708 257862 307760
rect 153286 302200 153292 302252
rect 153344 302240 153350 302252
rect 153470 302240 153476 302252
rect 153344 302212 153476 302240
rect 153344 302200 153350 302212
rect 153470 302200 153476 302212
rect 153528 302200 153534 302252
rect 288342 302240 288348 302252
rect 288303 302212 288348 302240
rect 288342 302200 288348 302212
rect 288400 302200 288406 302252
rect 128630 302064 128636 302116
rect 128688 302104 128694 302116
rect 128906 302104 128912 302116
rect 128688 302076 128912 302104
rect 128688 302064 128694 302076
rect 128906 302064 128912 302076
rect 128964 302064 128970 302116
rect 304258 301696 304264 301708
rect 304219 301668 304264 301696
rect 304258 301656 304264 301668
rect 304316 301656 304322 301708
rect 288342 299520 288348 299532
rect 288303 299492 288348 299520
rect 288342 299480 288348 299492
rect 288400 299480 288406 299532
rect 503622 299480 503628 299532
rect 503680 299520 503686 299532
rect 503806 299520 503812 299532
rect 503680 299492 503812 299520
rect 503680 299480 503686 299492
rect 503806 299480 503812 299492
rect 503864 299480 503870 299532
rect 504361 299523 504419 299529
rect 504361 299489 504373 299523
rect 504407 299520 504419 299523
rect 504450 299520 504456 299532
rect 504407 299492 504456 299520
rect 504407 299489 504419 299492
rect 504361 299483 504419 299489
rect 504450 299480 504456 299492
rect 504508 299480 504514 299532
rect 209774 299452 209780 299464
rect 209735 299424 209780 299452
rect 209774 299412 209780 299424
rect 209832 299412 209838 299464
rect 304258 299452 304264 299464
rect 304219 299424 304264 299452
rect 304258 299412 304264 299424
rect 304316 299412 304322 299464
rect 257801 298163 257859 298169
rect 257801 298129 257813 298163
rect 257847 298160 257859 298163
rect 257890 298160 257896 298172
rect 257847 298132 257896 298160
rect 257847 298129 257859 298132
rect 257801 298123 257859 298129
rect 257890 298120 257896 298132
rect 257948 298120 257954 298172
rect 504450 298092 504456 298104
rect 504411 298064 504456 298092
rect 504450 298052 504456 298064
rect 504508 298052 504514 298104
rect 126146 296692 126152 296744
rect 126204 296732 126210 296744
rect 126330 296732 126336 296744
rect 126204 296704 126336 296732
rect 126204 296692 126210 296704
rect 126330 296692 126336 296704
rect 126388 296692 126394 296744
rect 132678 296080 132684 296132
rect 132736 296120 132742 296132
rect 132862 296120 132868 296132
rect 132736 296092 132868 296120
rect 132736 296080 132742 296092
rect 132862 296080 132868 296092
rect 132920 296080 132926 296132
rect 288342 294080 288348 294092
rect 288303 294052 288348 294080
rect 288342 294040 288348 294052
rect 288400 294040 288406 294092
rect 3326 293972 3332 294024
rect 3384 294012 3390 294024
rect 434530 294012 434536 294024
rect 3384 293984 434536 294012
rect 3384 293972 3390 293984
rect 434530 293972 434536 293984
rect 434588 293972 434594 294024
rect 126054 292476 126060 292528
rect 126112 292516 126118 292528
rect 126330 292516 126336 292528
rect 126112 292488 126336 292516
rect 126112 292476 126118 292488
rect 126330 292476 126336 292488
rect 126388 292476 126394 292528
rect 304258 289932 304264 289944
rect 304219 289904 304264 289932
rect 304258 289892 304264 289904
rect 304316 289892 304322 289944
rect 209774 289864 209780 289876
rect 209735 289836 209780 289864
rect 209774 289824 209780 289836
rect 209832 289824 209838 289876
rect 288158 289824 288164 289876
rect 288216 289864 288222 289876
rect 288345 289867 288403 289873
rect 288345 289864 288357 289867
rect 288216 289836 288357 289864
rect 288216 289824 288222 289836
rect 288345 289833 288357 289836
rect 288391 289833 288403 289867
rect 288345 289827 288403 289833
rect 128814 289796 128820 289808
rect 128775 289768 128820 289796
rect 128814 289756 128820 289768
rect 128872 289756 128878 289808
rect 304258 289796 304264 289808
rect 304219 289768 304264 289796
rect 304258 289756 304264 289768
rect 304316 289756 304322 289808
rect 288158 289728 288164 289740
rect 288119 289700 288164 289728
rect 288158 289688 288164 289700
rect 288216 289688 288222 289740
rect 132678 288940 132684 288992
rect 132736 288980 132742 288992
rect 132862 288980 132868 288992
rect 132736 288952 132868 288980
rect 132736 288940 132742 288952
rect 132862 288940 132868 288952
rect 132920 288940 132926 288992
rect 257798 288396 257804 288448
rect 257856 288436 257862 288448
rect 257890 288436 257896 288448
rect 257856 288408 257896 288436
rect 257856 288396 257862 288408
rect 257890 288396 257896 288408
rect 257948 288396 257954 288448
rect 504453 288439 504511 288445
rect 504453 288405 504465 288439
rect 504499 288436 504511 288439
rect 504542 288436 504548 288448
rect 504499 288408 504548 288436
rect 504499 288405 504511 288408
rect 504453 288399 504511 288405
rect 504542 288396 504548 288408
rect 504600 288396 504606 288448
rect 257798 288300 257804 288312
rect 257759 288272 257804 288300
rect 257798 288260 257804 288272
rect 257856 288260 257862 288312
rect 503714 283024 503720 283076
rect 503772 283064 503778 283076
rect 503772 283036 503852 283064
rect 503772 283024 503778 283036
rect 503824 283008 503852 283036
rect 503806 282956 503812 283008
rect 503864 282956 503870 283008
rect 153286 282888 153292 282940
rect 153344 282928 153350 282940
rect 153470 282928 153476 282940
rect 153344 282900 153476 282928
rect 153344 282888 153350 282900
rect 153470 282888 153476 282900
rect 153528 282888 153534 282940
rect 304258 282792 304264 282804
rect 304219 282764 304264 282792
rect 304258 282752 304264 282764
rect 304316 282752 304322 282804
rect 128817 280211 128875 280217
rect 128817 280177 128829 280211
rect 128863 280208 128875 280211
rect 128906 280208 128912 280220
rect 128863 280180 128912 280208
rect 128863 280177 128875 280180
rect 128817 280171 128875 280177
rect 128906 280168 128912 280180
rect 128964 280168 128970 280220
rect 288161 280211 288219 280217
rect 288161 280177 288173 280211
rect 288207 280208 288219 280211
rect 288342 280208 288348 280220
rect 288207 280180 288348 280208
rect 288207 280177 288219 280180
rect 288161 280171 288219 280177
rect 288342 280168 288348 280180
rect 288400 280168 288406 280220
rect 126057 280143 126115 280149
rect 126057 280109 126069 280143
rect 126103 280140 126115 280143
rect 126146 280140 126152 280152
rect 126103 280112 126152 280140
rect 126103 280109 126115 280112
rect 126057 280103 126115 280109
rect 126146 280100 126152 280112
rect 126204 280100 126210 280152
rect 153378 280140 153384 280152
rect 153339 280112 153384 280140
rect 153378 280100 153384 280112
rect 153436 280100 153442 280152
rect 209774 280140 209780 280152
rect 209735 280112 209780 280140
rect 209774 280100 209780 280112
rect 209832 280100 209838 280152
rect 304258 280140 304264 280152
rect 304219 280112 304264 280140
rect 304258 280100 304264 280112
rect 304316 280100 304322 280152
rect 257801 278783 257859 278789
rect 257801 278749 257813 278783
rect 257847 278780 257859 278783
rect 257890 278780 257896 278792
rect 257847 278752 257896 278780
rect 257847 278749 257859 278752
rect 257801 278743 257859 278749
rect 257890 278740 257896 278752
rect 257948 278740 257954 278792
rect 504450 278712 504456 278724
rect 504411 278684 504456 278712
rect 504450 278672 504456 278684
rect 504508 278672 504514 278724
rect 132862 278060 132868 278112
rect 132920 278100 132926 278112
rect 133506 278100 133512 278112
rect 132920 278072 133512 278100
rect 132920 278060 132926 278072
rect 133506 278060 133512 278072
rect 133564 278060 133570 278112
rect 288342 274768 288348 274780
rect 288303 274740 288348 274768
rect 288342 274728 288348 274740
rect 288400 274728 288406 274780
rect 132678 274660 132684 274712
rect 132736 274700 132742 274712
rect 579614 274700 579620 274712
rect 132736 274672 579620 274700
rect 132736 274660 132742 274672
rect 579614 274660 579620 274672
rect 579672 274660 579678 274712
rect 503622 273300 503628 273352
rect 503680 273340 503686 273352
rect 503990 273340 503996 273352
rect 503680 273312 503996 273340
rect 503680 273300 503686 273312
rect 503990 273300 503996 273312
rect 504048 273300 504054 273352
rect 153381 273275 153439 273281
rect 153381 273241 153393 273275
rect 153427 273272 153439 273275
rect 153562 273272 153568 273284
rect 153427 273244 153568 273272
rect 153427 273241 153439 273244
rect 153381 273235 153439 273241
rect 153562 273232 153568 273244
rect 153620 273232 153626 273284
rect 503622 273164 503628 273216
rect 503680 273204 503686 273216
rect 503990 273204 503996 273216
rect 503680 273176 503996 273204
rect 503680 273164 503686 273176
rect 503990 273164 503996 273176
rect 504048 273164 504054 273216
rect 304258 270620 304264 270632
rect 304219 270592 304264 270620
rect 304258 270580 304264 270592
rect 304316 270580 304322 270632
rect 126054 270552 126060 270564
rect 126015 270524 126060 270552
rect 126054 270512 126060 270524
rect 126112 270512 126118 270564
rect 209774 270552 209780 270564
rect 209735 270524 209780 270552
rect 209774 270512 209780 270524
rect 209832 270512 209838 270564
rect 288158 270512 288164 270564
rect 288216 270552 288222 270564
rect 288345 270555 288403 270561
rect 288345 270552 288357 270555
rect 288216 270524 288357 270552
rect 288216 270512 288222 270524
rect 288345 270521 288357 270524
rect 288391 270521 288403 270555
rect 288345 270515 288403 270521
rect 153562 270484 153568 270496
rect 153523 270456 153568 270484
rect 153562 270444 153568 270456
rect 153620 270444 153626 270496
rect 257798 270484 257804 270496
rect 257759 270456 257804 270484
rect 257798 270444 257804 270456
rect 257856 270444 257862 270496
rect 304258 270444 304264 270496
rect 304316 270484 304322 270496
rect 304442 270484 304448 270496
rect 304316 270456 304448 270484
rect 304316 270444 304322 270456
rect 304442 270444 304448 270456
rect 304500 270444 304506 270496
rect 288158 270416 288164 270428
rect 288119 270388 288164 270416
rect 288158 270376 288164 270388
rect 288216 270376 288222 270428
rect 504453 269127 504511 269133
rect 504453 269093 504465 269127
rect 504499 269124 504511 269127
rect 504634 269124 504640 269136
rect 504499 269096 504640 269124
rect 504499 269093 504511 269096
rect 504453 269087 504511 269093
rect 504634 269084 504640 269096
rect 504692 269084 504698 269136
rect 132862 268404 132868 268456
rect 132920 268444 132926 268456
rect 133506 268444 133512 268456
rect 132920 268416 133512 268444
rect 132920 268404 132926 268416
rect 133506 268404 133512 268416
rect 133564 268404 133570 268456
rect 2774 264936 2780 264988
rect 2832 264976 2838 264988
rect 5442 264976 5448 264988
rect 2832 264948 5448 264976
rect 2832 264936 2838 264948
rect 5442 264936 5448 264948
rect 5500 264936 5506 264988
rect 503714 263644 503720 263696
rect 503772 263684 503778 263696
rect 503990 263684 503996 263696
rect 503772 263656 503996 263684
rect 503772 263644 503778 263656
rect 503990 263644 503996 263656
rect 504048 263644 504054 263696
rect 128906 263616 128912 263628
rect 128867 263588 128912 263616
rect 128906 263576 128912 263588
rect 128964 263576 128970 263628
rect 131574 263576 131580 263628
rect 131632 263616 131638 263628
rect 580166 263616 580172 263628
rect 131632 263588 580172 263616
rect 131632 263576 131638 263588
rect 580166 263576 580172 263588
rect 580224 263576 580230 263628
rect 257798 263548 257804 263560
rect 257759 263520 257804 263548
rect 257798 263508 257804 263520
rect 257856 263508 257862 263560
rect 503714 263508 503720 263560
rect 503772 263548 503778 263560
rect 503990 263548 503996 263560
rect 503772 263520 503996 263548
rect 503772 263508 503778 263520
rect 503990 263508 503996 263520
rect 504048 263508 504054 263560
rect 128906 260896 128912 260908
rect 128867 260868 128912 260896
rect 128906 260856 128912 260868
rect 128964 260856 128970 260908
rect 153565 260899 153623 260905
rect 153565 260865 153577 260899
rect 153611 260896 153623 260899
rect 153654 260896 153660 260908
rect 153611 260868 153660 260896
rect 153611 260865 153623 260868
rect 153565 260859 153623 260865
rect 153654 260856 153660 260868
rect 153712 260856 153718 260908
rect 288161 260899 288219 260905
rect 288161 260865 288173 260899
rect 288207 260896 288219 260899
rect 288342 260896 288348 260908
rect 288207 260868 288348 260896
rect 288207 260865 288219 260868
rect 288161 260859 288219 260865
rect 288342 260856 288348 260868
rect 288400 260856 288406 260908
rect 126057 260831 126115 260837
rect 126057 260797 126069 260831
rect 126103 260828 126115 260831
rect 126146 260828 126152 260840
rect 126103 260800 126152 260828
rect 126103 260797 126115 260800
rect 126057 260791 126115 260797
rect 126146 260788 126152 260800
rect 126204 260788 126210 260840
rect 209774 260828 209780 260840
rect 209735 260800 209780 260828
rect 209774 260788 209780 260800
rect 209832 260788 209838 260840
rect 257798 260828 257804 260840
rect 257759 260800 257804 260828
rect 257798 260788 257804 260800
rect 257856 260788 257862 260840
rect 304074 260828 304080 260840
rect 304035 260800 304080 260828
rect 304074 260788 304080 260800
rect 304132 260788 304138 260840
rect 504266 260828 504272 260840
rect 504227 260800 504272 260828
rect 504266 260788 504272 260800
rect 504324 260788 504330 260840
rect 128722 260720 128728 260772
rect 128780 260760 128786 260772
rect 128906 260760 128912 260772
rect 128780 260732 128912 260760
rect 128780 260720 128786 260732
rect 128906 260720 128912 260732
rect 128964 260720 128970 260772
rect 132862 258748 132868 258800
rect 132920 258788 132926 258800
rect 133506 258788 133512 258800
rect 132920 258760 133512 258788
rect 132920 258748 132926 258760
rect 133506 258748 133512 258760
rect 133564 258748 133570 258800
rect 153654 254028 153660 254040
rect 153580 254000 153660 254028
rect 153580 253904 153608 254000
rect 153654 253988 153660 254000
rect 153712 253988 153718 254040
rect 503622 253988 503628 254040
rect 503680 254028 503686 254040
rect 503990 254028 503996 254040
rect 503680 254000 503996 254028
rect 503680 253988 503686 254000
rect 503990 253988 503996 254000
rect 504048 253988 504054 254040
rect 153562 253852 153568 253904
rect 153620 253852 153626 253904
rect 503622 253852 503628 253904
rect 503680 253892 503686 253904
rect 503990 253892 503996 253904
rect 503680 253864 503996 253892
rect 503680 253852 503686 253864
rect 503990 253852 503996 253864
rect 504048 253852 504054 253904
rect 257798 253824 257804 253836
rect 257759 253796 257804 253824
rect 257798 253784 257804 253796
rect 257856 253784 257862 253836
rect 504266 253824 504272 253836
rect 504227 253796 504272 253824
rect 504266 253784 504272 253796
rect 504324 253784 504330 253836
rect 126054 251308 126060 251320
rect 126015 251280 126060 251308
rect 126054 251268 126060 251280
rect 126112 251268 126118 251320
rect 209774 251308 209780 251320
rect 209735 251280 209780 251308
rect 209774 251268 209780 251280
rect 209832 251268 209838 251320
rect 304077 251311 304135 251317
rect 284956 251280 288388 251308
rect 3326 251200 3332 251252
rect 3384 251240 3390 251252
rect 284956 251240 284984 251280
rect 3384 251212 284984 251240
rect 288360 251240 288388 251280
rect 304077 251277 304089 251311
rect 304123 251308 304135 251311
rect 304123 251280 304304 251308
rect 304123 251277 304135 251280
rect 304077 251271 304135 251277
rect 304276 251252 304304 251280
rect 304169 251243 304227 251249
rect 304169 251240 304181 251243
rect 288360 251212 304181 251240
rect 3384 251200 3390 251212
rect 304169 251209 304181 251212
rect 304215 251209 304227 251243
rect 304169 251203 304227 251209
rect 304258 251200 304264 251252
rect 304316 251200 304322 251252
rect 304353 251243 304411 251249
rect 304353 251209 304365 251243
rect 304399 251240 304411 251243
rect 435082 251240 435088 251252
rect 304399 251212 435088 251240
rect 304399 251209 304411 251212
rect 304353 251203 304411 251209
rect 435082 251200 435088 251212
rect 435140 251200 435146 251252
rect 257709 251175 257767 251181
rect 257709 251141 257721 251175
rect 257755 251172 257767 251175
rect 257798 251172 257804 251184
rect 257755 251144 257804 251172
rect 257755 251141 257767 251144
rect 257709 251135 257767 251141
rect 257798 251132 257804 251144
rect 257856 251132 257862 251184
rect 288250 251172 288256 251184
rect 288211 251144 288256 251172
rect 288250 251132 288256 251144
rect 288308 251132 288314 251184
rect 504266 251172 504272 251184
rect 504227 251144 504272 251172
rect 504266 251132 504272 251144
rect 504324 251132 504330 251184
rect 132862 249092 132868 249144
rect 132920 249132 132926 249144
rect 133506 249132 133512 249144
rect 132920 249104 133512 249132
rect 132920 249092 132926 249104
rect 133506 249092 133512 249104
rect 133564 249092 133570 249144
rect 503714 244400 503720 244452
rect 503772 244440 503778 244452
rect 503772 244412 503852 244440
rect 503772 244400 503778 244412
rect 503824 244384 503852 244412
rect 503806 244332 503812 244384
rect 503864 244332 503870 244384
rect 304166 244304 304172 244316
rect 304127 244276 304172 244304
rect 304166 244264 304172 244276
rect 304224 244264 304230 244316
rect 128814 244196 128820 244248
rect 128872 244236 128878 244248
rect 128998 244236 129004 244248
rect 128872 244208 129004 244236
rect 128872 244196 128878 244208
rect 128998 244196 129004 244208
rect 129056 244196 129062 244248
rect 257706 241516 257712 241528
rect 257667 241488 257712 241516
rect 257706 241476 257712 241488
rect 257764 241476 257770 241528
rect 288253 241519 288311 241525
rect 288253 241485 288265 241519
rect 288299 241516 288311 241519
rect 288342 241516 288348 241528
rect 288299 241488 288348 241516
rect 288299 241485 288311 241488
rect 288253 241479 288311 241485
rect 288342 241476 288348 241488
rect 288400 241476 288406 241528
rect 304166 241516 304172 241528
rect 304127 241488 304172 241516
rect 304166 241476 304172 241488
rect 304224 241476 304230 241528
rect 504269 241519 504327 241525
rect 504269 241485 504281 241519
rect 504315 241516 504327 241519
rect 504450 241516 504456 241528
rect 504315 241488 504456 241516
rect 504315 241485 504327 241488
rect 504269 241479 504327 241485
rect 504450 241476 504456 241488
rect 504508 241476 504514 241528
rect 304166 241380 304172 241392
rect 304127 241352 304172 241380
rect 304166 241340 304172 241352
rect 304224 241340 304230 241392
rect 132862 239436 132868 239488
rect 132920 239476 132926 239488
rect 133506 239476 133512 239488
rect 132920 239448 133512 239476
rect 132920 239436 132926 239448
rect 133506 239436 133512 239448
rect 133564 239436 133570 239488
rect 128998 236756 129004 236768
rect 128959 236728 129004 236756
rect 128998 236716 129004 236728
rect 129056 236716 129062 236768
rect 288342 236008 288348 236020
rect 288303 235980 288348 236008
rect 288342 235968 288348 235980
rect 288400 235968 288406 236020
rect 153286 234676 153292 234728
rect 153344 234676 153350 234728
rect 503622 234676 503628 234728
rect 503680 234716 503686 234728
rect 503990 234716 503996 234728
rect 503680 234688 503996 234716
rect 503680 234676 503686 234688
rect 503990 234676 503996 234688
rect 504048 234676 504054 234728
rect 504450 234716 504456 234728
rect 504376 234688 504456 234716
rect 126146 234608 126152 234660
rect 126204 234648 126210 234660
rect 126330 234648 126336 234660
rect 126204 234620 126336 234648
rect 126204 234608 126210 234620
rect 126330 234608 126336 234620
rect 126388 234608 126394 234660
rect 153304 234592 153332 234676
rect 257706 234608 257712 234660
rect 257764 234608 257770 234660
rect 153286 234540 153292 234592
rect 153344 234540 153350 234592
rect 257724 234512 257752 234608
rect 504376 234592 504404 234688
rect 504450 234676 504456 234688
rect 504508 234676 504514 234728
rect 503622 234540 503628 234592
rect 503680 234580 503686 234592
rect 503990 234580 503996 234592
rect 503680 234552 503996 234580
rect 503680 234540 503686 234552
rect 503990 234540 503996 234552
rect 504048 234540 504054 234592
rect 504358 234540 504364 234592
rect 504416 234540 504422 234592
rect 257798 234512 257804 234524
rect 257724 234484 257804 234512
rect 257798 234472 257804 234484
rect 257856 234472 257862 234524
rect 128998 231928 129004 231940
rect 128959 231900 129004 231928
rect 128998 231888 129004 231900
rect 129056 231888 129062 231940
rect 209774 231820 209780 231872
rect 209832 231860 209838 231872
rect 209958 231860 209964 231872
rect 209832 231832 209964 231860
rect 209832 231820 209838 231832
rect 209958 231820 209964 231832
rect 210016 231820 210022 231872
rect 288158 231820 288164 231872
rect 288216 231860 288222 231872
rect 288345 231863 288403 231869
rect 288345 231860 288357 231863
rect 288216 231832 288357 231860
rect 288216 231820 288222 231832
rect 288345 231829 288357 231832
rect 288391 231829 288403 231863
rect 304166 231860 304172 231872
rect 304127 231832 304172 231860
rect 288345 231823 288403 231829
rect 304166 231820 304172 231832
rect 304224 231820 304230 231872
rect 504358 231792 504364 231804
rect 504319 231764 504364 231792
rect 504358 231752 504364 231764
rect 504416 231752 504422 231804
rect 132862 229712 132868 229764
rect 132920 229752 132926 229764
rect 133506 229752 133512 229764
rect 132920 229724 133512 229752
rect 132920 229712 132926 229724
rect 133506 229712 133512 229724
rect 133564 229712 133570 229764
rect 131298 227740 131304 227792
rect 131356 227780 131362 227792
rect 580166 227780 580172 227792
rect 131356 227752 580172 227780
rect 131356 227740 131362 227752
rect 580166 227740 580172 227752
rect 580224 227740 580230 227792
rect 503714 225088 503720 225140
rect 503772 225128 503778 225140
rect 503772 225100 503852 225128
rect 503772 225088 503778 225100
rect 503824 225072 503852 225100
rect 257798 225060 257804 225072
rect 257724 225032 257804 225060
rect 153194 224992 153200 225004
rect 153155 224964 153200 224992
rect 153194 224952 153200 224964
rect 153252 224952 153258 225004
rect 257724 224936 257752 225032
rect 257798 225020 257804 225032
rect 257856 225020 257862 225072
rect 503806 225020 503812 225072
rect 503864 225020 503870 225072
rect 126146 224884 126152 224936
rect 126204 224924 126210 224936
rect 126330 224924 126336 224936
rect 126204 224896 126336 224924
rect 126204 224884 126210 224896
rect 126330 224884 126336 224896
rect 126388 224884 126394 224936
rect 257706 224884 257712 224936
rect 257764 224884 257770 224936
rect 2958 222164 2964 222216
rect 3016 222204 3022 222216
rect 14458 222204 14464 222216
rect 3016 222176 14464 222204
rect 3016 222164 3022 222176
rect 14458 222164 14464 222176
rect 14516 222164 14522 222216
rect 128630 222164 128636 222216
rect 128688 222204 128694 222216
rect 128998 222204 129004 222216
rect 128688 222176 129004 222204
rect 128688 222164 128694 222176
rect 128998 222164 129004 222176
rect 129056 222164 129062 222216
rect 153194 222204 153200 222216
rect 153155 222176 153200 222204
rect 153194 222164 153200 222176
rect 153252 222164 153258 222216
rect 288342 222164 288348 222216
rect 288400 222204 288406 222216
rect 288526 222204 288532 222216
rect 288400 222176 288532 222204
rect 288400 222164 288406 222176
rect 288526 222164 288532 222176
rect 288584 222164 288590 222216
rect 304350 222164 304356 222216
rect 304408 222204 304414 222216
rect 304534 222204 304540 222216
rect 304408 222176 304540 222204
rect 304408 222164 304414 222176
rect 304534 222164 304540 222176
rect 304592 222164 304598 222216
rect 504361 222207 504419 222213
rect 504361 222173 504373 222207
rect 504407 222204 504419 222207
rect 504450 222204 504456 222216
rect 504407 222176 504456 222204
rect 504407 222173 504419 222176
rect 504361 222167 504419 222173
rect 504450 222164 504456 222176
rect 504508 222164 504514 222216
rect 257706 222028 257712 222080
rect 257764 222068 257770 222080
rect 257982 222068 257988 222080
rect 257764 222040 257988 222068
rect 257764 222028 257770 222040
rect 257982 222028 257988 222040
rect 258040 222028 258046 222080
rect 132862 220056 132868 220108
rect 132920 220096 132926 220108
rect 133506 220096 133512 220108
rect 132920 220068 133512 220096
rect 132920 220056 132926 220068
rect 133506 220056 133512 220068
rect 133564 220056 133570 220108
rect 131482 216656 131488 216708
rect 131540 216696 131546 216708
rect 579614 216696 579620 216708
rect 131540 216668 579620 216696
rect 131540 216656 131546 216668
rect 579614 216656 579620 216668
rect 579672 216656 579678 216708
rect 503622 215364 503628 215416
rect 503680 215404 503686 215416
rect 503990 215404 503996 215416
rect 503680 215376 503996 215404
rect 503680 215364 503686 215376
rect 503990 215364 503996 215376
rect 504048 215364 504054 215416
rect 504450 215404 504456 215416
rect 504284 215376 504456 215404
rect 153194 215296 153200 215348
rect 153252 215296 153258 215348
rect 128630 215160 128636 215212
rect 128688 215200 128694 215212
rect 128998 215200 129004 215212
rect 128688 215172 129004 215200
rect 128688 215160 128694 215172
rect 128998 215160 129004 215172
rect 129056 215160 129062 215212
rect 153212 215200 153240 215296
rect 504284 215280 504312 215376
rect 504450 215364 504456 215376
rect 504508 215364 504514 215416
rect 503622 215228 503628 215280
rect 503680 215268 503686 215280
rect 503990 215268 503996 215280
rect 503680 215240 503996 215268
rect 503680 215228 503686 215240
rect 503990 215228 503996 215240
rect 504048 215228 504054 215280
rect 504266 215228 504272 215280
rect 504324 215228 504330 215280
rect 153286 215200 153292 215212
rect 153212 215172 153292 215200
rect 153286 215160 153292 215172
rect 153344 215160 153350 215212
rect 304166 213392 304172 213444
rect 304224 213432 304230 213444
rect 304350 213432 304356 213444
rect 304224 213404 304356 213432
rect 304224 213392 304230 213404
rect 304350 213392 304356 213404
rect 304408 213392 304414 213444
rect 209774 212508 209780 212560
rect 209832 212548 209838 212560
rect 209958 212548 209964 212560
rect 209832 212520 209964 212548
rect 209832 212508 209838 212520
rect 209958 212508 209964 212520
rect 210016 212508 210022 212560
rect 255314 212508 255320 212560
rect 255372 212548 255378 212560
rect 256234 212548 256240 212560
rect 255372 212520 256240 212548
rect 255372 212508 255378 212520
rect 256234 212508 256240 212520
rect 256292 212508 256298 212560
rect 288066 212508 288072 212560
rect 288124 212548 288130 212560
rect 288158 212548 288164 212560
rect 288124 212520 288164 212548
rect 288124 212508 288130 212520
rect 288158 212508 288164 212520
rect 288216 212508 288222 212560
rect 416406 212508 416412 212560
rect 416464 212548 416470 212560
rect 416682 212548 416688 212560
rect 416464 212520 416688 212548
rect 416464 212508 416470 212520
rect 416682 212508 416688 212520
rect 416740 212508 416746 212560
rect 153286 212480 153292 212492
rect 153247 212452 153292 212480
rect 153286 212440 153292 212452
rect 153344 212440 153350 212492
rect 132862 210400 132868 210452
rect 132920 210440 132926 210452
rect 133506 210440 133512 210452
rect 132920 210412 133512 210440
rect 132920 210400 132926 210412
rect 133506 210400 133512 210412
rect 133564 210400 133570 210452
rect 290918 210400 290924 210452
rect 290976 210440 290982 210452
rect 291102 210440 291108 210452
rect 290976 210412 291108 210440
rect 290976 210400 290982 210412
rect 291102 210400 291108 210412
rect 291160 210400 291166 210452
rect 243998 209720 244004 209772
rect 244056 209760 244062 209772
rect 244182 209760 244188 209772
rect 244056 209732 244188 209760
rect 244056 209720 244062 209732
rect 244182 209720 244188 209732
rect 244240 209720 244246 209772
rect 2958 207000 2964 207052
rect 3016 207040 3022 207052
rect 435174 207040 435180 207052
rect 3016 207012 435180 207040
rect 3016 207000 3022 207012
rect 435174 207000 435180 207012
rect 435232 207000 435238 207052
rect 503714 205776 503720 205828
rect 503772 205816 503778 205828
rect 503772 205788 503852 205816
rect 503772 205776 503778 205788
rect 503824 205760 503852 205788
rect 503806 205708 503812 205760
rect 503864 205708 503870 205760
rect 126422 205680 126428 205692
rect 126383 205652 126428 205680
rect 126422 205640 126428 205652
rect 126480 205640 126486 205692
rect 304074 205680 304080 205692
rect 304035 205652 304080 205680
rect 304074 205640 304080 205652
rect 304132 205640 304138 205692
rect 503714 205640 503720 205692
rect 503772 205680 503778 205692
rect 503990 205680 503996 205692
rect 503772 205652 503996 205680
rect 503772 205640 503778 205652
rect 503990 205640 503996 205652
rect 504048 205640 504054 205692
rect 504174 205680 504180 205692
rect 504135 205652 504180 205680
rect 504174 205640 504180 205652
rect 504232 205640 504238 205692
rect 126422 205544 126428 205556
rect 126383 205516 126428 205544
rect 126422 205504 126428 205516
rect 126480 205504 126486 205556
rect 196710 205300 196716 205352
rect 196768 205340 196774 205352
rect 226886 205340 226892 205352
rect 196768 205312 226892 205340
rect 196768 205300 196774 205312
rect 226886 205300 226892 205312
rect 226944 205300 226950 205352
rect 196618 205232 196624 205284
rect 196676 205272 196682 205284
rect 227898 205272 227904 205284
rect 196676 205244 227904 205272
rect 196676 205232 196682 205244
rect 227898 205232 227904 205244
rect 227956 205232 227962 205284
rect 195882 205164 195888 205216
rect 195940 205204 195946 205216
rect 228634 205204 228640 205216
rect 195940 205176 228640 205204
rect 195940 205164 195946 205176
rect 228634 205164 228640 205176
rect 228692 205164 228698 205216
rect 195698 205096 195704 205148
rect 195756 205136 195762 205148
rect 229554 205136 229560 205148
rect 195756 205108 229560 205136
rect 195756 205096 195762 205108
rect 229554 205096 229560 205108
rect 229612 205096 229618 205148
rect 195790 205028 195796 205080
rect 195848 205068 195854 205080
rect 230474 205068 230480 205080
rect 195848 205040 230480 205068
rect 195848 205028 195854 205040
rect 230474 205028 230480 205040
rect 230532 205028 230538 205080
rect 195514 204960 195520 205012
rect 195572 205000 195578 205012
rect 231210 205000 231216 205012
rect 195572 204972 231216 205000
rect 195572 204960 195578 204972
rect 231210 204960 231216 204972
rect 231268 204960 231274 205012
rect 195606 204892 195612 204944
rect 195664 204932 195670 204944
rect 233234 204932 233240 204944
rect 195664 204904 233240 204932
rect 195664 204892 195670 204904
rect 233234 204892 233240 204904
rect 233292 204892 233298 204944
rect 294414 204212 294420 204264
rect 294472 204252 294478 204264
rect 340874 204252 340880 204264
rect 294472 204224 340880 204252
rect 294472 204212 294478 204224
rect 340874 204212 340880 204224
rect 340932 204212 340938 204264
rect 345750 204212 345756 204264
rect 345808 204252 345814 204264
rect 417050 204252 417056 204264
rect 345808 204224 417056 204252
rect 345808 204212 345814 204224
rect 417050 204212 417056 204224
rect 417108 204212 417114 204264
rect 255774 204144 255780 204196
rect 255832 204184 255838 204196
rect 268194 204184 268200 204196
rect 255832 204156 268200 204184
rect 255832 204144 255838 204156
rect 268194 204144 268200 204156
rect 268252 204144 268258 204196
rect 297910 204144 297916 204196
rect 297968 204184 297974 204196
rect 304258 204184 304264 204196
rect 297968 204156 304264 204184
rect 297968 204144 297974 204156
rect 304258 204144 304264 204156
rect 304316 204144 304322 204196
rect 306650 204144 306656 204196
rect 306708 204184 306714 204196
rect 380434 204184 380440 204196
rect 306708 204156 380440 204184
rect 306708 204144 306714 204156
rect 380434 204144 380440 204156
rect 380492 204144 380498 204196
rect 253566 204076 253572 204128
rect 253624 204116 253630 204128
rect 269022 204116 269028 204128
rect 253624 204088 269028 204116
rect 253624 204076 253630 204088
rect 269022 204076 269028 204088
rect 269080 204076 269086 204128
rect 301406 204076 301412 204128
rect 301464 204116 301470 204128
rect 379606 204116 379612 204128
rect 301464 204088 379612 204116
rect 301464 204076 301470 204088
rect 379606 204076 379612 204088
rect 379664 204076 379670 204128
rect 250530 204008 250536 204060
rect 250588 204048 250594 204060
rect 267918 204048 267924 204060
rect 250588 204020 267924 204048
rect 250588 204008 250594 204020
rect 267918 204008 267924 204020
rect 267976 204008 267982 204060
rect 299014 204008 299020 204060
rect 299072 204048 299078 204060
rect 380342 204048 380348 204060
rect 299072 204020 380348 204048
rect 299072 204008 299078 204020
rect 380342 204008 380348 204020
rect 380400 204008 380406 204060
rect 199010 203940 199016 203992
rect 199068 203980 199074 203992
rect 238754 203980 238760 203992
rect 199068 203952 238760 203980
rect 199068 203940 199074 203952
rect 238754 203940 238760 203952
rect 238812 203940 238818 203992
rect 247586 203940 247592 203992
rect 247644 203980 247650 203992
rect 268102 203980 268108 203992
rect 247644 203952 268108 203980
rect 247644 203940 247650 203952
rect 268102 203940 268108 203952
rect 268160 203940 268166 203992
rect 294874 203940 294880 203992
rect 294932 203980 294938 203992
rect 377398 203980 377404 203992
rect 294932 203952 377404 203980
rect 294932 203940 294938 203952
rect 377398 203940 377404 203952
rect 377456 203940 377462 203992
rect 197722 203872 197728 203924
rect 197780 203912 197786 203924
rect 257154 203912 257160 203924
rect 197780 203884 257160 203912
rect 197780 203872 197786 203884
rect 257154 203872 257160 203884
rect 257212 203872 257218 203924
rect 292206 203872 292212 203924
rect 292264 203912 292270 203924
rect 379790 203912 379796 203924
rect 292264 203884 379796 203912
rect 292264 203872 292270 203884
rect 379790 203872 379796 203884
rect 379848 203872 379854 203924
rect 197998 203804 198004 203856
rect 198056 203844 198062 203856
rect 260374 203844 260380 203856
rect 198056 203816 260380 203844
rect 198056 203804 198062 203816
rect 260374 203804 260380 203816
rect 260432 203804 260438 203856
rect 292482 203804 292488 203856
rect 292540 203844 292546 203856
rect 379882 203844 379888 203856
rect 292540 203816 379888 203844
rect 292540 203804 292546 203816
rect 379882 203804 379888 203816
rect 379940 203804 379946 203856
rect 198458 203736 198464 203788
rect 198516 203776 198522 203788
rect 262766 203776 262772 203788
rect 198516 203748 262772 203776
rect 198516 203736 198522 203748
rect 262766 203736 262772 203748
rect 262824 203736 262830 203788
rect 286962 203736 286968 203788
rect 287020 203776 287026 203788
rect 377306 203776 377312 203788
rect 287020 203748 377312 203776
rect 287020 203736 287026 203748
rect 377306 203736 377312 203748
rect 377364 203736 377370 203788
rect 197446 203668 197452 203720
rect 197504 203708 197510 203720
rect 262950 203708 262956 203720
rect 197504 203680 262956 203708
rect 197504 203668 197510 203680
rect 262950 203668 262956 203680
rect 263008 203668 263014 203720
rect 287514 203668 287520 203720
rect 287572 203708 287578 203720
rect 379698 203708 379704 203720
rect 287572 203680 379704 203708
rect 287572 203668 287578 203680
rect 379698 203668 379704 203680
rect 379756 203668 379762 203720
rect 197814 203600 197820 203652
rect 197872 203640 197878 203652
rect 265250 203640 265256 203652
rect 197872 203612 265256 203640
rect 197872 203600 197878 203612
rect 265250 203600 265256 203612
rect 265308 203600 265314 203652
rect 271782 203600 271788 203652
rect 271840 203640 271846 203652
rect 369854 203640 369860 203652
rect 271840 203612 369860 203640
rect 271840 203600 271846 203612
rect 369854 203600 369860 203612
rect 369912 203600 369918 203652
rect 198366 203532 198372 203584
rect 198424 203572 198430 203584
rect 267550 203572 267556 203584
rect 198424 203544 267556 203572
rect 198424 203532 198430 203544
rect 267550 203532 267556 203544
rect 267608 203532 267614 203584
rect 280522 203532 280528 203584
rect 280580 203572 280586 203584
rect 379974 203572 379980 203584
rect 280580 203544 379980 203572
rect 280580 203532 280586 203544
rect 379974 203532 379980 203544
rect 380032 203532 380038 203584
rect 313550 203464 313556 203516
rect 313608 203504 313614 203516
rect 379514 203504 379520 203516
rect 313608 203476 379520 203504
rect 313608 203464 313614 203476
rect 379514 203464 379520 203476
rect 379572 203464 379578 203516
rect 296162 203396 296168 203448
rect 296220 203436 296226 203448
rect 353294 203436 353300 203448
rect 296220 203408 353300 203436
rect 296220 203396 296226 203408
rect 353294 203396 353300 203408
rect 353352 203396 353358 203448
rect 322934 203328 322940 203380
rect 322992 203368 322998 203380
rect 380158 203368 380164 203380
rect 322992 203340 380164 203368
rect 322992 203328 322998 203340
rect 380158 203328 380164 203340
rect 380216 203328 380222 203380
rect 302878 203260 302884 203312
rect 302936 203300 302942 203312
rect 331214 203300 331220 203312
rect 302936 203272 331220 203300
rect 302936 203260 302942 203272
rect 331214 203260 331220 203272
rect 331272 203260 331278 203312
rect 298002 203192 298008 203244
rect 298060 203232 298066 203244
rect 325142 203232 325148 203244
rect 298060 203204 325148 203232
rect 298060 203192 298066 203204
rect 325142 203192 325148 203204
rect 325200 203192 325206 203244
rect 128998 202960 129004 202972
rect 128924 202932 129004 202960
rect 126054 202852 126060 202904
rect 126112 202892 126118 202904
rect 126606 202892 126612 202904
rect 126112 202864 126612 202892
rect 126112 202852 126118 202864
rect 126606 202852 126612 202864
rect 126664 202852 126670 202904
rect 128924 202836 128952 202932
rect 128998 202920 129004 202932
rect 129056 202920 129062 202972
rect 153289 202895 153347 202901
rect 153289 202861 153301 202895
rect 153335 202892 153347 202895
rect 153378 202892 153384 202904
rect 153335 202864 153384 202892
rect 153335 202861 153347 202864
rect 153289 202855 153347 202861
rect 153378 202852 153384 202864
rect 153436 202852 153442 202904
rect 257706 202852 257712 202904
rect 257764 202892 257770 202904
rect 257982 202892 257988 202904
rect 257764 202864 257988 202892
rect 257764 202852 257770 202864
rect 257982 202852 257988 202864
rect 258040 202852 258046 202904
rect 304074 202892 304080 202904
rect 298848 202864 301636 202892
rect 304035 202864 304080 202892
rect 128906 202784 128912 202836
rect 128964 202784 128970 202836
rect 162118 202784 162124 202836
rect 162176 202824 162182 202836
rect 169110 202824 169116 202836
rect 162176 202796 169116 202824
rect 162176 202784 162182 202796
rect 169110 202784 169116 202796
rect 169168 202784 169174 202836
rect 199102 202784 199108 202836
rect 199160 202824 199166 202836
rect 199933 202827 199991 202833
rect 199933 202824 199945 202827
rect 199160 202796 199945 202824
rect 199160 202784 199166 202796
rect 199933 202793 199945 202796
rect 199979 202793 199991 202827
rect 199933 202787 199991 202793
rect 200022 202784 200028 202836
rect 200080 202824 200086 202836
rect 239585 202827 239643 202833
rect 239585 202824 239597 202827
rect 200080 202796 239597 202824
rect 200080 202784 200086 202796
rect 239585 202793 239597 202796
rect 239631 202793 239643 202827
rect 239585 202787 239643 202793
rect 239674 202784 239680 202836
rect 239732 202824 239738 202836
rect 240134 202824 240140 202836
rect 239732 202796 240140 202824
rect 239732 202784 239738 202796
rect 240134 202784 240140 202796
rect 240192 202784 240198 202836
rect 240502 202784 240508 202836
rect 240560 202824 240566 202836
rect 241422 202824 241428 202836
rect 240560 202796 241428 202824
rect 240560 202784 240566 202796
rect 241422 202784 241428 202796
rect 241480 202784 241486 202836
rect 242986 202784 242992 202836
rect 243044 202824 243050 202836
rect 244090 202824 244096 202836
rect 243044 202796 244096 202824
rect 243044 202784 243050 202796
rect 244090 202784 244096 202796
rect 244148 202784 244154 202836
rect 251818 202784 251824 202836
rect 251876 202824 251882 202836
rect 258813 202827 258871 202833
rect 251876 202796 258764 202824
rect 251876 202784 251882 202796
rect 196894 202716 196900 202768
rect 196952 202756 196958 202768
rect 241514 202756 241520 202768
rect 196952 202728 241520 202756
rect 196952 202716 196958 202728
rect 241514 202716 241520 202728
rect 241572 202716 241578 202768
rect 252370 202716 252376 202768
rect 252428 202756 252434 202768
rect 258629 202759 258687 202765
rect 258629 202756 258641 202759
rect 252428 202728 258641 202756
rect 252428 202716 252434 202728
rect 258629 202725 258641 202728
rect 258675 202725 258687 202759
rect 258736 202756 258764 202796
rect 258813 202793 258825 202827
rect 258859 202824 258871 202827
rect 266722 202824 266728 202836
rect 258859 202796 266728 202824
rect 258859 202793 258871 202796
rect 258813 202787 258871 202793
rect 266722 202784 266728 202796
rect 266780 202784 266786 202836
rect 272242 202784 272248 202836
rect 272300 202824 272306 202836
rect 273162 202824 273168 202836
rect 272300 202796 273168 202824
rect 272300 202784 272306 202796
rect 273162 202784 273168 202796
rect 273220 202784 273226 202836
rect 290550 202784 290556 202836
rect 290608 202824 290614 202836
rect 291010 202824 291016 202836
rect 290608 202796 291016 202824
rect 290608 202784 290614 202796
rect 291010 202784 291016 202796
rect 291068 202784 291074 202836
rect 291378 202784 291384 202836
rect 291436 202824 291442 202836
rect 292298 202824 292304 202836
rect 291436 202796 292304 202824
rect 291436 202784 291442 202796
rect 292298 202784 292304 202796
rect 292356 202784 292362 202836
rect 293126 202784 293132 202836
rect 293184 202824 293190 202836
rect 294598 202824 294604 202836
rect 293184 202796 294604 202824
rect 293184 202784 293190 202796
rect 294598 202784 294604 202796
rect 294656 202784 294662 202836
rect 295794 202784 295800 202836
rect 295852 202824 295858 202836
rect 296438 202824 296444 202836
rect 295852 202796 296444 202824
rect 295852 202784 295858 202796
rect 296438 202784 296444 202796
rect 296496 202784 296502 202836
rect 296548 202796 297864 202824
rect 267826 202756 267832 202768
rect 258736 202728 267832 202756
rect 258629 202719 258687 202725
rect 267826 202716 267832 202728
rect 267884 202716 267890 202768
rect 289262 202716 289268 202768
rect 289320 202756 289326 202768
rect 291838 202756 291844 202768
rect 289320 202728 291844 202756
rect 289320 202716 289326 202728
rect 291838 202716 291844 202728
rect 291896 202716 291902 202768
rect 199838 202648 199844 202700
rect 199896 202688 199902 202700
rect 239493 202691 239551 202697
rect 239493 202688 239505 202691
rect 199896 202660 239505 202688
rect 199896 202648 199902 202660
rect 239493 202657 239505 202660
rect 239539 202657 239551 202691
rect 239493 202651 239551 202657
rect 239585 202691 239643 202697
rect 239585 202657 239597 202691
rect 239631 202688 239643 202691
rect 245194 202688 245200 202700
rect 239631 202660 245200 202688
rect 239631 202657 239643 202660
rect 239585 202651 239643 202657
rect 245194 202648 245200 202660
rect 245252 202648 245258 202700
rect 247494 202648 247500 202700
rect 247552 202688 247558 202700
rect 253845 202691 253903 202697
rect 253845 202688 253857 202691
rect 247552 202660 253857 202688
rect 247552 202648 247558 202660
rect 253845 202657 253857 202660
rect 253891 202657 253903 202691
rect 266630 202688 266636 202700
rect 253845 202651 253903 202657
rect 255240 202660 266636 202688
rect 197630 202580 197636 202632
rect 197688 202620 197694 202632
rect 244734 202620 244740 202632
rect 197688 202592 244740 202620
rect 197688 202580 197694 202592
rect 244734 202580 244740 202592
rect 244792 202580 244798 202632
rect 250898 202580 250904 202632
rect 250956 202620 250962 202632
rect 255240 202620 255268 202660
rect 266630 202648 266636 202660
rect 266688 202648 266694 202700
rect 250956 202592 255268 202620
rect 255593 202623 255651 202629
rect 250956 202580 250962 202592
rect 255593 202589 255605 202623
rect 255639 202620 255651 202623
rect 268286 202620 268292 202632
rect 255639 202592 268292 202620
rect 255639 202589 255651 202592
rect 255593 202583 255651 202589
rect 268286 202580 268292 202592
rect 268344 202580 268350 202632
rect 288802 202580 288808 202632
rect 288860 202620 288866 202632
rect 296548 202620 296576 202796
rect 297836 202756 297864 202796
rect 297910 202784 297916 202836
rect 297968 202824 297974 202836
rect 298738 202824 298744 202836
rect 297968 202796 298744 202824
rect 297968 202784 297974 202796
rect 298738 202784 298744 202796
rect 298796 202784 298802 202836
rect 298848 202756 298876 202864
rect 298922 202784 298928 202836
rect 298980 202824 298986 202836
rect 301498 202824 301504 202836
rect 298980 202796 301504 202824
rect 298980 202784 298986 202796
rect 301498 202784 301504 202796
rect 301556 202784 301562 202836
rect 301608 202824 301636 202864
rect 304074 202852 304080 202864
rect 304132 202852 304138 202904
rect 504174 202892 504180 202904
rect 504135 202864 504180 202892
rect 504174 202852 504180 202864
rect 504232 202852 504238 202904
rect 305638 202824 305644 202836
rect 301608 202796 305644 202824
rect 305638 202784 305644 202796
rect 305696 202784 305702 202836
rect 309134 202784 309140 202836
rect 309192 202824 309198 202836
rect 309594 202824 309600 202836
rect 309192 202796 309600 202824
rect 309192 202784 309198 202796
rect 309594 202784 309600 202796
rect 309652 202784 309658 202836
rect 311894 202784 311900 202836
rect 311952 202824 311958 202836
rect 312538 202824 312544 202836
rect 311952 202796 312544 202824
rect 311952 202784 311958 202796
rect 312538 202784 312544 202796
rect 312596 202784 312602 202836
rect 314838 202784 314844 202836
rect 314896 202824 314902 202836
rect 315574 202824 315580 202836
rect 314896 202796 315580 202824
rect 314896 202784 314902 202796
rect 315574 202784 315580 202796
rect 315632 202784 315638 202836
rect 315669 202827 315727 202833
rect 315669 202793 315681 202827
rect 315715 202824 315727 202827
rect 375561 202827 375619 202833
rect 375561 202824 375573 202827
rect 315715 202796 375573 202824
rect 315715 202793 315727 202796
rect 315669 202787 315727 202793
rect 375561 202793 375573 202796
rect 375607 202793 375619 202827
rect 375561 202787 375619 202793
rect 375742 202784 375748 202836
rect 375800 202824 375806 202836
rect 378778 202824 378784 202836
rect 375800 202796 378784 202824
rect 375800 202784 375806 202796
rect 378778 202784 378784 202796
rect 378836 202784 378842 202836
rect 400582 202784 400588 202836
rect 400640 202824 400646 202836
rect 401502 202824 401508 202836
rect 400640 202796 401508 202824
rect 400640 202784 400646 202796
rect 401502 202784 401508 202796
rect 401560 202784 401566 202836
rect 297836 202728 298876 202756
rect 299106 202716 299112 202768
rect 299164 202756 299170 202768
rect 302421 202759 302479 202765
rect 299164 202728 302372 202756
rect 299164 202716 299170 202728
rect 299198 202648 299204 202700
rect 299256 202688 299262 202700
rect 302237 202691 302295 202697
rect 302237 202688 302249 202691
rect 299256 202660 302249 202688
rect 299256 202648 299262 202660
rect 302237 202657 302249 202660
rect 302283 202657 302295 202691
rect 302344 202688 302372 202728
rect 302421 202725 302433 202759
rect 302467 202756 302479 202759
rect 318337 202759 318395 202765
rect 318337 202756 318349 202759
rect 302467 202728 318349 202756
rect 302467 202725 302479 202728
rect 302421 202719 302479 202725
rect 318337 202725 318349 202728
rect 318383 202725 318395 202759
rect 318337 202719 318395 202725
rect 319254 202716 319260 202768
rect 319312 202756 319318 202768
rect 320082 202756 320088 202768
rect 319312 202728 320088 202756
rect 319312 202716 319318 202728
rect 320082 202716 320088 202728
rect 320140 202716 320146 202768
rect 320542 202716 320548 202768
rect 320600 202756 320606 202768
rect 321462 202756 321468 202768
rect 320600 202728 321468 202756
rect 320600 202716 320606 202728
rect 321462 202716 321468 202728
rect 321520 202716 321526 202768
rect 333146 202716 333152 202768
rect 333204 202756 333210 202768
rect 333882 202756 333888 202768
rect 333204 202728 333888 202756
rect 333204 202716 333210 202728
rect 333882 202716 333888 202728
rect 333940 202716 333946 202768
rect 342070 202716 342076 202768
rect 342128 202756 342134 202768
rect 347685 202759 347743 202765
rect 347685 202756 347697 202759
rect 342128 202728 347697 202756
rect 342128 202716 342134 202728
rect 347685 202725 347697 202728
rect 347731 202725 347743 202759
rect 347685 202719 347743 202725
rect 349982 202716 349988 202768
rect 350040 202756 350046 202768
rect 350442 202756 350448 202768
rect 350040 202728 350448 202756
rect 350040 202716 350046 202728
rect 350442 202716 350448 202728
rect 350500 202716 350506 202768
rect 350994 202716 351000 202768
rect 351052 202756 351058 202768
rect 351822 202756 351828 202768
rect 351052 202728 351828 202756
rect 351052 202716 351058 202728
rect 351822 202716 351828 202728
rect 351880 202716 351886 202768
rect 351917 202759 351975 202765
rect 351917 202725 351929 202759
rect 351963 202756 351975 202759
rect 417142 202756 417148 202768
rect 351963 202728 417148 202756
rect 351963 202725 351975 202728
rect 351917 202719 351975 202725
rect 417142 202716 417148 202728
rect 417200 202716 417206 202768
rect 302970 202688 302976 202700
rect 302344 202660 302976 202688
rect 302237 202651 302295 202657
rect 302970 202648 302976 202660
rect 303028 202648 303034 202700
rect 325694 202688 325700 202700
rect 304368 202660 325700 202688
rect 288860 202592 296576 202620
rect 288860 202580 288866 202592
rect 299658 202580 299664 202632
rect 299716 202620 299722 202632
rect 304368 202620 304396 202660
rect 325694 202648 325700 202660
rect 325752 202648 325758 202700
rect 344002 202648 344008 202700
rect 344060 202688 344066 202700
rect 416866 202688 416872 202700
rect 344060 202660 416872 202688
rect 344060 202648 344066 202660
rect 416866 202648 416872 202660
rect 416924 202648 416930 202700
rect 299716 202592 304396 202620
rect 304905 202623 304963 202629
rect 299716 202580 299722 202592
rect 304905 202589 304917 202623
rect 304951 202620 304963 202623
rect 338758 202620 338764 202632
rect 304951 202592 338764 202620
rect 304951 202589 304963 202592
rect 304905 202583 304963 202589
rect 338758 202580 338764 202592
rect 338816 202580 338822 202632
rect 341426 202580 341432 202632
rect 341484 202620 341490 202632
rect 342162 202620 342168 202632
rect 341484 202592 342168 202620
rect 341484 202580 341490 202592
rect 342162 202580 342168 202592
rect 342220 202580 342226 202632
rect 343082 202580 343088 202632
rect 343140 202620 343146 202632
rect 343542 202620 343548 202632
rect 343140 202592 343548 202620
rect 343140 202580 343146 202592
rect 343542 202580 343548 202592
rect 343600 202580 343606 202632
rect 346670 202580 346676 202632
rect 346728 202620 346734 202632
rect 347590 202620 347596 202632
rect 346728 202592 347596 202620
rect 346728 202580 346734 202592
rect 347590 202580 347596 202592
rect 347648 202580 347654 202632
rect 347685 202623 347743 202629
rect 347685 202589 347697 202623
rect 347731 202620 347743 202623
rect 415394 202620 415400 202632
rect 347731 202592 415400 202620
rect 347731 202589 347743 202592
rect 347685 202583 347743 202589
rect 415394 202580 415400 202592
rect 415452 202580 415458 202632
rect 159358 202512 159364 202564
rect 159416 202552 159422 202564
rect 176930 202552 176936 202564
rect 159416 202524 176936 202552
rect 159416 202512 159422 202524
rect 176930 202512 176936 202524
rect 176988 202512 176994 202564
rect 197538 202512 197544 202564
rect 197596 202552 197602 202564
rect 245654 202552 245660 202564
rect 197596 202524 245660 202552
rect 197596 202512 197602 202524
rect 245654 202512 245660 202524
rect 245712 202512 245718 202564
rect 248785 202555 248843 202561
rect 248785 202521 248797 202555
rect 248831 202552 248843 202555
rect 253845 202555 253903 202561
rect 248831 202524 253796 202552
rect 248831 202521 248843 202524
rect 248785 202515 248843 202521
rect 160738 202444 160744 202496
rect 160796 202484 160802 202496
rect 178034 202484 178040 202496
rect 160796 202456 178040 202484
rect 160796 202444 160802 202456
rect 178034 202444 178040 202456
rect 178092 202444 178098 202496
rect 197354 202444 197360 202496
rect 197412 202484 197418 202496
rect 244829 202487 244887 202493
rect 244829 202484 244841 202487
rect 197412 202456 244841 202484
rect 197412 202444 197418 202456
rect 244829 202453 244841 202456
rect 244875 202453 244887 202487
rect 244829 202447 244887 202453
rect 244918 202444 244924 202496
rect 244976 202484 244982 202496
rect 246022 202484 246028 202496
rect 244976 202456 246028 202484
rect 244976 202444 244982 202456
rect 246022 202444 246028 202456
rect 246080 202444 246086 202496
rect 250070 202444 250076 202496
rect 250128 202484 250134 202496
rect 250990 202484 250996 202496
rect 250128 202456 250996 202484
rect 250128 202444 250134 202456
rect 250990 202444 250996 202456
rect 251048 202444 251054 202496
rect 253768 202484 253796 202524
rect 253845 202521 253857 202555
rect 253891 202552 253903 202555
rect 267734 202552 267740 202564
rect 253891 202524 258028 202552
rect 253891 202521 253903 202524
rect 253845 202515 253903 202521
rect 258000 202484 258028 202524
rect 258184 202524 267740 202552
rect 258184 202484 258212 202524
rect 267734 202512 267740 202524
rect 267792 202512 267798 202564
rect 271414 202512 271420 202564
rect 271472 202552 271478 202564
rect 272518 202552 272524 202564
rect 271472 202524 272524 202552
rect 271472 202512 271478 202524
rect 272518 202512 272524 202524
rect 272576 202512 272582 202564
rect 299382 202512 299388 202564
rect 299440 202552 299446 202564
rect 302421 202555 302479 202561
rect 302421 202552 302433 202555
rect 299440 202524 302433 202552
rect 299440 202512 299446 202524
rect 302421 202521 302433 202524
rect 302467 202521 302479 202555
rect 302421 202515 302479 202521
rect 302881 202555 302939 202561
rect 302881 202521 302893 202555
rect 302927 202552 302939 202555
rect 375469 202555 375527 202561
rect 375469 202552 375481 202555
rect 302927 202524 375481 202552
rect 302927 202521 302939 202524
rect 302881 202515 302939 202521
rect 375469 202521 375481 202524
rect 375515 202521 375527 202555
rect 375469 202515 375527 202521
rect 375561 202555 375619 202561
rect 375561 202521 375573 202555
rect 375607 202552 375619 202555
rect 377214 202552 377220 202564
rect 375607 202524 377220 202552
rect 375607 202521 375619 202524
rect 375561 202515 375619 202521
rect 377214 202512 377220 202524
rect 377272 202512 377278 202564
rect 400950 202512 400956 202564
rect 401008 202552 401014 202564
rect 414658 202552 414664 202564
rect 401008 202524 414664 202552
rect 401008 202512 401014 202524
rect 414658 202512 414664 202524
rect 414716 202512 414722 202564
rect 253768 202456 257108 202484
rect 258000 202456 258212 202484
rect 258629 202487 258687 202493
rect 157978 202376 157984 202428
rect 158036 202416 158042 202428
rect 182174 202416 182180 202428
rect 158036 202388 182180 202416
rect 158036 202376 158042 202388
rect 182174 202376 182180 202388
rect 182232 202376 182238 202428
rect 199194 202376 199200 202428
rect 199252 202416 199258 202428
rect 254026 202416 254032 202428
rect 199252 202388 254032 202416
rect 199252 202376 199258 202388
rect 254026 202376 254032 202388
rect 254084 202376 254090 202428
rect 153838 202308 153844 202360
rect 153896 202348 153902 202360
rect 181254 202348 181260 202360
rect 153896 202320 181260 202348
rect 153896 202308 153902 202320
rect 181254 202308 181260 202320
rect 181312 202308 181318 202360
rect 200025 202351 200083 202357
rect 200025 202317 200037 202351
rect 200071 202348 200083 202351
rect 211801 202351 211859 202357
rect 211801 202348 211813 202351
rect 200071 202320 211813 202348
rect 200071 202317 200083 202320
rect 200025 202311 200083 202317
rect 211801 202317 211813 202320
rect 211847 202317 211859 202351
rect 211801 202311 211859 202317
rect 219345 202351 219403 202357
rect 219345 202317 219357 202351
rect 219391 202348 219403 202351
rect 229097 202351 229155 202357
rect 229097 202348 229109 202351
rect 219391 202320 229109 202348
rect 219391 202317 219403 202320
rect 219345 202311 219403 202317
rect 229097 202317 229109 202320
rect 229143 202317 229155 202351
rect 229097 202311 229155 202317
rect 238665 202351 238723 202357
rect 238665 202317 238677 202351
rect 238711 202348 238723 202351
rect 238711 202320 248920 202348
rect 238711 202317 238723 202320
rect 238665 202311 238723 202317
rect 140038 202240 140044 202292
rect 140096 202280 140102 202292
rect 168374 202280 168380 202292
rect 140096 202252 168380 202280
rect 140096 202240 140102 202252
rect 168374 202240 168380 202252
rect 168432 202240 168438 202292
rect 199933 202283 199991 202289
rect 199933 202249 199945 202283
rect 199979 202280 199991 202283
rect 215205 202283 215263 202289
rect 215205 202280 215217 202283
rect 199979 202252 215217 202280
rect 199979 202249 199991 202252
rect 199933 202243 199991 202249
rect 215205 202249 215217 202252
rect 215251 202249 215263 202283
rect 215205 202243 215263 202249
rect 219253 202283 219311 202289
rect 219253 202249 219265 202283
rect 219299 202280 219311 202283
rect 229189 202283 229247 202289
rect 229189 202280 229201 202283
rect 219299 202252 229201 202280
rect 219299 202249 219311 202252
rect 219253 202243 219311 202249
rect 229189 202249 229201 202252
rect 229235 202249 229247 202283
rect 229189 202243 229247 202249
rect 238573 202283 238631 202289
rect 238573 202249 238585 202283
rect 238619 202280 238631 202283
rect 248785 202283 248843 202289
rect 248785 202280 248797 202283
rect 238619 202252 248797 202280
rect 238619 202249 238631 202252
rect 238573 202243 238631 202249
rect 248785 202249 248797 202252
rect 248831 202249 248843 202283
rect 248892 202280 248920 202320
rect 248966 202308 248972 202360
rect 249024 202348 249030 202360
rect 255593 202351 255651 202357
rect 255593 202348 255605 202351
rect 249024 202320 255605 202348
rect 249024 202308 249030 202320
rect 255593 202317 255605 202320
rect 255639 202317 255651 202351
rect 257080 202348 257108 202456
rect 258629 202453 258641 202487
rect 258675 202484 258687 202487
rect 268378 202484 268384 202496
rect 258675 202456 268384 202484
rect 258675 202453 258687 202456
rect 258629 202447 258687 202453
rect 268378 202444 268384 202456
rect 268436 202444 268442 202496
rect 273990 202444 273996 202496
rect 274048 202484 274054 202496
rect 274542 202484 274548 202496
rect 274048 202456 274548 202484
rect 274048 202444 274054 202456
rect 274542 202444 274548 202456
rect 274600 202444 274606 202496
rect 276934 202444 276940 202496
rect 276992 202484 276998 202496
rect 277302 202484 277308 202496
rect 276992 202456 277308 202484
rect 276992 202444 276998 202456
rect 277302 202444 277308 202456
rect 277360 202444 277366 202496
rect 278682 202444 278688 202496
rect 278740 202484 278746 202496
rect 279418 202484 279424 202496
rect 278740 202456 279424 202484
rect 278740 202444 278746 202456
rect 279418 202444 279424 202456
rect 279476 202444 279482 202496
rect 280982 202444 280988 202496
rect 281040 202484 281046 202496
rect 281350 202484 281356 202496
rect 281040 202456 281356 202484
rect 281040 202444 281046 202456
rect 281350 202444 281356 202456
rect 281408 202444 281414 202496
rect 297726 202444 297732 202496
rect 297784 202484 297790 202496
rect 303890 202484 303896 202496
rect 297784 202456 303896 202484
rect 297784 202444 297790 202456
rect 303890 202444 303896 202456
rect 303948 202444 303954 202496
rect 304902 202444 304908 202496
rect 304960 202484 304966 202496
rect 309134 202484 309140 202496
rect 304960 202456 309140 202484
rect 304960 202444 304966 202456
rect 309134 202444 309140 202456
rect 309192 202444 309198 202496
rect 310606 202444 310612 202496
rect 310664 202484 310670 202496
rect 311250 202484 311256 202496
rect 310664 202456 311256 202484
rect 310664 202444 310670 202456
rect 311250 202444 311256 202456
rect 311308 202444 311314 202496
rect 311345 202487 311403 202493
rect 311345 202453 311357 202487
rect 311391 202484 311403 202487
rect 377490 202484 377496 202496
rect 311391 202456 377496 202484
rect 311391 202453 311403 202456
rect 311345 202447 311403 202453
rect 377490 202444 377496 202456
rect 377548 202444 377554 202496
rect 413186 202444 413192 202496
rect 413244 202484 413250 202496
rect 416038 202484 416044 202496
rect 413244 202456 416044 202484
rect 413244 202444 413250 202456
rect 416038 202444 416044 202456
rect 416096 202444 416102 202496
rect 416133 202487 416191 202493
rect 416133 202453 416145 202487
rect 416179 202484 416191 202487
rect 457438 202484 457444 202496
rect 416179 202456 457444 202484
rect 416179 202453 416191 202456
rect 416133 202447 416191 202453
rect 457438 202444 457444 202456
rect 457496 202444 457502 202496
rect 260190 202416 260196 202428
rect 258184 202388 260196 202416
rect 258184 202348 258212 202388
rect 260190 202376 260196 202388
rect 260248 202376 260254 202428
rect 268470 202416 268476 202428
rect 260300 202388 268476 202416
rect 257080 202320 258212 202348
rect 258353 202351 258411 202357
rect 255593 202311 255651 202317
rect 258353 202317 258365 202351
rect 258399 202348 258411 202351
rect 260300 202348 260328 202388
rect 268470 202376 268476 202388
rect 268528 202376 268534 202428
rect 275278 202376 275284 202428
rect 275336 202416 275342 202428
rect 286410 202416 286416 202428
rect 275336 202388 286416 202416
rect 275336 202376 275342 202388
rect 286410 202376 286416 202388
rect 286468 202376 286474 202428
rect 301866 202376 301872 202428
rect 301924 202416 301930 202428
rect 302881 202419 302939 202425
rect 302881 202416 302893 202419
rect 301924 202388 302893 202416
rect 301924 202376 301930 202388
rect 302881 202385 302893 202388
rect 302927 202385 302939 202419
rect 302881 202379 302939 202385
rect 302973 202419 303031 202425
rect 302973 202385 302985 202419
rect 303019 202416 303031 202419
rect 304074 202416 304080 202428
rect 303019 202388 304080 202416
rect 303019 202385 303031 202388
rect 302973 202379 303031 202385
rect 304074 202376 304080 202388
rect 304132 202376 304138 202428
rect 307018 202376 307024 202428
rect 307076 202416 307082 202428
rect 308398 202416 308404 202428
rect 307076 202388 308404 202416
rect 307076 202376 307082 202388
rect 308398 202376 308404 202388
rect 308456 202376 308462 202428
rect 308493 202419 308551 202425
rect 308493 202385 308505 202419
rect 308539 202416 308551 202419
rect 322934 202416 322940 202428
rect 308539 202388 322940 202416
rect 308539 202385 308551 202388
rect 308493 202379 308551 202385
rect 322934 202376 322940 202388
rect 322992 202376 322998 202428
rect 332502 202376 332508 202428
rect 332560 202416 332566 202428
rect 332560 202388 412220 202416
rect 332560 202376 332566 202388
rect 258399 202320 260328 202348
rect 258399 202317 258411 202320
rect 258353 202311 258411 202317
rect 261662 202308 261668 202360
rect 261720 202348 261726 202360
rect 262122 202348 262128 202360
rect 261720 202320 262128 202348
rect 261720 202308 261726 202320
rect 262122 202308 262128 202320
rect 262180 202308 262186 202360
rect 262217 202351 262275 202357
rect 262217 202317 262229 202351
rect 262263 202348 262275 202351
rect 266814 202348 266820 202360
rect 262263 202320 266820 202348
rect 262263 202317 262275 202320
rect 262217 202311 262275 202317
rect 266814 202308 266820 202320
rect 266872 202308 266878 202360
rect 275738 202308 275744 202360
rect 275796 202348 275802 202360
rect 286318 202348 286324 202360
rect 275796 202320 286324 202348
rect 275796 202308 275802 202320
rect 286318 202308 286324 202320
rect 286376 202308 286382 202360
rect 300118 202308 300124 202360
rect 300176 202348 300182 202360
rect 374365 202351 374423 202357
rect 374365 202348 374377 202351
rect 300176 202320 374377 202348
rect 300176 202308 300182 202320
rect 374365 202317 374377 202320
rect 374411 202317 374423 202351
rect 374365 202311 374423 202317
rect 374454 202308 374460 202360
rect 374512 202348 374518 202360
rect 375282 202348 375288 202360
rect 374512 202320 375288 202348
rect 374512 202308 374518 202320
rect 375282 202308 375288 202320
rect 375340 202308 375346 202360
rect 375469 202351 375527 202357
rect 375469 202317 375481 202351
rect 375515 202348 375527 202351
rect 378962 202348 378968 202360
rect 375515 202320 378968 202348
rect 375515 202317 375527 202320
rect 375469 202311 375527 202317
rect 378962 202308 378968 202320
rect 379020 202308 379026 202360
rect 412192 202348 412220 202388
rect 415762 202376 415768 202428
rect 415820 202416 415826 202428
rect 416590 202416 416596 202428
rect 415820 202388 416596 202416
rect 415820 202376 415826 202388
rect 416590 202376 416596 202388
rect 416648 202376 416654 202428
rect 417510 202376 417516 202428
rect 417568 202416 417574 202428
rect 418062 202416 418068 202428
rect 417568 202388 418068 202416
rect 417568 202376 417574 202388
rect 418062 202376 418068 202388
rect 418120 202376 418126 202428
rect 416774 202348 416780 202360
rect 412192 202320 416780 202348
rect 416774 202308 416780 202320
rect 416832 202308 416838 202360
rect 503898 202348 503904 202360
rect 416884 202320 503904 202348
rect 258166 202280 258172 202292
rect 248892 202252 258172 202280
rect 248785 202243 248843 202249
rect 258166 202240 258172 202252
rect 258224 202240 258230 202292
rect 258261 202283 258319 202289
rect 258261 202249 258273 202283
rect 258307 202280 258319 202283
rect 261938 202280 261944 202292
rect 258307 202252 261944 202280
rect 258307 202249 258319 202252
rect 258261 202243 258319 202249
rect 261938 202240 261944 202252
rect 261996 202240 262002 202292
rect 277302 202240 277308 202292
rect 277360 202280 277366 202292
rect 378134 202280 378140 202292
rect 277360 202252 378140 202280
rect 277360 202240 277366 202252
rect 378134 202240 378140 202252
rect 378192 202240 378198 202292
rect 414934 202240 414940 202292
rect 414992 202280 414998 202292
rect 416884 202280 416912 202320
rect 503898 202308 503904 202320
rect 503956 202308 503962 202360
rect 503806 202280 503812 202292
rect 414992 202252 416912 202280
rect 416976 202252 503812 202280
rect 414992 202240 414998 202252
rect 103422 202172 103428 202224
rect 103480 202212 103486 202224
rect 142522 202212 142528 202224
rect 103480 202184 142528 202212
rect 103480 202172 103486 202184
rect 142522 202172 142528 202184
rect 142580 202172 142586 202224
rect 151078 202172 151084 202224
rect 151136 202212 151142 202224
rect 180334 202212 180340 202224
rect 151136 202184 180340 202212
rect 151136 202172 151142 202184
rect 180334 202172 180340 202184
rect 180392 202172 180398 202224
rect 198826 202172 198832 202224
rect 198884 202212 198890 202224
rect 257985 202215 258043 202221
rect 257985 202212 257997 202215
rect 198884 202184 257997 202212
rect 198884 202172 198890 202184
rect 257985 202181 257997 202184
rect 258031 202181 258043 202215
rect 257985 202175 258043 202181
rect 264057 202215 264115 202221
rect 264057 202181 264069 202215
rect 264103 202212 264115 202215
rect 268562 202212 268568 202224
rect 264103 202184 268568 202212
rect 264103 202181 264115 202184
rect 264057 202175 264115 202181
rect 268562 202172 268568 202184
rect 268620 202172 268626 202224
rect 270954 202172 270960 202224
rect 271012 202212 271018 202224
rect 374273 202215 374331 202221
rect 374273 202212 374285 202215
rect 271012 202184 374285 202212
rect 271012 202172 271018 202184
rect 374273 202181 374285 202184
rect 374319 202181 374331 202215
rect 374273 202175 374331 202181
rect 374365 202215 374423 202221
rect 374365 202181 374377 202215
rect 374411 202212 374423 202215
rect 378318 202212 378324 202224
rect 374411 202184 378324 202212
rect 374411 202181 374423 202184
rect 374365 202175 374423 202181
rect 378318 202172 378324 202184
rect 378376 202172 378382 202224
rect 411070 202172 411076 202224
rect 411128 202212 411134 202224
rect 416976 202212 417004 202252
rect 503806 202240 503812 202252
rect 503864 202240 503870 202292
rect 411128 202184 417004 202212
rect 417053 202215 417111 202221
rect 411128 202172 411134 202184
rect 417053 202181 417065 202215
rect 417099 202212 417111 202215
rect 503714 202212 503720 202224
rect 417099 202184 503720 202212
rect 417099 202181 417111 202184
rect 417053 202175 417111 202181
rect 503714 202172 503720 202184
rect 503772 202172 503778 202224
rect 93762 202104 93768 202156
rect 93820 202144 93826 202156
rect 134702 202144 134708 202156
rect 93820 202116 134708 202144
rect 93820 202104 93826 202116
rect 134702 202104 134708 202116
rect 134760 202104 134766 202156
rect 146938 202104 146944 202156
rect 146996 202144 147002 202156
rect 178678 202144 178684 202156
rect 146996 202116 178684 202144
rect 146996 202104 147002 202116
rect 178678 202104 178684 202116
rect 178736 202104 178742 202156
rect 197906 202104 197912 202156
rect 197964 202144 197970 202156
rect 269482 202144 269488 202156
rect 197964 202116 269488 202144
rect 197964 202104 197970 202116
rect 269482 202104 269488 202116
rect 269540 202104 269546 202156
rect 283558 202104 283564 202156
rect 283616 202144 283622 202156
rect 340138 202144 340144 202156
rect 283616 202116 340144 202144
rect 283616 202104 283622 202116
rect 340138 202104 340144 202116
rect 340196 202104 340202 202156
rect 348326 202104 348332 202156
rect 348384 202144 348390 202156
rect 351917 202147 351975 202153
rect 351917 202144 351929 202147
rect 348384 202116 351929 202144
rect 348384 202104 348390 202116
rect 351917 202113 351929 202116
rect 351963 202113 351975 202147
rect 351917 202107 351975 202113
rect 353570 202104 353576 202156
rect 353628 202144 353634 202156
rect 354582 202144 354588 202156
rect 353628 202116 354588 202144
rect 353628 202104 353634 202116
rect 354582 202104 354588 202116
rect 354640 202104 354646 202156
rect 366174 202104 366180 202156
rect 366232 202144 366238 202156
rect 367002 202144 367008 202156
rect 366232 202116 367008 202144
rect 366232 202104 366238 202116
rect 367002 202104 367008 202116
rect 367060 202104 367066 202156
rect 376478 202104 376484 202156
rect 376536 202144 376542 202156
rect 506474 202144 506480 202156
rect 376536 202116 506480 202144
rect 376536 202104 376542 202116
rect 506474 202104 506480 202116
rect 506532 202104 506538 202156
rect 198918 202036 198924 202088
rect 198976 202076 198982 202088
rect 199841 202079 199899 202085
rect 199841 202076 199853 202079
rect 198976 202048 199853 202076
rect 198976 202036 198982 202048
rect 199841 202045 199853 202048
rect 199887 202045 199899 202079
rect 199841 202039 199899 202045
rect 199930 202036 199936 202088
rect 199988 202076 199994 202088
rect 229094 202076 229100 202088
rect 199988 202048 229100 202076
rect 199988 202036 199994 202048
rect 229094 202036 229100 202048
rect 229152 202036 229158 202088
rect 240962 202036 240968 202088
rect 241020 202076 241026 202088
rect 267366 202076 267372 202088
rect 241020 202048 267372 202076
rect 241020 202036 241026 202048
rect 267366 202036 267372 202048
rect 267424 202036 267430 202088
rect 289538 202036 289544 202088
rect 289596 202076 289602 202088
rect 302973 202079 303031 202085
rect 302973 202076 302985 202079
rect 289596 202048 302985 202076
rect 289596 202036 289602 202048
rect 302973 202045 302985 202048
rect 303019 202045 303031 202079
rect 311345 202079 311403 202085
rect 311345 202076 311357 202079
rect 302973 202039 303031 202045
rect 303080 202048 311357 202076
rect 199746 201968 199752 202020
rect 199804 202008 199810 202020
rect 233605 202011 233663 202017
rect 233605 202008 233617 202011
rect 199804 201980 233617 202008
rect 199804 201968 199810 201980
rect 233605 201977 233617 201980
rect 233651 201977 233663 202011
rect 233605 201971 233663 201977
rect 233697 202011 233755 202017
rect 233697 201977 233709 202011
rect 233743 202008 233755 202011
rect 236549 202011 236607 202017
rect 236549 202008 236561 202011
rect 233743 201980 236561 202008
rect 233743 201977 233755 201980
rect 233697 201971 233755 201977
rect 236549 201977 236561 201980
rect 236595 201977 236607 202011
rect 236549 201971 236607 201977
rect 236638 201968 236644 202020
rect 236696 202008 236702 202020
rect 237282 202008 237288 202020
rect 236696 201980 237288 202008
rect 236696 201968 236702 201980
rect 237282 201968 237288 201980
rect 237340 201968 237346 202020
rect 237377 202011 237435 202017
rect 237377 201977 237389 202011
rect 237423 202008 237435 202011
rect 238573 202011 238631 202017
rect 238573 202008 238585 202011
rect 237423 201980 238585 202008
rect 237423 201977 237435 201980
rect 237377 201971 237435 201977
rect 238573 201977 238585 201980
rect 238619 201977 238631 202011
rect 238573 201971 238631 201977
rect 238662 201968 238668 202020
rect 238720 202008 238726 202020
rect 241054 202008 241060 202020
rect 238720 201980 241060 202008
rect 238720 201968 238726 201980
rect 241054 201968 241060 201980
rect 241112 201968 241118 202020
rect 244642 201968 244648 202020
rect 244700 202008 244706 202020
rect 268010 202008 268016 202020
rect 244700 201980 268016 202008
rect 244700 201968 244706 201980
rect 268010 201968 268016 201980
rect 268068 201968 268074 202020
rect 300762 201968 300768 202020
rect 300820 202008 300826 202020
rect 303080 202008 303108 202048
rect 311345 202045 311357 202048
rect 311391 202045 311403 202079
rect 311345 202039 311403 202045
rect 315298 202036 315304 202088
rect 315356 202076 315362 202088
rect 315942 202076 315948 202088
rect 315356 202048 315948 202076
rect 315356 202036 315362 202048
rect 315942 202036 315948 202048
rect 316000 202036 316006 202088
rect 316034 202036 316040 202088
rect 316092 202076 316098 202088
rect 317138 202076 317144 202088
rect 316092 202048 317144 202076
rect 316092 202036 316098 202048
rect 317138 202036 317144 202048
rect 317196 202036 317202 202088
rect 318610 202036 318616 202088
rect 318668 202076 318674 202088
rect 337378 202076 337384 202088
rect 318668 202048 337384 202076
rect 318668 202036 318674 202048
rect 337378 202036 337384 202048
rect 337436 202036 337442 202088
rect 352742 202036 352748 202088
rect 352800 202076 352806 202088
rect 353202 202076 353208 202088
rect 352800 202048 353208 202076
rect 352800 202036 352806 202048
rect 353202 202036 353208 202048
rect 353260 202036 353266 202088
rect 417234 202076 417240 202088
rect 353312 202048 417240 202076
rect 305638 202008 305644 202020
rect 300820 201980 303108 202008
rect 303632 201980 305644 202008
rect 300820 201968 300826 201980
rect 198642 201900 198648 201952
rect 198700 201940 198706 201952
rect 216030 201940 216036 201952
rect 198700 201912 216036 201940
rect 198700 201900 198706 201912
rect 216030 201900 216036 201912
rect 216088 201900 216094 201952
rect 239125 201943 239183 201949
rect 239125 201940 239137 201943
rect 216140 201912 239137 201940
rect 198734 201832 198740 201884
rect 198792 201872 198798 201884
rect 211706 201872 211712 201884
rect 198792 201844 211712 201872
rect 198792 201832 198798 201844
rect 211706 201832 211712 201844
rect 211764 201832 211770 201884
rect 211801 201875 211859 201881
rect 211801 201841 211813 201875
rect 211847 201872 211859 201875
rect 215849 201875 215907 201881
rect 215849 201872 215861 201875
rect 211847 201844 215861 201872
rect 211847 201841 211859 201844
rect 211801 201835 211859 201841
rect 215849 201841 215861 201844
rect 215895 201841 215907 201875
rect 215849 201835 215907 201841
rect 215938 201832 215944 201884
rect 215996 201872 216002 201884
rect 216140 201872 216168 201912
rect 239125 201909 239137 201912
rect 239171 201909 239183 201943
rect 239125 201903 239183 201909
rect 239214 201900 239220 201952
rect 239272 201940 239278 201952
rect 240042 201940 240048 201952
rect 239272 201912 240048 201940
rect 239272 201900 239278 201912
rect 240042 201900 240048 201912
rect 240100 201900 240106 201952
rect 242066 201900 242072 201952
rect 242124 201940 242130 201952
rect 247678 201940 247684 201952
rect 242124 201912 247684 201940
rect 242124 201900 242130 201912
rect 247678 201900 247684 201912
rect 247736 201900 247742 201952
rect 253106 201900 253112 201952
rect 253164 201940 253170 201952
rect 253750 201940 253756 201952
rect 253164 201912 253756 201940
rect 253164 201900 253170 201912
rect 253750 201900 253756 201912
rect 253808 201900 253814 201952
rect 254854 201900 254860 201952
rect 254912 201940 254918 201952
rect 266906 201940 266912 201952
rect 254912 201912 266912 201940
rect 254912 201900 254918 201912
rect 266906 201900 266912 201912
rect 266964 201900 266970 201952
rect 297818 201900 297824 201952
rect 297876 201940 297882 201952
rect 303632 201940 303660 201980
rect 305638 201968 305644 201980
rect 305696 201968 305702 202020
rect 306285 202011 306343 202017
rect 306285 201977 306297 202011
rect 306331 202008 306343 202011
rect 315390 202008 315396 202020
rect 306331 201980 315396 202008
rect 306331 201977 306343 201980
rect 306285 201971 306343 201977
rect 315390 201968 315396 201980
rect 315448 201968 315454 202020
rect 318337 202011 318395 202017
rect 318337 201977 318349 202011
rect 318383 202008 318395 202011
rect 320634 202008 320640 202020
rect 318383 201980 320640 202008
rect 318383 201977 318395 201980
rect 318337 201971 318395 201977
rect 320634 201968 320640 201980
rect 320692 201968 320698 202020
rect 351730 201968 351736 202020
rect 351788 202008 351794 202020
rect 353312 202008 353340 202048
rect 417234 202036 417240 202048
rect 417292 202036 417298 202088
rect 351788 201980 353340 202008
rect 351788 201968 351794 201980
rect 365346 201968 365352 202020
rect 365404 202008 365410 202020
rect 369118 202008 369124 202020
rect 365404 201980 369124 202008
rect 365404 201968 365410 201980
rect 369118 201968 369124 201980
rect 369176 201968 369182 202020
rect 308493 201943 308551 201949
rect 308493 201940 308505 201943
rect 297876 201912 303660 201940
rect 306300 201912 308505 201940
rect 297876 201900 297882 201912
rect 215996 201844 216168 201872
rect 216217 201875 216275 201881
rect 215996 201832 216002 201844
rect 216217 201841 216229 201875
rect 216263 201872 216275 201875
rect 242158 201872 242164 201884
rect 216263 201844 242164 201872
rect 216263 201841 216275 201844
rect 216217 201835 216275 201841
rect 242158 201832 242164 201844
rect 242216 201832 242222 201884
rect 244829 201875 244887 201881
rect 244829 201841 244841 201875
rect 244875 201872 244887 201875
rect 251910 201872 251916 201884
rect 244875 201844 251916 201872
rect 244875 201841 244887 201844
rect 244829 201835 244887 201841
rect 251910 201832 251916 201844
rect 251968 201832 251974 201884
rect 256142 201832 256148 201884
rect 256200 201872 256206 201884
rect 264057 201875 264115 201881
rect 264057 201872 264069 201875
rect 256200 201844 264069 201872
rect 256200 201832 256206 201844
rect 264057 201841 264069 201844
rect 264103 201841 264115 201875
rect 267458 201872 267464 201884
rect 264057 201835 264115 201841
rect 264164 201844 267464 201872
rect 196802 201764 196808 201816
rect 196860 201804 196866 201816
rect 196860 201776 220492 201804
rect 196860 201764 196866 201776
rect 199286 201696 199292 201748
rect 199344 201736 199350 201748
rect 219526 201736 219532 201748
rect 199344 201708 219532 201736
rect 199344 201696 199350 201708
rect 219526 201696 219532 201708
rect 219584 201696 219590 201748
rect 220464 201736 220492 201776
rect 220814 201764 220820 201816
rect 220872 201804 220878 201816
rect 221274 201804 221280 201816
rect 220872 201776 221280 201804
rect 220872 201764 220878 201776
rect 221274 201764 221280 201776
rect 221332 201764 221338 201816
rect 229094 201764 229100 201816
rect 229152 201804 229158 201816
rect 232406 201804 232412 201816
rect 229152 201776 232412 201804
rect 229152 201764 229158 201776
rect 232406 201764 232412 201776
rect 232464 201764 232470 201816
rect 232498 201764 232504 201816
rect 232556 201804 232562 201816
rect 236730 201804 236736 201816
rect 232556 201776 236736 201804
rect 232556 201764 232562 201776
rect 236730 201764 236736 201776
rect 236788 201764 236794 201816
rect 236825 201807 236883 201813
rect 236825 201773 236837 201807
rect 236871 201804 236883 201807
rect 237377 201807 237435 201813
rect 237377 201804 237389 201807
rect 236871 201776 237389 201804
rect 236871 201773 236883 201776
rect 236825 201767 236883 201773
rect 237377 201773 237389 201776
rect 237423 201773 237435 201807
rect 237377 201767 237435 201773
rect 238110 201764 238116 201816
rect 238168 201804 238174 201816
rect 260834 201804 260840 201816
rect 238168 201776 260840 201804
rect 238168 201764 238174 201776
rect 260834 201764 260840 201776
rect 260892 201764 260898 201816
rect 223022 201736 223028 201748
rect 220464 201708 223028 201736
rect 223022 201696 223028 201708
rect 223080 201696 223086 201748
rect 223117 201739 223175 201745
rect 223117 201705 223129 201739
rect 223163 201736 223175 201739
rect 243170 201736 243176 201748
rect 223163 201708 243176 201736
rect 223163 201705 223175 201708
rect 223117 201699 223175 201705
rect 243170 201696 243176 201708
rect 243228 201696 243234 201748
rect 252462 201696 252468 201748
rect 252520 201736 252526 201748
rect 263594 201736 263600 201748
rect 252520 201708 263600 201736
rect 252520 201696 252526 201708
rect 263594 201696 263600 201708
rect 263652 201696 263658 201748
rect 199562 201628 199568 201680
rect 199620 201668 199626 201680
rect 218606 201668 218612 201680
rect 199620 201640 218612 201668
rect 199620 201628 199626 201640
rect 218606 201628 218612 201640
rect 218664 201628 218670 201680
rect 229738 201628 229744 201680
rect 229796 201668 229802 201680
rect 237374 201668 237380 201680
rect 229796 201640 237380 201668
rect 229796 201628 229802 201640
rect 237374 201628 237380 201640
rect 237432 201628 237438 201680
rect 238018 201628 238024 201680
rect 238076 201668 238082 201680
rect 259454 201668 259460 201680
rect 238076 201640 259460 201668
rect 238076 201628 238082 201640
rect 259454 201628 259460 201640
rect 259512 201628 259518 201680
rect 260098 201628 260104 201680
rect 260156 201668 260162 201680
rect 264164 201668 264192 201844
rect 267458 201832 267464 201844
rect 267516 201832 267522 201884
rect 297542 201832 297548 201884
rect 297600 201872 297606 201884
rect 306300 201872 306328 201912
rect 308493 201909 308505 201912
rect 308539 201909 308551 201943
rect 308493 201903 308551 201909
rect 311158 201900 311164 201952
rect 311216 201940 311222 201952
rect 330478 201940 330484 201952
rect 311216 201912 330484 201940
rect 311216 201900 311222 201912
rect 330478 201900 330484 201912
rect 330536 201900 330542 201952
rect 357894 201900 357900 201952
rect 357952 201940 357958 201952
rect 416958 201940 416964 201952
rect 357952 201912 416964 201940
rect 357952 201900 357958 201912
rect 416958 201900 416964 201912
rect 417016 201900 417022 201952
rect 313642 201872 313648 201884
rect 297600 201844 306328 201872
rect 306392 201844 313648 201872
rect 297600 201832 297606 201844
rect 266262 201764 266268 201816
rect 266320 201804 266326 201816
rect 269114 201804 269120 201816
rect 266320 201776 269120 201804
rect 266320 201764 266326 201776
rect 269114 201764 269120 201776
rect 269172 201764 269178 201816
rect 299566 201764 299572 201816
rect 299624 201804 299630 201816
rect 306285 201807 306343 201813
rect 306285 201804 306297 201807
rect 299624 201776 306297 201804
rect 299624 201764 299630 201776
rect 306285 201773 306297 201776
rect 306331 201773 306343 201807
rect 306285 201767 306343 201773
rect 265158 201696 265164 201748
rect 265216 201736 265222 201748
rect 267182 201736 267188 201748
rect 265216 201708 267188 201736
rect 265216 201696 265222 201708
rect 267182 201696 267188 201708
rect 267240 201696 267246 201748
rect 298370 201696 298376 201748
rect 298428 201736 298434 201748
rect 304905 201739 304963 201745
rect 304905 201736 304917 201739
rect 298428 201708 304917 201736
rect 298428 201696 298434 201708
rect 304905 201705 304917 201708
rect 304951 201705 304963 201739
rect 304905 201699 304963 201705
rect 260156 201640 264192 201668
rect 260156 201628 260162 201640
rect 267090 201628 267096 201680
rect 267148 201668 267154 201680
rect 268194 201668 268200 201680
rect 267148 201640 268200 201668
rect 267148 201628 267154 201640
rect 268194 201628 268200 201640
rect 268252 201628 268258 201680
rect 273622 201628 273628 201680
rect 273680 201668 273686 201680
rect 276658 201668 276664 201680
rect 273680 201640 276664 201668
rect 273680 201628 273686 201640
rect 276658 201628 276664 201640
rect 276716 201628 276722 201680
rect 299474 201628 299480 201680
rect 299532 201668 299538 201680
rect 306392 201668 306420 201844
rect 313642 201832 313648 201844
rect 313700 201832 313706 201884
rect 322750 201832 322756 201884
rect 322808 201872 322814 201884
rect 378226 201872 378232 201884
rect 322808 201844 378232 201872
rect 322808 201832 322814 201844
rect 378226 201832 378232 201844
rect 378284 201832 378290 201884
rect 412266 201832 412272 201884
rect 412324 201872 412330 201884
rect 416133 201875 416191 201881
rect 416133 201872 416145 201875
rect 412324 201844 416145 201872
rect 412324 201832 412330 201844
rect 416133 201841 416145 201844
rect 416179 201841 416191 201875
rect 416133 201835 416191 201841
rect 311986 201804 311992 201816
rect 307404 201776 311992 201804
rect 306466 201696 306472 201748
rect 306524 201736 306530 201748
rect 307294 201736 307300 201748
rect 306524 201708 307300 201736
rect 306524 201696 306530 201708
rect 307294 201696 307300 201708
rect 307352 201696 307358 201748
rect 299532 201640 306420 201668
rect 299532 201628 299538 201640
rect 126422 201560 126428 201612
rect 126480 201600 126486 201612
rect 134150 201600 134156 201612
rect 126480 201572 134156 201600
rect 126480 201560 126486 201572
rect 134150 201560 134156 201572
rect 134208 201560 134214 201612
rect 199654 201560 199660 201612
rect 199712 201600 199718 201612
rect 216858 201600 216864 201612
rect 199712 201572 216864 201600
rect 199712 201560 199718 201572
rect 216858 201560 216864 201572
rect 216916 201560 216922 201612
rect 216953 201603 217011 201609
rect 216953 201569 216965 201603
rect 216999 201600 217011 201603
rect 219253 201603 219311 201609
rect 219253 201600 219265 201603
rect 216999 201572 219265 201600
rect 216999 201569 217011 201572
rect 216953 201563 217011 201569
rect 219253 201569 219265 201572
rect 219299 201569 219311 201603
rect 219253 201563 219311 201569
rect 229189 201603 229247 201609
rect 229189 201569 229201 201603
rect 229235 201600 229247 201603
rect 233513 201603 233571 201609
rect 233513 201600 233525 201603
rect 229235 201572 233525 201600
rect 229235 201569 229247 201572
rect 229189 201563 229247 201569
rect 233513 201569 233525 201572
rect 233559 201569 233571 201603
rect 233513 201563 233571 201569
rect 233605 201603 233663 201609
rect 233605 201569 233617 201603
rect 233651 201600 233663 201603
rect 238202 201600 238208 201612
rect 233651 201572 238208 201600
rect 233651 201569 233663 201572
rect 233605 201563 233663 201569
rect 238202 201560 238208 201572
rect 238260 201560 238266 201612
rect 239125 201603 239183 201609
rect 239125 201569 239137 201603
rect 239171 201600 239183 201603
rect 247770 201600 247776 201612
rect 239171 201572 247776 201600
rect 239171 201569 239183 201572
rect 239125 201563 239183 201569
rect 247770 201560 247776 201572
rect 247828 201560 247834 201612
rect 255222 201560 255228 201612
rect 255280 201600 255286 201612
rect 258353 201603 258411 201609
rect 258353 201600 258365 201603
rect 255280 201572 258365 201600
rect 255280 201560 255286 201572
rect 258353 201569 258365 201572
rect 258399 201569 258411 201603
rect 258353 201563 258411 201569
rect 258718 201560 258724 201612
rect 258776 201600 258782 201612
rect 263870 201600 263876 201612
rect 258776 201572 263876 201600
rect 258776 201560 258782 201572
rect 263870 201560 263876 201572
rect 263928 201560 263934 201612
rect 266998 201560 267004 201612
rect 267056 201600 267062 201612
rect 267734 201600 267740 201612
rect 267056 201572 267740 201600
rect 267056 201560 267062 201572
rect 267734 201560 267740 201572
rect 267792 201560 267798 201612
rect 279234 201560 279240 201612
rect 279292 201600 279298 201612
rect 280062 201600 280068 201612
rect 279292 201572 280068 201600
rect 279292 201560 279298 201572
rect 280062 201560 280068 201572
rect 280120 201560 280126 201612
rect 282638 201560 282644 201612
rect 282696 201600 282702 201612
rect 287698 201600 287704 201612
rect 282696 201572 287704 201600
rect 282696 201560 282702 201572
rect 287698 201560 287704 201572
rect 287756 201560 287762 201612
rect 299290 201560 299296 201612
rect 299348 201600 299354 201612
rect 307404 201600 307432 201776
rect 311986 201764 311992 201776
rect 312044 201764 312050 201816
rect 366910 201764 366916 201816
rect 366968 201804 366974 201816
rect 420178 201804 420184 201816
rect 366968 201776 420184 201804
rect 366968 201764 366974 201776
rect 420178 201764 420184 201776
rect 420236 201764 420242 201816
rect 308398 201696 308404 201748
rect 308456 201736 308462 201748
rect 315669 201739 315727 201745
rect 315669 201736 315681 201739
rect 308456 201708 315681 201736
rect 308456 201696 308462 201708
rect 315669 201705 315681 201708
rect 315715 201705 315727 201739
rect 315669 201699 315727 201705
rect 364886 201696 364892 201748
rect 364944 201736 364950 201748
rect 381538 201736 381544 201748
rect 364944 201708 381544 201736
rect 364944 201696 364950 201708
rect 381538 201696 381544 201708
rect 381596 201696 381602 201748
rect 410150 201696 410156 201748
rect 410208 201736 410214 201748
rect 411162 201736 411168 201748
rect 410208 201708 411168 201736
rect 410208 201696 410214 201708
rect 411162 201696 411168 201708
rect 411220 201696 411226 201748
rect 374273 201671 374331 201677
rect 374273 201637 374285 201671
rect 374319 201668 374331 201671
rect 380066 201668 380072 201680
rect 374319 201640 380072 201668
rect 374319 201637 374331 201640
rect 374273 201631 374331 201637
rect 380066 201628 380072 201640
rect 380124 201628 380130 201680
rect 409230 201628 409236 201680
rect 409288 201668 409294 201680
rect 417053 201671 417111 201677
rect 417053 201668 417065 201671
rect 409288 201640 417065 201668
rect 409288 201628 409294 201640
rect 417053 201637 417065 201640
rect 417099 201637 417111 201671
rect 417053 201631 417111 201637
rect 299348 201572 307432 201600
rect 299348 201560 299354 201572
rect 314930 201560 314936 201612
rect 314988 201600 314994 201612
rect 380250 201600 380256 201612
rect 314988 201572 380256 201600
rect 314988 201560 314994 201572
rect 380250 201560 380256 201572
rect 380308 201560 380314 201612
rect 127618 201492 127624 201544
rect 127676 201532 127682 201544
rect 134334 201532 134340 201544
rect 127676 201504 134340 201532
rect 127676 201492 127682 201504
rect 134334 201492 134340 201504
rect 134392 201492 134398 201544
rect 198550 201492 198556 201544
rect 198608 201532 198614 201544
rect 202874 201532 202880 201544
rect 198608 201504 202880 201532
rect 198608 201492 198614 201504
rect 202874 201492 202880 201504
rect 202932 201492 202938 201544
rect 212442 201492 212448 201544
rect 212500 201532 212506 201544
rect 216217 201535 216275 201541
rect 216217 201532 216229 201535
rect 212500 201504 216229 201532
rect 212500 201492 212506 201504
rect 216217 201501 216229 201504
rect 216263 201501 216275 201535
rect 219345 201535 219403 201541
rect 219345 201532 219357 201535
rect 216217 201495 216275 201501
rect 216324 201504 219357 201532
rect 215849 201467 215907 201473
rect 215849 201433 215861 201467
rect 215895 201464 215907 201467
rect 216324 201464 216352 201504
rect 219345 201501 219357 201504
rect 219391 201501 219403 201535
rect 219345 201495 219403 201501
rect 220078 201492 220084 201544
rect 220136 201532 220142 201544
rect 223117 201535 223175 201541
rect 223117 201532 223129 201535
rect 220136 201504 223129 201532
rect 220136 201492 220142 201504
rect 223117 201501 223129 201504
rect 223163 201501 223175 201535
rect 223117 201495 223175 201501
rect 229097 201535 229155 201541
rect 229097 201501 229109 201535
rect 229143 201532 229155 201535
rect 238665 201535 238723 201541
rect 238665 201532 238677 201535
rect 229143 201504 238677 201532
rect 229143 201501 229155 201504
rect 229097 201495 229155 201501
rect 238665 201501 238677 201504
rect 238711 201501 238723 201535
rect 238665 201495 238723 201501
rect 239493 201535 239551 201541
rect 239493 201501 239505 201535
rect 239539 201532 239551 201535
rect 246482 201532 246488 201544
rect 239539 201504 246488 201532
rect 239539 201501 239551 201504
rect 239493 201495 239551 201501
rect 246482 201492 246488 201504
rect 246540 201492 246546 201544
rect 251450 201492 251456 201544
rect 251508 201532 251514 201544
rect 258813 201535 258871 201541
rect 258813 201532 258825 201535
rect 251508 201504 258825 201532
rect 251508 201492 251514 201504
rect 258813 201501 258825 201504
rect 258859 201501 258871 201535
rect 262217 201535 262275 201541
rect 262217 201532 262229 201535
rect 258813 201495 258871 201501
rect 258920 201504 262229 201532
rect 215895 201436 216352 201464
rect 215895 201433 215907 201436
rect 215849 201427 215907 201433
rect 258074 201424 258080 201476
rect 258132 201464 258138 201476
rect 258920 201464 258948 201504
rect 262217 201501 262229 201504
rect 262263 201501 262275 201535
rect 262217 201495 262275 201501
rect 264882 201492 264888 201544
rect 264940 201532 264946 201544
rect 266538 201532 266544 201544
rect 264940 201504 266544 201532
rect 264940 201492 264946 201504
rect 266538 201492 266544 201504
rect 266596 201492 266602 201544
rect 266630 201492 266636 201544
rect 266688 201532 266694 201544
rect 267274 201532 267280 201544
rect 266688 201504 267280 201532
rect 266688 201492 266694 201504
rect 267274 201492 267280 201504
rect 267332 201492 267338 201544
rect 282270 201492 282276 201544
rect 282328 201532 282334 201544
rect 284938 201532 284944 201544
rect 282328 201504 284944 201532
rect 282328 201492 282334 201504
rect 284938 201492 284944 201504
rect 284996 201492 285002 201544
rect 286226 201492 286232 201544
rect 286284 201532 286290 201544
rect 286962 201532 286968 201544
rect 286284 201504 286968 201532
rect 286284 201492 286290 201504
rect 286962 201492 286968 201504
rect 287020 201492 287026 201544
rect 302237 201535 302295 201541
rect 302237 201501 302249 201535
rect 302283 201532 302295 201535
rect 304994 201532 305000 201544
rect 302283 201504 305000 201532
rect 302283 201501 302295 201504
rect 302237 201495 302295 201501
rect 304994 201492 305000 201504
rect 305052 201492 305058 201544
rect 324038 201492 324044 201544
rect 324096 201532 324102 201544
rect 327074 201532 327080 201544
rect 324096 201504 327080 201532
rect 324096 201492 324102 201504
rect 327074 201492 327080 201504
rect 327132 201492 327138 201544
rect 355318 201492 355324 201544
rect 355376 201532 355382 201544
rect 355962 201532 355968 201544
rect 355376 201504 355968 201532
rect 355376 201492 355382 201504
rect 355962 201492 355968 201504
rect 356020 201492 356026 201544
rect 359642 201492 359648 201544
rect 359700 201532 359706 201544
rect 360102 201532 360108 201544
rect 359700 201504 360108 201532
rect 359700 201492 359706 201504
rect 360102 201492 360108 201504
rect 360160 201492 360166 201544
rect 360562 201492 360568 201544
rect 360620 201532 360626 201544
rect 361390 201532 361396 201544
rect 360620 201504 361396 201532
rect 360620 201492 360626 201504
rect 361390 201492 361396 201504
rect 361448 201492 361454 201544
rect 362310 201492 362316 201544
rect 362368 201532 362374 201544
rect 362770 201532 362776 201544
rect 362368 201504 362776 201532
rect 362368 201492 362374 201504
rect 362770 201492 362776 201504
rect 362828 201492 362834 201544
rect 258132 201436 258948 201464
rect 258132 201424 258138 201436
rect 215205 201399 215263 201405
rect 215205 201365 215217 201399
rect 215251 201396 215263 201399
rect 216953 201399 217011 201405
rect 216953 201396 216965 201399
rect 215251 201368 216965 201396
rect 215251 201365 215263 201368
rect 215205 201359 215263 201365
rect 216953 201365 216965 201368
rect 216999 201365 217011 201399
rect 216953 201359 217011 201365
rect 130562 201220 130568 201272
rect 130620 201260 130626 201272
rect 145558 201260 145564 201272
rect 130620 201232 145564 201260
rect 130620 201220 130626 201232
rect 145558 201220 145564 201232
rect 145616 201220 145622 201272
rect 133506 201152 133512 201204
rect 133564 201192 133570 201204
rect 153378 201192 153384 201204
rect 133564 201164 153384 201192
rect 133564 201152 133570 201164
rect 153378 201152 153384 201164
rect 153436 201152 153442 201204
rect 266446 201152 266452 201204
rect 266504 201192 266510 201204
rect 267642 201192 267648 201204
rect 266504 201164 267648 201192
rect 266504 201152 266510 201164
rect 267642 201152 267648 201164
rect 267700 201152 267706 201204
rect 3878 201084 3884 201136
rect 3936 201124 3942 201136
rect 436554 201124 436560 201136
rect 3936 201096 436560 201124
rect 3936 201084 3942 201096
rect 436554 201084 436560 201096
rect 436612 201084 436618 201136
rect 3602 201016 3608 201068
rect 3660 201056 3666 201068
rect 436462 201056 436468 201068
rect 3660 201028 436468 201056
rect 3660 201016 3666 201028
rect 436462 201016 436468 201028
rect 436520 201016 436526 201068
rect 3418 200948 3424 201000
rect 3476 200988 3482 201000
rect 436370 200988 436376 201000
rect 3476 200960 436376 200988
rect 3476 200948 3482 200960
rect 436370 200948 436376 200960
rect 436428 200948 436434 201000
rect 132402 200880 132408 200932
rect 132460 200920 132466 200932
rect 580258 200920 580264 200932
rect 132460 200892 580264 200920
rect 132460 200880 132466 200892
rect 580258 200880 580264 200892
rect 580316 200880 580322 200932
rect 132218 200812 132224 200864
rect 132276 200852 132282 200864
rect 580442 200852 580448 200864
rect 132276 200824 580448 200852
rect 132276 200812 132282 200824
rect 580442 200812 580448 200824
rect 580500 200812 580506 200864
rect 131390 200744 131396 200796
rect 131448 200784 131454 200796
rect 580350 200784 580356 200796
rect 131448 200756 580356 200784
rect 131448 200744 131454 200756
rect 580350 200744 580356 200756
rect 580408 200744 580414 200796
rect 504174 200404 504180 200456
rect 504232 200444 504238 200456
rect 504450 200444 504456 200456
rect 504232 200416 504456 200444
rect 504232 200404 504238 200416
rect 504450 200404 504456 200416
rect 504508 200404 504514 200456
rect 209866 200200 209872 200252
rect 209924 200240 209930 200252
rect 210280 200240 210286 200252
rect 209924 200212 210286 200240
rect 209924 200200 209930 200212
rect 210280 200200 210286 200212
rect 210338 200200 210344 200252
rect 213914 200200 213920 200252
rect 213972 200240 213978 200252
rect 214604 200240 214610 200252
rect 213972 200212 214610 200240
rect 213972 200200 213978 200212
rect 214604 200200 214610 200212
rect 214662 200200 214668 200252
rect 3234 200132 3240 200184
rect 3292 200172 3298 200184
rect 436646 200172 436652 200184
rect 3292 200144 436652 200172
rect 3292 200132 3298 200144
rect 436646 200132 436652 200144
rect 436704 200132 436710 200184
rect 128538 200064 128544 200116
rect 128596 200104 128602 200116
rect 128906 200104 128912 200116
rect 128596 200076 128912 200104
rect 128596 200064 128602 200076
rect 128906 200064 128912 200076
rect 128964 200064 128970 200116
rect 266446 200064 266452 200116
rect 266504 200104 266510 200116
rect 266722 200104 266728 200116
rect 266504 200076 266728 200104
rect 266504 200064 266510 200076
rect 266722 200064 266728 200076
rect 266780 200064 266786 200116
rect 238754 199860 238760 199912
rect 238812 199900 238818 199912
rect 239490 199900 239496 199912
rect 238812 199872 239496 199900
rect 238812 199860 238818 199872
rect 239490 199860 239496 199872
rect 239548 199860 239554 199912
rect 243078 199860 243084 199912
rect 243136 199900 243142 199912
rect 243814 199900 243820 199912
rect 243136 199872 243820 199900
rect 243136 199860 243142 199872
rect 243814 199860 243820 199872
rect 243872 199860 243878 199912
rect 133598 199792 133604 199844
rect 133656 199832 133662 199844
rect 580258 199832 580264 199844
rect 133656 199804 580264 199832
rect 133656 199792 133662 199804
rect 580258 199792 580264 199804
rect 580316 199792 580322 199844
rect 131390 198296 131396 198348
rect 131448 198336 131454 198348
rect 131485 198339 131543 198345
rect 131485 198336 131497 198339
rect 131448 198308 131497 198336
rect 131448 198296 131454 198308
rect 131485 198305 131497 198308
rect 131531 198305 131543 198339
rect 131485 198299 131543 198305
rect 3418 197344 3424 197396
rect 3476 197384 3482 197396
rect 131390 197384 131396 197396
rect 3476 197356 131396 197384
rect 3476 197344 3482 197356
rect 131390 197344 131396 197356
rect 131448 197344 131454 197396
rect 5350 196256 5356 196308
rect 5408 196296 5414 196308
rect 131390 196296 131396 196308
rect 5408 196268 131396 196296
rect 5408 196256 5414 196268
rect 131390 196256 131396 196268
rect 131448 196256 131454 196308
rect 17218 196052 17224 196104
rect 17276 196092 17282 196104
rect 130470 196092 130476 196104
rect 17276 196064 130476 196092
rect 17276 196052 17282 196064
rect 130470 196052 130476 196064
rect 130528 196052 130534 196104
rect 131758 196092 131764 196104
rect 131719 196064 131764 196092
rect 131758 196052 131764 196064
rect 131816 196052 131822 196104
rect 132862 196092 132868 196104
rect 132823 196064 132868 196092
rect 132862 196052 132868 196064
rect 132920 196052 132926 196104
rect 131390 195984 131396 196036
rect 131448 196024 131454 196036
rect 131485 196027 131543 196033
rect 131485 196024 131497 196027
rect 131448 195996 131497 196024
rect 131448 195984 131454 195996
rect 131485 195993 131497 195996
rect 131531 195993 131543 196027
rect 131485 195987 131543 195993
rect 126422 195916 126428 195968
rect 126480 195956 126486 195968
rect 126606 195956 126612 195968
rect 126480 195928 126612 195956
rect 126480 195916 126486 195928
rect 126606 195916 126612 195928
rect 126664 195916 126670 195968
rect 131758 195956 131764 195968
rect 131719 195928 131764 195956
rect 131758 195916 131764 195928
rect 131816 195916 131822 195968
rect 132862 195956 132868 195968
rect 132823 195928 132868 195956
rect 132862 195916 132868 195928
rect 132920 195916 132926 195968
rect 15838 194556 15844 194608
rect 15896 194596 15902 194608
rect 130470 194596 130476 194608
rect 15896 194568 130476 194596
rect 15896 194556 15902 194568
rect 130470 194556 130476 194568
rect 130528 194556 130534 194608
rect 14458 194420 14464 194472
rect 14516 194460 14522 194472
rect 130470 194460 130476 194472
rect 14516 194432 130476 194460
rect 14516 194420 14522 194432
rect 130470 194420 130476 194432
rect 130528 194420 130534 194472
rect 5258 193128 5264 193180
rect 5316 193168 5322 193180
rect 130378 193168 130384 193180
rect 5316 193140 130384 193168
rect 5316 193128 5322 193140
rect 130378 193128 130384 193140
rect 130436 193128 130442 193180
rect 5442 193060 5448 193112
rect 5500 193100 5506 193112
rect 130470 193100 130476 193112
rect 5500 193072 130476 193100
rect 5500 193060 5506 193072
rect 130470 193060 130476 193072
rect 130528 193060 130534 193112
rect 5166 191768 5172 191820
rect 5224 191808 5230 191820
rect 130470 191808 130476 191820
rect 5224 191780 130476 191808
rect 5224 191768 5230 191780
rect 130470 191768 130476 191780
rect 130528 191768 130534 191820
rect 5074 190408 5080 190460
rect 5132 190448 5138 190460
rect 130470 190448 130476 190460
rect 5132 190420 130476 190448
rect 5132 190408 5138 190420
rect 130470 190408 130476 190420
rect 130528 190408 130534 190460
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 130378 189020 130384 189032
rect 3568 188992 130384 189020
rect 3568 188980 3574 188992
rect 130378 188980 130384 188992
rect 130436 188980 130442 189032
rect 4982 188912 4988 188964
rect 5040 188952 5046 188964
rect 130470 188952 130476 188964
rect 5040 188924 130476 188952
rect 5040 188912 5046 188924
rect 130470 188912 130476 188924
rect 130528 188912 130534 188964
rect 4890 187620 4896 187672
rect 4948 187660 4954 187672
rect 130470 187660 130476 187672
rect 4948 187632 130476 187660
rect 4948 187620 4954 187632
rect 130470 187620 130476 187632
rect 130528 187620 130534 187672
rect 4798 186260 4804 186312
rect 4856 186300 4862 186312
rect 131117 186303 131175 186309
rect 4856 186272 131068 186300
rect 4856 186260 4862 186272
rect 131040 186232 131068 186272
rect 131117 186269 131129 186303
rect 131163 186300 131175 186303
rect 131206 186300 131212 186312
rect 131163 186272 131212 186300
rect 131163 186269 131175 186272
rect 131117 186263 131175 186269
rect 131206 186260 131212 186272
rect 131264 186260 131270 186312
rect 131040 186204 131252 186232
rect 131224 186176 131252 186204
rect 131206 186124 131212 186176
rect 131264 186124 131270 186176
rect 13078 184832 13084 184884
rect 13136 184872 13142 184884
rect 131206 184872 131212 184884
rect 13136 184844 131212 184872
rect 13136 184832 13142 184844
rect 131206 184832 131212 184844
rect 131264 184832 131270 184884
rect 72418 183472 72424 183524
rect 72476 183512 72482 183524
rect 131206 183512 131212 183524
rect 72476 183484 131212 183512
rect 72476 183472 72482 183484
rect 131206 183472 131212 183484
rect 131264 183472 131270 183524
rect 131117 183379 131175 183385
rect 131117 183345 131129 183379
rect 131163 183376 131175 183379
rect 131206 183376 131212 183388
rect 131163 183348 131212 183376
rect 131163 183345 131175 183348
rect 131117 183339 131175 183345
rect 131206 183336 131212 183348
rect 131264 183336 131270 183388
rect 132862 181432 132868 181484
rect 132920 181472 132926 181484
rect 133322 181472 133328 181484
rect 132920 181444 133328 181472
rect 132920 181432 132926 181444
rect 133322 181432 133328 181444
rect 133380 181432 133386 181484
rect 2866 180752 2872 180804
rect 2924 180792 2930 180804
rect 15838 180792 15844 180804
rect 2924 180764 15844 180792
rect 2924 180752 2930 180764
rect 15838 180752 15844 180764
rect 15896 180752 15902 180804
rect 128906 180792 128912 180804
rect 128867 180764 128912 180792
rect 128906 180752 128912 180764
rect 128964 180752 128970 180804
rect 126422 176604 126428 176656
rect 126480 176644 126486 176656
rect 126606 176644 126612 176656
rect 126480 176616 126612 176644
rect 126480 176604 126486 176616
rect 126606 176604 126612 176616
rect 126664 176604 126670 176656
rect 504450 173884 504456 173936
rect 504508 173924 504514 173936
rect 504634 173924 504640 173936
rect 504508 173896 504640 173924
rect 504508 173884 504514 173896
rect 504634 173884 504640 173896
rect 504692 173884 504698 173936
rect 128909 171139 128967 171145
rect 128909 171105 128921 171139
rect 128955 171136 128967 171139
rect 128998 171136 129004 171148
rect 128955 171108 129004 171136
rect 128955 171105 128967 171108
rect 128909 171099 128967 171105
rect 128998 171096 129004 171108
rect 129056 171096 129062 171148
rect 132954 168580 132960 168632
rect 133012 168620 133018 168632
rect 133322 168620 133328 168632
rect 133012 168592 133328 168620
rect 133012 168580 133018 168592
rect 133322 168580 133328 168592
rect 133380 168580 133386 168632
rect 128906 164228 128912 164280
rect 128964 164268 128970 164280
rect 128998 164268 129004 164280
rect 128964 164240 129004 164268
rect 128964 164228 128970 164240
rect 128998 164228 129004 164240
rect 129056 164228 129062 164280
rect 504174 164160 504180 164212
rect 504232 164200 504238 164212
rect 504358 164200 504364 164212
rect 504232 164172 504364 164200
rect 504232 164160 504238 164172
rect 504358 164160 504364 164172
rect 504416 164160 504422 164212
rect 126514 161440 126520 161492
rect 126572 161480 126578 161492
rect 126606 161480 126612 161492
rect 126572 161452 126612 161480
rect 126572 161440 126578 161452
rect 126606 161440 126612 161452
rect 126664 161440 126670 161492
rect 128906 157468 128912 157480
rect 128832 157440 128912 157468
rect 128832 157276 128860 157440
rect 128906 157428 128912 157440
rect 128964 157428 128970 157480
rect 436830 157360 436836 157412
rect 436888 157400 436894 157412
rect 580166 157400 580172 157412
rect 436888 157372 580172 157400
rect 436888 157360 436894 157372
rect 580166 157360 580172 157372
rect 580224 157360 580230 157412
rect 131206 157332 131212 157344
rect 131167 157304 131212 157332
rect 131206 157292 131212 157304
rect 131264 157292 131270 157344
rect 128814 157224 128820 157276
rect 128872 157224 128878 157276
rect 131114 156272 131120 156324
rect 131172 156312 131178 156324
rect 131172 156284 131436 156312
rect 131172 156272 131178 156284
rect 3510 156068 3516 156120
rect 3568 156108 3574 156120
rect 131298 156108 131304 156120
rect 3568 156080 131304 156108
rect 3568 156068 3574 156080
rect 131298 156068 131304 156080
rect 131356 156068 131362 156120
rect 3234 156000 3240 156052
rect 3292 156040 3298 156052
rect 131114 156040 131120 156052
rect 3292 156012 131120 156040
rect 3292 156000 3298 156012
rect 131114 156000 131120 156012
rect 131172 156000 131178 156052
rect 131298 155932 131304 155984
rect 131356 155972 131362 155984
rect 131408 155972 131436 156284
rect 131356 155944 131436 155972
rect 131356 155932 131362 155944
rect 3602 155864 3608 155916
rect 3660 155904 3666 155916
rect 131114 155904 131120 155916
rect 3660 155876 131120 155904
rect 3660 155864 3666 155876
rect 131114 155864 131120 155876
rect 131172 155864 131178 155916
rect 436094 155184 436100 155236
rect 436152 155224 436158 155236
rect 438118 155224 438124 155236
rect 436152 155196 438124 155224
rect 436152 155184 436158 155196
rect 438118 155184 438124 155196
rect 438176 155184 438182 155236
rect 57977 154547 58035 154553
rect 57977 154544 57989 154547
rect 31680 154516 57989 154544
rect 31680 154476 31708 154516
rect 57977 154513 57989 154516
rect 58023 154513 58035 154547
rect 99285 154547 99343 154553
rect 99285 154544 99297 154547
rect 57977 154507 58035 154513
rect 89640 154516 99297 154544
rect 22112 154448 31708 154476
rect 67545 154479 67603 154485
rect 22112 154408 22140 154448
rect 67545 154445 67557 154479
rect 67591 154476 67603 154479
rect 89640 154476 89668 154516
rect 99285 154513 99297 154516
rect 99331 154513 99343 154547
rect 99285 154507 99343 154513
rect 67591 154448 70348 154476
rect 67591 154445 67603 154448
rect 67545 154439 67603 154445
rect 14476 154380 22140 154408
rect 70320 154408 70348 154448
rect 86880 154448 89668 154476
rect 99469 154479 99527 154485
rect 80057 154411 80115 154417
rect 80057 154408 80069 154411
rect 70320 154380 80069 154408
rect 9600 154312 9720 154340
rect 3326 154232 3332 154284
rect 3384 154272 3390 154284
rect 9600 154272 9628 154312
rect 3384 154244 9628 154272
rect 9692 154272 9720 154312
rect 14476 154272 14504 154380
rect 80057 154377 80069 154380
rect 80103 154377 80115 154411
rect 80057 154371 80115 154377
rect 80149 154411 80207 154417
rect 80149 154377 80161 154411
rect 80195 154408 80207 154411
rect 86880 154408 86908 154448
rect 99469 154445 99481 154479
rect 99515 154476 99527 154479
rect 118605 154479 118663 154485
rect 118605 154476 118617 154479
rect 99515 154448 118617 154476
rect 99515 154445 99527 154448
rect 99469 154439 99527 154445
rect 118605 154445 118617 154448
rect 118651 154445 118663 154479
rect 118605 154439 118663 154445
rect 80195 154380 86908 154408
rect 118789 154411 118847 154417
rect 80195 154377 80207 154380
rect 80149 154371 80207 154377
rect 118789 154377 118801 154411
rect 118835 154408 118847 154411
rect 124214 154408 124220 154420
rect 118835 154380 124220 154408
rect 118835 154377 118847 154380
rect 118789 154371 118847 154377
rect 124214 154368 124220 154380
rect 124272 154368 124278 154420
rect 57977 154343 58035 154349
rect 57977 154309 57989 154343
rect 58023 154340 58035 154343
rect 67545 154343 67603 154349
rect 67545 154340 67557 154343
rect 58023 154312 67557 154340
rect 58023 154309 58035 154312
rect 57977 154303 58035 154309
rect 67545 154309 67557 154312
rect 67591 154309 67603 154343
rect 67545 154303 67603 154309
rect 9692 154244 14504 154272
rect 3384 154232 3390 154244
rect 4062 153144 4068 153196
rect 4120 153184 4126 153196
rect 131114 153184 131120 153196
rect 4120 153156 131120 153184
rect 4120 153144 4126 153156
rect 131114 153144 131120 153156
rect 131172 153144 131178 153196
rect 437382 153144 437388 153196
rect 437440 153184 437446 153196
rect 447778 153184 447784 153196
rect 437440 153156 447784 153184
rect 437440 153144 437446 153156
rect 447778 153144 447784 153156
rect 447836 153144 447842 153196
rect 32401 153119 32459 153125
rect 32401 153085 32413 153119
rect 32447 153116 32459 153119
rect 108945 153119 109003 153125
rect 108945 153116 108957 153119
rect 32447 153088 60780 153116
rect 32447 153085 32459 153088
rect 32401 153079 32459 153085
rect 22741 153051 22799 153057
rect 22741 153017 22753 153051
rect 22787 153048 22799 153051
rect 27617 153051 27675 153057
rect 27617 153048 27629 153051
rect 22787 153020 27629 153048
rect 22787 153017 22799 153020
rect 22741 153011 22799 153017
rect 27617 153017 27629 153020
rect 27663 153017 27675 153051
rect 60752 153048 60780 153088
rect 89640 153088 108957 153116
rect 86865 153051 86923 153057
rect 60752 153020 70348 153048
rect 27617 153011 27675 153017
rect 3970 152940 3976 152992
rect 4028 152980 4034 152992
rect 70320 152980 70348 153020
rect 86865 153017 86877 153051
rect 86911 153048 86923 153051
rect 89640 153048 89668 153088
rect 108945 153085 108957 153088
rect 108991 153085 109003 153119
rect 108945 153079 109003 153085
rect 109037 153119 109095 153125
rect 109037 153085 109049 153119
rect 109083 153116 109095 153119
rect 131298 153116 131304 153128
rect 109083 153088 118740 153116
rect 131259 153088 131304 153116
rect 109083 153085 109095 153088
rect 109037 153079 109095 153085
rect 86911 153020 89668 153048
rect 118712 153048 118740 153088
rect 131298 153076 131304 153088
rect 131356 153076 131362 153128
rect 118712 153020 128308 153048
rect 86911 153017 86923 153020
rect 86865 153011 86923 153017
rect 77297 152983 77355 152989
rect 77297 152980 77309 152983
rect 4028 152952 12204 152980
rect 70320 152952 77309 152980
rect 4028 152940 4034 152952
rect 12176 152912 12204 152952
rect 77297 152949 77309 152952
rect 77343 152949 77355 152983
rect 77297 152943 77355 152949
rect 17957 152915 18015 152921
rect 17957 152912 17969 152915
rect 12176 152884 17969 152912
rect 17957 152881 17969 152884
rect 18003 152881 18015 152915
rect 17957 152875 18015 152881
rect 27617 152915 27675 152921
rect 27617 152881 27629 152915
rect 27663 152912 27675 152915
rect 32401 152915 32459 152921
rect 32401 152912 32413 152915
rect 27663 152884 32413 152912
rect 27663 152881 27675 152884
rect 27617 152875 27675 152881
rect 32401 152881 32413 152884
rect 32447 152881 32459 152915
rect 128280 152912 128308 153020
rect 131206 152912 131212 152924
rect 128280 152884 131212 152912
rect 32401 152875 32459 152881
rect 131206 152872 131212 152884
rect 131264 152872 131270 152924
rect 77297 152847 77355 152853
rect 77297 152813 77309 152847
rect 77343 152844 77355 152847
rect 86865 152847 86923 152853
rect 86865 152844 86877 152847
rect 77343 152816 86877 152844
rect 77343 152813 77355 152816
rect 77297 152807 77355 152813
rect 86865 152813 86877 152816
rect 86911 152813 86923 152847
rect 86865 152807 86923 152813
rect 17957 152779 18015 152785
rect 17957 152745 17969 152779
rect 18003 152776 18015 152779
rect 22741 152779 22799 152785
rect 22741 152776 22753 152779
rect 18003 152748 22753 152776
rect 18003 152745 18015 152748
rect 17957 152739 18015 152745
rect 22741 152745 22753 152748
rect 22787 152745 22799 152779
rect 22741 152739 22799 152745
rect 131298 151892 131304 151904
rect 131259 151864 131304 151892
rect 131298 151852 131304 151864
rect 131356 151852 131362 151904
rect 3786 151716 3792 151768
rect 3844 151756 3850 151768
rect 131114 151756 131120 151768
rect 3844 151728 131120 151756
rect 3844 151716 3850 151728
rect 131114 151716 131120 151728
rect 131172 151716 131178 151768
rect 3694 150356 3700 150408
rect 3752 150396 3758 150408
rect 131114 150396 131120 150408
rect 3752 150368 131120 150396
rect 3752 150356 3758 150368
rect 131114 150356 131120 150368
rect 131172 150356 131178 150408
rect 437382 150356 437388 150408
rect 437440 150396 437446 150408
rect 446398 150396 446404 150408
rect 437440 150368 446404 150396
rect 437440 150356 437446 150368
rect 446398 150356 446404 150368
rect 446456 150356 446462 150408
rect 28258 148996 28264 149048
rect 28316 149036 28322 149048
rect 28316 149008 131252 149036
rect 28316 148996 28322 149008
rect 31018 148928 31024 148980
rect 31076 148968 31082 148980
rect 131114 148968 131120 148980
rect 31076 148940 131120 148968
rect 31076 148928 31082 148940
rect 131114 148928 131120 148940
rect 131172 148928 131178 148980
rect 131224 148900 131252 149008
rect 436094 148996 436100 149048
rect 436152 149036 436158 149048
rect 445018 149036 445024 149048
rect 436152 149008 445024 149036
rect 436152 148996 436158 149008
rect 445018 148996 445024 149008
rect 445076 148996 445082 149048
rect 131132 148872 131252 148900
rect 131132 148640 131160 148872
rect 131114 148588 131120 148640
rect 131172 148588 131178 148640
rect 131206 147676 131212 147688
rect 131167 147648 131212 147676
rect 131206 147636 131212 147648
rect 131264 147636 131270 147688
rect 21358 147568 21364 147620
rect 21416 147608 21422 147620
rect 131114 147608 131120 147620
rect 21416 147580 131120 147608
rect 21416 147568 21422 147580
rect 131114 147568 131120 147580
rect 131172 147568 131178 147620
rect 19978 146208 19984 146260
rect 20036 146248 20042 146260
rect 131114 146248 131120 146260
rect 20036 146220 131120 146248
rect 20036 146208 20042 146220
rect 131114 146208 131120 146220
rect 131172 146208 131178 146260
rect 437382 146140 437388 146192
rect 437440 146180 437446 146192
rect 442258 146180 442264 146192
rect 437440 146152 442264 146180
rect 437440 146140 437446 146152
rect 442258 146140 442264 146152
rect 442316 146140 442322 146192
rect 67637 144891 67695 144897
rect 67637 144857 67649 144891
rect 67683 144888 67695 144891
rect 79965 144891 80023 144897
rect 79965 144888 79977 144891
rect 67683 144860 79977 144888
rect 67683 144857 67695 144860
rect 67637 144851 67695 144857
rect 79965 144857 79977 144860
rect 80011 144857 80023 144891
rect 79965 144851 80023 144857
rect 96525 144891 96583 144897
rect 96525 144857 96537 144891
rect 96571 144888 96583 144891
rect 99285 144891 99343 144897
rect 99285 144888 99297 144891
rect 96571 144860 99297 144888
rect 96571 144857 96583 144860
rect 96525 144851 96583 144857
rect 99285 144857 99297 144860
rect 99331 144857 99343 144891
rect 99285 144851 99343 144857
rect 109037 144891 109095 144897
rect 109037 144857 109049 144891
rect 109083 144888 109095 144891
rect 118605 144891 118663 144897
rect 118605 144888 118617 144891
rect 109083 144860 118617 144888
rect 109083 144857 109095 144860
rect 109037 144851 109095 144857
rect 118605 144857 118617 144860
rect 118651 144857 118663 144891
rect 118605 144851 118663 144857
rect 437014 144848 437020 144900
rect 437072 144888 437078 144900
rect 514018 144888 514024 144900
rect 437072 144860 514024 144888
rect 437072 144848 437078 144860
rect 514018 144848 514024 144860
rect 514076 144848 514082 144900
rect 99469 144823 99527 144829
rect 99469 144789 99481 144823
rect 99515 144820 99527 144823
rect 99515 144792 108988 144820
rect 99515 144789 99527 144792
rect 99469 144783 99527 144789
rect 38565 144755 38623 144761
rect 38565 144721 38577 144755
rect 38611 144752 38623 144755
rect 41325 144755 41383 144761
rect 41325 144752 41337 144755
rect 38611 144724 41337 144752
rect 38611 144721 38623 144724
rect 38565 144715 38623 144721
rect 41325 144721 41337 144724
rect 41371 144721 41383 144755
rect 41325 144715 41383 144721
rect 41417 144755 41475 144761
rect 41417 144721 41429 144755
rect 41463 144752 41475 144755
rect 57885 144755 57943 144761
rect 41463 144724 42656 144752
rect 41463 144721 41475 144724
rect 41417 144715 41475 144721
rect 24762 144644 24768 144696
rect 24820 144684 24826 144696
rect 28997 144687 29055 144693
rect 28997 144684 29009 144687
rect 24820 144656 29009 144684
rect 24820 144644 24826 144656
rect 28997 144653 29009 144656
rect 29043 144653 29055 144687
rect 42628 144684 42656 144724
rect 57885 144721 57897 144755
rect 57931 144752 57943 144755
rect 60645 144755 60703 144761
rect 60645 144752 60657 144755
rect 57931 144724 60657 144752
rect 57931 144721 57943 144724
rect 57885 144715 57943 144721
rect 60645 144721 60657 144724
rect 60691 144721 60703 144755
rect 60645 144715 60703 144721
rect 60737 144755 60795 144761
rect 60737 144721 60749 144755
rect 60783 144752 60795 144755
rect 80149 144755 80207 144761
rect 60783 144724 61976 144752
rect 60783 144721 60795 144724
rect 60737 144715 60795 144721
rect 48317 144687 48375 144693
rect 48317 144684 48329 144687
rect 42628 144656 48329 144684
rect 28997 144647 29055 144653
rect 48317 144653 48329 144656
rect 48363 144653 48375 144687
rect 61948 144684 61976 144724
rect 80149 144721 80161 144755
rect 80195 144752 80207 144755
rect 86957 144755 87015 144761
rect 86957 144752 86969 144755
rect 80195 144724 86969 144752
rect 80195 144721 80207 144724
rect 80149 144715 80207 144721
rect 86957 144721 86969 144724
rect 87003 144721 87015 144755
rect 108960 144752 108988 144792
rect 109037 144755 109095 144761
rect 109037 144752 109049 144755
rect 108960 144724 109049 144752
rect 86957 144715 87015 144721
rect 109037 144721 109049 144724
rect 109083 144721 109095 144755
rect 109037 144715 109095 144721
rect 118789 144755 118847 144761
rect 118789 144721 118801 144755
rect 118835 144752 118847 144755
rect 128170 144752 128176 144764
rect 118835 144724 128176 144752
rect 118835 144721 118847 144724
rect 118789 144715 118847 144721
rect 128170 144712 128176 144724
rect 128228 144712 128234 144764
rect 67637 144687 67695 144693
rect 67637 144684 67649 144687
rect 61948 144656 67649 144684
rect 48317 144647 48375 144653
rect 67637 144653 67649 144656
rect 67683 144653 67695 144687
rect 67637 144647 67695 144653
rect 86957 144619 87015 144625
rect 86957 144585 86969 144619
rect 87003 144616 87015 144619
rect 96525 144619 96583 144625
rect 96525 144616 96537 144619
rect 87003 144588 96537 144616
rect 87003 144585 87015 144588
rect 86957 144579 87015 144585
rect 96525 144585 96537 144588
rect 96571 144585 96583 144619
rect 96525 144579 96583 144585
rect 28997 144551 29055 144557
rect 28997 144517 29009 144551
rect 29043 144548 29055 144551
rect 38565 144551 38623 144557
rect 38565 144548 38577 144551
rect 29043 144520 38577 144548
rect 29043 144517 29055 144520
rect 28997 144511 29055 144517
rect 38565 144517 38577 144520
rect 38611 144517 38623 144551
rect 38565 144511 38623 144517
rect 48317 144551 48375 144557
rect 48317 144517 48329 144551
rect 48363 144548 48375 144551
rect 57885 144551 57943 144557
rect 57885 144548 57897 144551
rect 48363 144520 57897 144548
rect 48363 144517 48375 144520
rect 48317 144511 48375 144517
rect 57885 144517 57897 144520
rect 57931 144517 57943 144551
rect 57885 144511 57943 144517
rect 126238 144372 126244 144424
rect 126296 144412 126302 144424
rect 131114 144412 131120 144424
rect 126296 144384 131120 144412
rect 126296 144372 126302 144384
rect 131114 144372 131120 144384
rect 131172 144372 131178 144424
rect 132773 143599 132831 143605
rect 132773 143565 132785 143599
rect 132819 143596 132831 143599
rect 132862 143596 132868 143608
rect 132819 143568 132868 143596
rect 132819 143565 132831 143568
rect 132773 143559 132831 143565
rect 132862 143556 132868 143568
rect 132920 143556 132926 143608
rect 132770 142168 132776 142180
rect 132731 142140 132776 142168
rect 132770 142128 132776 142140
rect 132828 142128 132834 142180
rect 128814 142100 128820 142112
rect 128775 142072 128820 142100
rect 128814 142060 128820 142072
rect 128872 142060 128878 142112
rect 436094 142060 436100 142112
rect 436152 142100 436158 142112
rect 438210 142100 438216 142112
rect 436152 142072 438216 142100
rect 436152 142060 436158 142072
rect 438210 142060 438216 142072
rect 438268 142060 438274 142112
rect 437382 137912 437388 137964
rect 437440 137952 437446 137964
rect 580534 137952 580540 137964
rect 437440 137924 580540 137952
rect 437440 137912 437446 137924
rect 580534 137912 580540 137924
rect 580592 137912 580598 137964
rect 3326 136552 3332 136604
rect 3384 136592 3390 136604
rect 17218 136592 17224 136604
rect 3384 136564 17224 136592
rect 3384 136552 3390 136564
rect 17218 136552 17224 136564
rect 17276 136552 17282 136604
rect 437014 136552 437020 136604
rect 437072 136592 437078 136604
rect 504450 136592 504456 136604
rect 437072 136564 504456 136592
rect 437072 136552 437078 136564
rect 504450 136552 504456 136564
rect 504508 136552 504514 136604
rect 130654 135532 130660 135584
rect 130712 135572 130718 135584
rect 132310 135572 132316 135584
rect 130712 135544 132316 135572
rect 130712 135532 130718 135544
rect 132310 135532 132316 135544
rect 132368 135532 132374 135584
rect 128814 133872 128820 133884
rect 128775 133844 128820 133872
rect 128814 133832 128820 133844
rect 128872 133832 128878 133884
rect 131114 133832 131120 133884
rect 131172 133872 131178 133884
rect 131298 133872 131304 133884
rect 131172 133844 131304 133872
rect 131172 133832 131178 133844
rect 131298 133832 131304 133844
rect 131356 133832 131362 133884
rect 437382 133832 437388 133884
rect 437440 133872 437446 133884
rect 580626 133872 580632 133884
rect 437440 133844 580632 133872
rect 437440 133832 437446 133844
rect 580626 133832 580632 133844
rect 580684 133832 580690 133884
rect 132310 132404 132316 132456
rect 132368 132444 132374 132456
rect 132368 132416 132540 132444
rect 132368 132404 132374 132416
rect 132512 132376 132540 132416
rect 437382 132404 437388 132456
rect 437440 132444 437446 132456
rect 580718 132444 580724 132456
rect 437440 132416 580724 132444
rect 437440 132404 437446 132416
rect 580718 132404 580724 132416
rect 580776 132404 580782 132456
rect 133138 132376 133144 132388
rect 132512 132348 133144 132376
rect 133138 132336 133144 132348
rect 133196 132336 133202 132388
rect 437382 129684 437388 129736
rect 437440 129724 437446 129736
rect 580810 129724 580816 129736
rect 437440 129696 580816 129724
rect 437440 129684 437446 129696
rect 580810 129684 580816 129696
rect 580868 129684 580874 129736
rect 126054 124108 126060 124160
rect 126112 124148 126118 124160
rect 126422 124148 126428 124160
rect 126112 124120 126428 124148
rect 126112 124108 126118 124120
rect 126422 124108 126428 124120
rect 126480 124108 126486 124160
rect 131114 124108 131120 124160
rect 131172 124148 131178 124160
rect 131390 124148 131396 124160
rect 131172 124120 131396 124148
rect 131172 124108 131178 124120
rect 131390 124108 131396 124120
rect 131448 124108 131454 124160
rect 134058 122380 134064 122392
rect 134019 122352 134064 122380
rect 134058 122340 134064 122352
rect 134116 122340 134122 122392
rect 134058 120776 134064 120828
rect 134116 120816 134122 120828
rect 580902 120816 580908 120828
rect 134116 120788 580908 120816
rect 134116 120776 134122 120788
rect 580902 120776 580908 120788
rect 580960 120776 580966 120828
rect 132402 120708 132408 120760
rect 132460 120748 132466 120760
rect 580350 120748 580356 120760
rect 132460 120720 580356 120748
rect 132460 120708 132466 120720
rect 580350 120708 580356 120720
rect 580408 120708 580414 120760
rect 133966 120640 133972 120692
rect 134024 120680 134030 120692
rect 580258 120680 580264 120692
rect 134024 120652 580264 120680
rect 134024 120640 134030 120652
rect 580258 120640 580264 120652
rect 580316 120640 580322 120692
rect 3326 120572 3332 120624
rect 3384 120612 3390 120624
rect 138569 120615 138627 120621
rect 138569 120612 138581 120615
rect 3384 120584 138581 120612
rect 3384 120572 3390 120584
rect 138569 120581 138581 120584
rect 138615 120581 138627 120615
rect 138569 120575 138627 120581
rect 143445 120615 143503 120621
rect 143445 120581 143457 120615
rect 143491 120612 143503 120615
rect 436278 120612 436284 120624
rect 143491 120584 436284 120612
rect 143491 120581 143503 120584
rect 143445 120575 143503 120581
rect 436278 120572 436284 120584
rect 436336 120572 436342 120624
rect 143537 120547 143595 120553
rect 143537 120544 143549 120547
rect 143460 120516 143549 120544
rect 134061 120479 134119 120485
rect 134061 120445 134073 120479
rect 134107 120476 134119 120479
rect 143460 120476 143488 120516
rect 143537 120513 143549 120516
rect 143583 120513 143595 120547
rect 143537 120507 143595 120513
rect 134107 120448 143488 120476
rect 161385 120479 161443 120485
rect 134107 120445 134119 120448
rect 134061 120439 134119 120445
rect 161385 120445 161397 120479
rect 161431 120476 161443 120479
rect 171137 120479 171195 120485
rect 171137 120476 171149 120479
rect 161431 120448 171149 120476
rect 161431 120445 161443 120448
rect 161385 120439 161443 120445
rect 171137 120445 171149 120448
rect 171183 120445 171195 120479
rect 171137 120439 171195 120445
rect 180705 120479 180763 120485
rect 180705 120445 180717 120479
rect 180751 120476 180763 120479
rect 182177 120479 182235 120485
rect 182177 120476 182189 120479
rect 180751 120448 182189 120476
rect 180751 120445 180763 120448
rect 180705 120439 180763 120445
rect 182177 120445 182189 120448
rect 182223 120445 182235 120479
rect 182177 120439 182235 120445
rect 138569 120411 138627 120417
rect 138569 120377 138581 120411
rect 138615 120408 138627 120411
rect 143445 120411 143503 120417
rect 143445 120408 143457 120411
rect 138615 120380 143457 120408
rect 138615 120377 138627 120380
rect 138569 120371 138627 120377
rect 143445 120377 143457 120380
rect 143491 120377 143503 120411
rect 143445 120371 143503 120377
rect 133138 120300 133144 120352
rect 133196 120340 133202 120352
rect 135162 120340 135168 120352
rect 133196 120312 135168 120340
rect 133196 120300 133202 120312
rect 135162 120300 135168 120312
rect 135220 120300 135226 120352
rect 143537 120343 143595 120349
rect 143537 120309 143549 120343
rect 143583 120340 143595 120343
rect 151817 120343 151875 120349
rect 151817 120340 151829 120343
rect 143583 120312 151829 120340
rect 143583 120309 143595 120312
rect 143537 120303 143595 120309
rect 151817 120309 151829 120312
rect 151863 120309 151875 120343
rect 151817 120303 151875 120309
rect 171137 120343 171195 120349
rect 171137 120309 171149 120343
rect 171183 120340 171195 120343
rect 180705 120343 180763 120349
rect 180705 120340 180717 120343
rect 171183 120312 180717 120340
rect 171183 120309 171195 120312
rect 171137 120303 171195 120309
rect 180705 120309 180717 120312
rect 180751 120309 180763 120343
rect 180705 120303 180763 120309
rect 182177 120275 182235 120281
rect 182177 120241 182189 120275
rect 182223 120272 182235 120275
rect 186590 120272 186596 120284
rect 182223 120244 186596 120272
rect 182223 120241 182235 120244
rect 182177 120235 182235 120241
rect 186590 120232 186596 120244
rect 186648 120232 186654 120284
rect 151817 120207 151875 120213
rect 151817 120173 151829 120207
rect 151863 120204 151875 120207
rect 161385 120207 161443 120213
rect 161385 120204 161397 120207
rect 151863 120176 161397 120204
rect 151863 120173 151875 120176
rect 151817 120167 151875 120173
rect 161385 120173 161397 120176
rect 161431 120173 161443 120207
rect 161385 120167 161443 120173
rect 145006 120136 145012 120148
rect 144967 120108 145012 120136
rect 145006 120096 145012 120108
rect 145064 120096 145070 120148
rect 395108 119756 395114 119808
rect 395166 119796 395172 119808
rect 395982 119796 395988 119808
rect 395166 119768 395988 119796
rect 395166 119756 395172 119768
rect 395982 119756 395988 119768
rect 396040 119756 396046 119808
rect 135162 119348 135168 119400
rect 135220 119388 135226 119400
rect 192110 119388 192116 119400
rect 135220 119360 192116 119388
rect 135220 119348 135226 119360
rect 192110 119348 192116 119360
rect 192168 119348 192174 119400
rect 138290 119280 138296 119332
rect 138348 119320 138354 119332
rect 138842 119320 138848 119332
rect 138348 119292 138848 119320
rect 138348 119280 138354 119292
rect 138842 119280 138848 119292
rect 138900 119280 138906 119332
rect 130746 118940 130752 118992
rect 130804 118980 130810 118992
rect 140774 118980 140780 118992
rect 130804 118952 140780 118980
rect 130804 118940 130810 118952
rect 140774 118940 140780 118952
rect 140832 118940 140838 118992
rect 130930 118872 130936 118924
rect 130988 118912 130994 118924
rect 142246 118912 142252 118924
rect 130988 118884 142252 118912
rect 130988 118872 130994 118884
rect 142246 118872 142252 118884
rect 142304 118912 142310 118924
rect 142522 118912 142528 118924
rect 142304 118884 142528 118912
rect 142304 118872 142310 118884
rect 142522 118872 142528 118884
rect 142580 118872 142586 118924
rect 129550 118804 129556 118856
rect 129608 118844 129614 118856
rect 145009 118847 145067 118853
rect 145009 118844 145021 118847
rect 129608 118816 145021 118844
rect 129608 118804 129614 118816
rect 145009 118813 145021 118816
rect 145055 118813 145067 118847
rect 145009 118807 145067 118813
rect 131022 118736 131028 118788
rect 131080 118776 131086 118788
rect 149054 118776 149060 118788
rect 131080 118748 149060 118776
rect 131080 118736 131086 118748
rect 149054 118736 149060 118748
rect 149112 118736 149118 118788
rect 129642 118668 129648 118720
rect 129700 118708 129706 118720
rect 147766 118708 147772 118720
rect 129700 118680 147772 118708
rect 129700 118668 129706 118680
rect 147766 118668 147772 118680
rect 147824 118668 147830 118720
rect 424778 118668 424784 118720
rect 424836 118708 424842 118720
rect 424836 118680 425468 118708
rect 424836 118668 424842 118680
rect 42702 118600 42708 118652
rect 42760 118640 42766 118652
rect 129734 118640 129740 118652
rect 42760 118612 129740 118640
rect 42760 118600 42766 118612
rect 129734 118600 129740 118612
rect 129792 118640 129798 118652
rect 155310 118640 155316 118652
rect 129792 118612 155316 118640
rect 129792 118600 129798 118612
rect 155310 118600 155316 118612
rect 155368 118600 155374 118652
rect 210421 118643 210479 118649
rect 210421 118609 210433 118643
rect 210467 118640 210479 118643
rect 218422 118640 218428 118652
rect 210467 118612 218428 118640
rect 210467 118609 210479 118612
rect 210421 118603 210479 118609
rect 218422 118600 218428 118612
rect 218480 118600 218486 118652
rect 220081 118643 220139 118649
rect 220081 118609 220093 118643
rect 220127 118640 220139 118643
rect 243538 118640 243544 118652
rect 220127 118612 243544 118640
rect 220127 118609 220139 118612
rect 220081 118603 220139 118609
rect 243538 118600 243544 118612
rect 243596 118600 243602 118652
rect 243633 118643 243691 118649
rect 243633 118609 243645 118643
rect 243679 118640 243691 118643
rect 253290 118640 253296 118652
rect 243679 118612 253296 118640
rect 243679 118609 243691 118612
rect 243633 118603 243691 118609
rect 253290 118600 253296 118612
rect 253348 118600 253354 118652
rect 253385 118643 253443 118649
rect 253385 118609 253397 118643
rect 253431 118640 253443 118643
rect 258258 118640 258264 118652
rect 253431 118612 258264 118640
rect 253431 118609 253443 118612
rect 253385 118603 253443 118609
rect 258258 118600 258264 118612
rect 258316 118600 258322 118652
rect 306006 118600 306012 118652
rect 306064 118640 306070 118652
rect 332870 118640 332876 118652
rect 306064 118612 332876 118640
rect 306064 118600 306070 118612
rect 332870 118600 332876 118612
rect 332928 118600 332934 118652
rect 353110 118600 353116 118652
rect 353168 118640 353174 118652
rect 425330 118640 425336 118652
rect 353168 118612 425336 118640
rect 353168 118600 353174 118612
rect 425330 118600 425336 118612
rect 425388 118600 425394 118652
rect 425440 118640 425468 118680
rect 426268 118680 429976 118708
rect 426268 118640 426296 118680
rect 425440 118612 426296 118640
rect 426342 118600 426348 118652
rect 426400 118640 426406 118652
rect 429838 118640 429844 118652
rect 426400 118612 429844 118640
rect 426400 118600 426406 118612
rect 429838 118600 429844 118612
rect 429896 118600 429902 118652
rect 429948 118640 429976 118680
rect 431681 118643 431739 118649
rect 431681 118640 431693 118643
rect 429948 118612 431693 118640
rect 431681 118609 431693 118612
rect 431727 118609 431739 118643
rect 431681 118603 431739 118609
rect 431770 118600 431776 118652
rect 431828 118640 431834 118652
rect 511258 118640 511264 118652
rect 431828 118612 511264 118640
rect 431828 118600 431834 118612
rect 511258 118600 511264 118612
rect 511316 118600 511322 118652
rect 97902 118532 97908 118584
rect 97960 118572 97966 118584
rect 181070 118572 181076 118584
rect 97960 118544 181076 118572
rect 97960 118532 97966 118544
rect 181070 118532 181076 118544
rect 181128 118532 181134 118584
rect 190362 118532 190368 118584
rect 190420 118572 190426 118584
rect 231302 118572 231308 118584
rect 190420 118544 231308 118572
rect 190420 118532 190426 118544
rect 231302 118532 231308 118544
rect 231360 118532 231366 118584
rect 237190 118532 237196 118584
rect 237248 118572 237254 118584
rect 255314 118572 255320 118584
rect 237248 118544 255320 118572
rect 237248 118532 237254 118544
rect 255314 118532 255320 118544
rect 255372 118532 255378 118584
rect 257338 118532 257344 118584
rect 257396 118572 257402 118584
rect 264330 118572 264336 118584
rect 257396 118544 264336 118572
rect 257396 118532 257402 118544
rect 264330 118532 264336 118544
rect 264388 118532 264394 118584
rect 308490 118532 308496 118584
rect 308548 118572 308554 118584
rect 338390 118572 338396 118584
rect 308548 118544 338396 118572
rect 308548 118532 308554 118544
rect 338390 118532 338396 118544
rect 338448 118532 338454 118584
rect 362310 118532 362316 118584
rect 362368 118572 362374 118584
rect 442994 118572 443000 118584
rect 362368 118544 443000 118572
rect 362368 118532 362374 118544
rect 442994 118532 443000 118544
rect 443052 118532 443058 118584
rect 82722 118464 82728 118516
rect 82780 118504 82786 118516
rect 164510 118504 164516 118516
rect 82780 118476 164516 118504
rect 82780 118464 82786 118476
rect 164510 118464 164516 118476
rect 164568 118464 164574 118516
rect 175918 118464 175924 118516
rect 175976 118504 175982 118516
rect 210421 118507 210479 118513
rect 210421 118504 210433 118507
rect 175976 118476 210433 118504
rect 175976 118464 175982 118476
rect 210421 118473 210433 118476
rect 210467 118473 210479 118507
rect 210421 118467 210479 118473
rect 210513 118507 210571 118513
rect 210513 118473 210525 118507
rect 210559 118504 210571 118507
rect 220262 118504 220268 118516
rect 210559 118476 220268 118504
rect 210559 118473 210571 118476
rect 210513 118467 210571 118473
rect 220262 118464 220268 118476
rect 220320 118464 220326 118516
rect 220357 118507 220415 118513
rect 220357 118473 220369 118507
rect 220403 118504 220415 118507
rect 227714 118504 227720 118516
rect 220403 118476 227720 118504
rect 220403 118473 220415 118476
rect 220357 118467 220415 118473
rect 227714 118464 227720 118476
rect 227772 118464 227778 118516
rect 232498 118464 232504 118516
rect 232556 118504 232562 118516
rect 240226 118504 240232 118516
rect 232556 118476 240232 118504
rect 232556 118464 232562 118476
rect 240226 118464 240232 118476
rect 240284 118464 240290 118516
rect 240962 118464 240968 118516
rect 241020 118504 241026 118516
rect 247770 118504 247776 118516
rect 241020 118476 247776 118504
rect 241020 118464 241026 118476
rect 247770 118464 247776 118476
rect 247828 118464 247834 118516
rect 249061 118507 249119 118513
rect 249061 118473 249073 118507
rect 249107 118504 249119 118507
rect 253385 118507 253443 118513
rect 253385 118504 253397 118507
rect 249107 118476 253397 118504
rect 249107 118473 249119 118476
rect 249061 118467 249119 118473
rect 253385 118473 253397 118476
rect 253431 118473 253443 118507
rect 253385 118467 253443 118473
rect 310882 118464 310888 118516
rect 310940 118504 310946 118516
rect 341426 118504 341432 118516
rect 310940 118476 341432 118504
rect 310940 118464 310946 118476
rect 341426 118464 341432 118476
rect 341484 118464 341490 118516
rect 347590 118464 347596 118516
rect 347648 118504 347654 118516
rect 376018 118504 376024 118516
rect 347648 118476 376024 118504
rect 347648 118464 347654 118476
rect 376018 118464 376024 118476
rect 376076 118464 376082 118516
rect 393590 118464 393596 118516
rect 393648 118504 393654 118516
rect 475378 118504 475384 118516
rect 393648 118476 475384 118504
rect 393648 118464 393654 118476
rect 475378 118464 475384 118476
rect 475436 118464 475442 118516
rect 71498 118396 71504 118448
rect 71556 118436 71562 118448
rect 88334 118436 88340 118448
rect 71556 118408 88340 118436
rect 71556 118396 71562 118408
rect 88334 118396 88340 118408
rect 88392 118396 88398 118448
rect 124122 118396 124128 118448
rect 124180 118436 124186 118448
rect 190454 118436 190460 118448
rect 124180 118408 190460 118436
rect 124180 118396 124186 118408
rect 190454 118396 190460 118408
rect 190512 118396 190518 118448
rect 194502 118396 194508 118448
rect 194560 118436 194566 118448
rect 233234 118436 233240 118448
rect 194560 118408 233240 118436
rect 194560 118396 194566 118408
rect 233234 118396 233240 118408
rect 233292 118396 233298 118448
rect 234522 118396 234528 118448
rect 234580 118436 234586 118448
rect 253934 118436 253940 118448
rect 234580 118408 253940 118436
rect 234580 118396 234586 118408
rect 253934 118396 253940 118408
rect 253992 118396 253998 118448
rect 256602 118396 256608 118448
rect 256660 118436 256666 118448
rect 265526 118436 265532 118448
rect 256660 118408 265532 118436
rect 256660 118396 256666 118408
rect 265526 118396 265532 118408
rect 265584 118396 265590 118448
rect 309686 118396 309692 118448
rect 309744 118436 309750 118448
rect 339586 118436 339592 118448
rect 309744 118408 339592 118436
rect 309744 118396 309750 118408
rect 339586 118396 339592 118408
rect 339644 118396 339650 118448
rect 342162 118396 342168 118448
rect 342220 118436 342226 118448
rect 389818 118436 389824 118448
rect 342220 118408 389824 118436
rect 342220 118396 342226 118408
rect 389818 118396 389824 118408
rect 389876 118396 389882 118448
rect 397270 118396 397276 118448
rect 397328 118436 397334 118448
rect 478138 118436 478144 118448
rect 397328 118408 478144 118436
rect 397328 118396 397334 118408
rect 478138 118396 478144 118408
rect 478196 118396 478202 118448
rect 56502 118328 56508 118380
rect 56560 118368 56566 118380
rect 125778 118368 125784 118380
rect 56560 118340 125784 118368
rect 56560 118328 56566 118340
rect 125778 118328 125784 118340
rect 125836 118328 125842 118380
rect 129274 118328 129280 118380
rect 129332 118368 129338 118380
rect 182910 118368 182916 118380
rect 129332 118340 182916 118368
rect 129332 118328 129338 118340
rect 182910 118328 182916 118340
rect 182968 118328 182974 118380
rect 186038 118328 186044 118380
rect 186096 118368 186102 118380
rect 229462 118368 229468 118380
rect 186096 118340 229468 118368
rect 186096 118328 186102 118340
rect 229462 118328 229468 118340
rect 229520 118328 229526 118380
rect 231762 118328 231768 118380
rect 231820 118368 231826 118380
rect 252738 118368 252744 118380
rect 231820 118340 252744 118368
rect 231820 118328 231826 118340
rect 252738 118328 252744 118340
rect 252796 118328 252802 118380
rect 257982 118328 257988 118380
rect 258040 118368 258046 118380
rect 266354 118368 266360 118380
rect 258040 118340 266360 118368
rect 258040 118328 258046 118340
rect 266354 118328 266360 118340
rect 266412 118328 266418 118380
rect 311526 118328 311532 118380
rect 311584 118368 311590 118380
rect 343910 118368 343916 118380
rect 311584 118340 343916 118368
rect 311584 118328 311590 118340
rect 343910 118328 343916 118340
rect 343968 118328 343974 118380
rect 365990 118328 365996 118380
rect 366048 118368 366054 118380
rect 449894 118368 449900 118380
rect 366048 118340 449900 118368
rect 366048 118328 366054 118340
rect 449894 118328 449900 118340
rect 449952 118328 449958 118380
rect 31662 118260 31668 118312
rect 31720 118300 31726 118312
rect 107562 118300 107568 118312
rect 31720 118272 107568 118300
rect 31720 118260 31726 118272
rect 107562 118260 107568 118272
rect 107620 118260 107626 118312
rect 109034 118260 109040 118312
rect 109092 118300 109098 118312
rect 109092 118272 111840 118300
rect 109092 118260 109098 118272
rect 28902 118192 28908 118244
rect 28960 118232 28966 118244
rect 111702 118232 111708 118244
rect 28960 118204 111708 118232
rect 28960 118192 28966 118204
rect 111702 118192 111708 118204
rect 111760 118192 111766 118244
rect 23382 118124 23388 118176
rect 23440 118164 23446 118176
rect 110322 118164 110328 118176
rect 23440 118136 110328 118164
rect 23440 118124 23446 118136
rect 110322 118124 110328 118136
rect 110380 118124 110386 118176
rect 111812 118164 111840 118272
rect 113082 118260 113088 118312
rect 113140 118300 113146 118312
rect 175642 118300 175648 118312
rect 113140 118272 175648 118300
rect 113140 118260 113146 118272
rect 175642 118260 175648 118272
rect 175700 118260 175706 118312
rect 176010 118260 176016 118312
rect 176068 118300 176074 118312
rect 210513 118303 210571 118309
rect 210513 118300 210525 118303
rect 176068 118272 210525 118300
rect 176068 118260 176074 118272
rect 210513 118269 210525 118272
rect 210559 118269 210571 118303
rect 210513 118263 210571 118269
rect 213822 118260 213828 118312
rect 213880 118300 213886 118312
rect 220081 118303 220139 118309
rect 220081 118300 220093 118303
rect 213880 118272 220093 118300
rect 213880 118260 213886 118272
rect 220081 118269 220093 118272
rect 220127 118269 220139 118303
rect 220081 118263 220139 118269
rect 220265 118303 220323 118309
rect 220265 118269 220277 118303
rect 220311 118300 220323 118303
rect 223666 118300 223672 118312
rect 220311 118272 223672 118300
rect 220311 118269 220323 118272
rect 220265 118263 220323 118269
rect 223666 118260 223672 118272
rect 223724 118260 223730 118312
rect 227622 118260 227628 118312
rect 227680 118300 227686 118312
rect 250254 118300 250260 118312
rect 227680 118272 250260 118300
rect 227680 118260 227686 118272
rect 250254 118260 250260 118272
rect 250312 118260 250318 118312
rect 250530 118260 250536 118312
rect 250588 118300 250594 118312
rect 260834 118300 260840 118312
rect 250588 118272 260840 118300
rect 250588 118260 250594 118272
rect 260834 118260 260840 118272
rect 260892 118260 260898 118312
rect 296162 118260 296168 118312
rect 296220 118300 296226 118312
rect 305638 118300 305644 118312
rect 296220 118272 305644 118300
rect 296220 118260 296226 118272
rect 305638 118260 305644 118272
rect 305696 118260 305702 118312
rect 307202 118260 307208 118312
rect 307260 118300 307266 118312
rect 334618 118300 334624 118312
rect 307260 118272 334624 118300
rect 307260 118260 307266 118272
rect 334618 118260 334624 118272
rect 334676 118260 334682 118312
rect 336642 118260 336648 118312
rect 336700 118300 336706 118312
rect 374638 118300 374644 118312
rect 336700 118272 374644 118300
rect 336700 118260 336706 118272
rect 374638 118260 374644 118272
rect 374696 118260 374702 118312
rect 377030 118260 377036 118312
rect 377088 118300 377094 118312
rect 384301 118303 384359 118309
rect 384301 118300 384313 118303
rect 377088 118272 384313 118300
rect 377088 118260 377094 118272
rect 384301 118269 384313 118272
rect 384347 118269 384359 118303
rect 384301 118263 384359 118269
rect 389910 118260 389916 118312
rect 389968 118300 389974 118312
rect 473998 118300 474004 118312
rect 389968 118272 474004 118300
rect 389968 118260 389974 118272
rect 473998 118260 474004 118272
rect 474056 118260 474062 118312
rect 129182 118192 129188 118244
rect 129240 118232 129246 118244
rect 177390 118232 177396 118244
rect 129240 118204 177396 118232
rect 129240 118192 129246 118204
rect 177390 118192 177396 118204
rect 177448 118192 177454 118244
rect 179322 118192 179328 118244
rect 179380 118232 179386 118244
rect 219986 118232 219992 118244
rect 179380 118204 219992 118232
rect 179380 118192 179386 118204
rect 219986 118192 219992 118204
rect 220044 118192 220050 118244
rect 220173 118235 220231 118241
rect 220173 118201 220185 118235
rect 220219 118232 220231 118235
rect 222194 118232 222200 118244
rect 220219 118204 222200 118232
rect 220219 118201 220231 118204
rect 220173 118195 220231 118201
rect 222194 118192 222200 118204
rect 222252 118192 222258 118244
rect 231118 118192 231124 118244
rect 231176 118232 231182 118244
rect 238018 118232 238024 118244
rect 231176 118204 238024 118232
rect 231176 118192 231182 118204
rect 238018 118192 238024 118204
rect 238076 118192 238082 118244
rect 238113 118235 238171 118241
rect 238113 118201 238125 118235
rect 238159 118232 238171 118235
rect 252094 118232 252100 118244
rect 238159 118204 252100 118232
rect 238159 118201 238171 118204
rect 238113 118195 238171 118201
rect 252094 118192 252100 118204
rect 252152 118192 252158 118244
rect 254670 118192 254676 118244
rect 254728 118232 254734 118244
rect 263686 118232 263692 118244
rect 254728 118204 263692 118232
rect 254728 118192 254734 118204
rect 263686 118192 263692 118204
rect 263744 118192 263750 118244
rect 293770 118192 293776 118244
rect 293828 118232 293834 118244
rect 302878 118232 302884 118244
rect 293828 118204 302884 118232
rect 293828 118192 293834 118204
rect 302878 118192 302884 118204
rect 302936 118192 302942 118244
rect 307662 118192 307668 118244
rect 307720 118232 307726 118244
rect 336918 118232 336924 118244
rect 307720 118204 336924 118232
rect 307720 118192 307726 118204
rect 336918 118192 336924 118204
rect 336976 118192 336982 118244
rect 338482 118192 338488 118244
rect 338540 118232 338546 118244
rect 384206 118232 384212 118244
rect 338540 118204 384212 118232
rect 338540 118192 338546 118204
rect 384206 118192 384212 118204
rect 384264 118192 384270 118244
rect 386230 118192 386236 118244
rect 386288 118232 386294 118244
rect 469858 118232 469864 118244
rect 386288 118204 469864 118232
rect 386288 118192 386294 118204
rect 469858 118192 469864 118204
rect 469916 118192 469922 118244
rect 123849 118167 123907 118173
rect 123849 118164 123861 118167
rect 111812 118136 123861 118164
rect 123849 118133 123861 118136
rect 123895 118133 123907 118167
rect 123849 118127 123907 118133
rect 129090 118124 129096 118176
rect 129148 118164 129154 118176
rect 173894 118164 173900 118176
rect 129148 118136 173900 118164
rect 129148 118124 129154 118136
rect 173894 118124 173900 118136
rect 173952 118124 173958 118176
rect 177298 118124 177304 118176
rect 177356 118164 177362 118176
rect 223942 118164 223948 118176
rect 177356 118136 223948 118164
rect 177356 118124 177362 118136
rect 223942 118124 223948 118136
rect 224000 118124 224006 118176
rect 226242 118124 226248 118176
rect 226300 118164 226306 118176
rect 249794 118164 249800 118176
rect 226300 118136 249800 118164
rect 226300 118124 226306 118136
rect 249794 118124 249800 118136
rect 249852 118124 249858 118176
rect 251082 118124 251088 118176
rect 251140 118164 251146 118176
rect 262490 118164 262496 118176
rect 251140 118136 262496 118164
rect 251140 118124 251146 118136
rect 262490 118124 262496 118136
rect 262548 118124 262554 118176
rect 283926 118124 283932 118176
rect 283984 118164 283990 118176
rect 290090 118164 290096 118176
rect 283984 118136 290096 118164
rect 283984 118124 283990 118136
rect 290090 118124 290096 118136
rect 290148 118124 290154 118176
rect 295610 118124 295616 118176
rect 295668 118164 295674 118176
rect 308398 118164 308404 118176
rect 295668 118136 308404 118164
rect 295668 118124 295674 118136
rect 308398 118124 308404 118136
rect 308456 118124 308462 118176
rect 311710 118124 311716 118176
rect 311768 118164 311774 118176
rect 345198 118164 345204 118176
rect 311768 118136 345204 118164
rect 311768 118124 311774 118136
rect 345198 118124 345204 118136
rect 345256 118124 345262 118176
rect 349430 118124 349436 118176
rect 349488 118164 349494 118176
rect 359461 118167 359519 118173
rect 359461 118164 359473 118167
rect 349488 118136 359473 118164
rect 349488 118124 349494 118136
rect 359461 118133 359473 118136
rect 359507 118133 359519 118167
rect 359461 118127 359519 118133
rect 369670 118124 369676 118176
rect 369728 118164 369734 118176
rect 456794 118164 456800 118176
rect 369728 118136 456800 118164
rect 369728 118124 369734 118136
rect 456794 118124 456800 118136
rect 456852 118124 456858 118176
rect 71682 118056 71688 118108
rect 71740 118096 71746 118108
rect 73798 118096 73804 118108
rect 71740 118068 73804 118096
rect 71740 118056 71746 118068
rect 73798 118056 73804 118068
rect 73856 118096 73862 118108
rect 73982 118096 73988 118108
rect 73856 118068 73988 118096
rect 73856 118056 73862 118068
rect 73982 118056 73988 118068
rect 74040 118056 74046 118108
rect 125686 118056 125692 118108
rect 125744 118096 125750 118108
rect 170030 118096 170036 118108
rect 125744 118068 170036 118096
rect 125744 118056 125750 118068
rect 170030 118056 170036 118068
rect 170088 118056 170094 118108
rect 170398 118056 170404 118108
rect 170456 118096 170462 118108
rect 216674 118096 216680 118108
rect 170456 118068 216680 118096
rect 170456 118056 170462 118068
rect 216674 118056 216680 118068
rect 216732 118056 216738 118108
rect 219250 118056 219256 118108
rect 219308 118096 219314 118108
rect 245930 118096 245936 118108
rect 219308 118068 245936 118096
rect 219308 118056 219314 118068
rect 245930 118056 245936 118068
rect 245988 118056 245994 118108
rect 248322 118056 248328 118108
rect 248380 118096 248386 118108
rect 261294 118096 261300 118108
rect 248380 118068 261300 118096
rect 248380 118056 248386 118068
rect 261294 118056 261300 118068
rect 261352 118056 261358 118108
rect 264974 118096 264980 118108
rect 261680 118068 264980 118096
rect 60642 117988 60648 118040
rect 60700 118028 60706 118040
rect 82722 118028 82728 118040
rect 60700 118000 82728 118028
rect 60700 117988 60706 118000
rect 82722 117988 82728 118000
rect 82780 117988 82786 118040
rect 88334 117988 88340 118040
rect 88392 118028 88398 118040
rect 115937 118031 115995 118037
rect 115937 118028 115949 118031
rect 88392 118000 115949 118028
rect 88392 117988 88398 118000
rect 115937 117997 115949 118000
rect 115983 117997 115995 118031
rect 115937 117991 115995 117997
rect 123757 118031 123815 118037
rect 123757 117997 123769 118031
rect 123803 118028 123815 118031
rect 179414 118028 179420 118040
rect 123803 118000 179420 118028
rect 123803 117997 123815 118000
rect 123757 117991 123815 117997
rect 179414 117988 179420 118000
rect 179472 117988 179478 118040
rect 183462 117988 183468 118040
rect 183520 118028 183526 118040
rect 183520 118000 220032 118028
rect 183520 117988 183526 118000
rect 38470 117920 38476 117972
rect 38528 117960 38534 117972
rect 69658 117960 69664 117972
rect 38528 117932 69664 117960
rect 38528 117920 38534 117932
rect 69658 117920 69664 117932
rect 69716 117920 69722 117972
rect 73982 117920 73988 117972
rect 74040 117960 74046 117972
rect 89717 117963 89775 117969
rect 89717 117960 89729 117963
rect 74040 117932 89729 117960
rect 74040 117920 74046 117932
rect 89717 117929 89729 117932
rect 89763 117929 89775 117963
rect 89717 117923 89775 117929
rect 108945 117963 109003 117969
rect 108945 117929 108957 117963
rect 108991 117960 109003 117963
rect 109034 117960 109040 117972
rect 108991 117932 109040 117960
rect 108991 117929 109003 117932
rect 108945 117923 109003 117929
rect 109034 117920 109040 117932
rect 109092 117920 109098 117972
rect 123849 117963 123907 117969
rect 123849 117929 123861 117963
rect 123895 117960 123907 117963
rect 137925 117963 137983 117969
rect 137925 117960 137937 117963
rect 123895 117932 137937 117960
rect 123895 117929 123907 117932
rect 123849 117923 123907 117929
rect 137925 117929 137937 117932
rect 137971 117929 137983 117963
rect 137925 117923 137983 117929
rect 138017 117963 138075 117969
rect 138017 117929 138029 117963
rect 138063 117960 138075 117963
rect 147677 117963 147735 117969
rect 147677 117960 147689 117963
rect 138063 117932 147689 117960
rect 138063 117929 138075 117932
rect 138017 117923 138075 117929
rect 147677 117929 147689 117932
rect 147723 117929 147735 117963
rect 147677 117923 147735 117929
rect 164145 117963 164203 117969
rect 164145 117929 164157 117963
rect 164191 117960 164203 117963
rect 171870 117960 171876 117972
rect 164191 117932 171876 117960
rect 164191 117929 164203 117932
rect 164145 117923 164203 117929
rect 171870 117920 171876 117932
rect 171928 117920 171934 117972
rect 174538 117920 174544 117972
rect 174596 117960 174602 117972
rect 219897 117963 219955 117969
rect 219897 117960 219909 117963
rect 174596 117932 219909 117960
rect 174596 117920 174602 117932
rect 219897 117929 219909 117932
rect 219943 117929 219955 117963
rect 220004 117960 220032 118000
rect 220078 117988 220084 118040
rect 220136 118028 220142 118040
rect 225782 118028 225788 118040
rect 220136 118000 225788 118028
rect 220136 117988 220142 118000
rect 225782 117988 225788 118000
rect 225840 117988 225846 118040
rect 229002 117988 229008 118040
rect 229060 118028 229066 118040
rect 251266 118028 251272 118040
rect 229060 118000 251272 118028
rect 229060 117988 229066 118000
rect 251266 117988 251272 118000
rect 251324 117988 251330 118040
rect 255222 117988 255228 118040
rect 255280 118028 255286 118040
rect 261680 118028 261708 118068
rect 264974 118056 264980 118068
rect 265032 118056 265038 118108
rect 284570 118056 284576 118108
rect 284628 118096 284634 118108
rect 291378 118096 291384 118108
rect 284628 118068 291384 118096
rect 284628 118056 284634 118068
rect 291378 118056 291384 118068
rect 291436 118056 291442 118108
rect 296622 118056 296628 118108
rect 296680 118096 296686 118108
rect 314838 118096 314844 118108
rect 296680 118068 314844 118096
rect 296680 118056 296686 118068
rect 314838 118056 314844 118068
rect 314896 118056 314902 118108
rect 324869 118099 324927 118105
rect 324869 118065 324881 118099
rect 324915 118096 324927 118099
rect 357986 118096 357992 118108
rect 324915 118068 357992 118096
rect 324915 118065 324927 118068
rect 324869 118059 324927 118065
rect 357986 118056 357992 118068
rect 358044 118056 358050 118108
rect 373350 118056 373356 118108
rect 373408 118096 373414 118108
rect 463694 118096 463700 118108
rect 373408 118068 463700 118096
rect 373408 118056 373414 118068
rect 463694 118056 463700 118068
rect 463752 118056 463758 118108
rect 255280 118000 261708 118028
rect 255280 117988 255286 118000
rect 262122 117988 262128 118040
rect 262180 118028 262186 118040
rect 268010 118028 268016 118040
rect 262180 118000 268016 118028
rect 262180 117988 262186 118000
rect 268010 117988 268016 118000
rect 268068 117988 268074 118040
rect 298646 117988 298652 118040
rect 298704 118028 298710 118040
rect 318978 118028 318984 118040
rect 298704 118000 318984 118028
rect 298704 117988 298710 118000
rect 318978 117988 318984 118000
rect 319036 117988 319042 118040
rect 321922 117988 321928 118040
rect 321980 118028 321986 118040
rect 363506 118028 363512 118040
rect 321980 118000 363512 118028
rect 321980 117988 321986 118000
rect 363506 117988 363512 118000
rect 363564 117988 363570 118040
rect 384301 118031 384359 118037
rect 384301 117997 384313 118031
rect 384347 118028 384359 118031
rect 470594 118028 470600 118040
rect 384347 118000 470600 118028
rect 384347 117997 384359 118000
rect 384301 117991 384359 117997
rect 470594 117988 470600 118000
rect 470652 117988 470658 118040
rect 220357 117963 220415 117969
rect 220357 117960 220369 117963
rect 220004 117932 220369 117960
rect 219897 117923 219955 117929
rect 220357 117929 220369 117932
rect 220403 117929 220415 117963
rect 220357 117923 220415 117929
rect 223482 117920 223488 117972
rect 223540 117960 223546 117972
rect 248506 117960 248512 117972
rect 223540 117932 248512 117960
rect 223540 117920 223546 117932
rect 248506 117920 248512 117932
rect 248564 117920 248570 117972
rect 249702 117920 249708 117972
rect 249760 117960 249766 117972
rect 262214 117960 262220 117972
rect 249760 117932 262220 117960
rect 249760 117920 249766 117932
rect 262214 117920 262220 117932
rect 262272 117920 262278 117972
rect 263502 117920 263508 117972
rect 263560 117960 263566 117972
rect 268654 117960 268660 117972
rect 263560 117932 268660 117960
rect 263560 117920 263566 117932
rect 268654 117920 268660 117932
rect 268712 117920 268718 117972
rect 294322 117920 294328 117972
rect 294380 117960 294386 117972
rect 295242 117960 295248 117972
rect 294380 117932 295248 117960
rect 294380 117920 294386 117932
rect 295242 117920 295248 117932
rect 295300 117920 295306 117972
rect 297450 117920 297456 117972
rect 297508 117960 297514 117972
rect 298002 117960 298008 117972
rect 297508 117932 298008 117960
rect 297508 117920 297514 117932
rect 298002 117920 298008 117932
rect 298060 117920 298066 117972
rect 300486 117920 300492 117972
rect 300544 117960 300550 117972
rect 321738 117960 321744 117972
rect 300544 117932 321744 117960
rect 300544 117920 300550 117932
rect 321738 117920 321744 117932
rect 321796 117920 321802 117972
rect 325418 117920 325424 117972
rect 325476 117960 325482 117972
rect 369118 117960 369124 117972
rect 325476 117932 369124 117960
rect 325476 117920 325482 117932
rect 369118 117920 369124 117932
rect 369176 117920 369182 117972
rect 380710 117920 380716 117972
rect 380768 117960 380774 117972
rect 477494 117960 477500 117972
rect 380768 117932 477500 117960
rect 380768 117920 380774 117932
rect 477494 117920 477500 117932
rect 477552 117920 477558 117972
rect 99190 117852 99196 117904
rect 99248 117892 99254 117904
rect 101214 117892 101220 117904
rect 99248 117864 101220 117892
rect 99248 117852 99254 117864
rect 101214 117852 101220 117864
rect 101272 117852 101278 117904
rect 107562 117852 107568 117904
rect 107620 117892 107626 117904
rect 149882 117892 149888 117904
rect 107620 117864 149888 117892
rect 107620 117852 107626 117864
rect 149882 117852 149888 117864
rect 149940 117852 149946 117904
rect 150437 117895 150495 117901
rect 150437 117861 150449 117895
rect 150483 117892 150495 117895
rect 154577 117895 154635 117901
rect 154577 117892 154589 117895
rect 150483 117864 154589 117892
rect 150483 117861 150495 117864
rect 150437 117855 150495 117861
rect 154577 117861 154589 117864
rect 154623 117861 154635 117895
rect 154577 117855 154635 117861
rect 185670 117852 185676 117904
rect 185728 117892 185734 117904
rect 225138 117892 225144 117904
rect 185728 117864 225144 117892
rect 185728 117852 185734 117864
rect 225138 117852 225144 117864
rect 225196 117852 225202 117904
rect 226245 117895 226303 117901
rect 226245 117861 226257 117895
rect 226291 117892 226303 117895
rect 229186 117892 229192 117904
rect 226291 117864 229192 117892
rect 226291 117861 226303 117864
rect 226245 117855 226303 117861
rect 229186 117852 229192 117864
rect 229244 117852 229250 117904
rect 229281 117895 229339 117901
rect 229281 117861 229293 117895
rect 229327 117892 229339 117895
rect 236178 117892 236184 117904
rect 229327 117864 236184 117892
rect 229327 117861 229339 117864
rect 229281 117855 229339 117861
rect 236178 117852 236184 117864
rect 236236 117852 236242 117904
rect 237282 117852 237288 117904
rect 237340 117892 237346 117904
rect 255774 117892 255780 117904
rect 237340 117864 255780 117892
rect 237340 117852 237346 117864
rect 255774 117852 255780 117864
rect 255832 117852 255838 117904
rect 263410 117852 263416 117904
rect 263468 117892 263474 117904
rect 269206 117892 269212 117904
rect 263468 117864 269212 117892
rect 263468 117852 263474 117864
rect 269206 117852 269212 117864
rect 269264 117852 269270 117904
rect 288894 117852 288900 117904
rect 288952 117892 288958 117904
rect 288952 117864 293080 117892
rect 288952 117852 288958 117864
rect 82722 117784 82728 117836
rect 82780 117824 82786 117836
rect 113082 117824 113088 117836
rect 82780 117796 113088 117824
rect 82780 117784 82786 117796
rect 113082 117784 113088 117796
rect 113140 117784 113146 117836
rect 122742 117784 122748 117836
rect 122800 117824 122806 117836
rect 160830 117824 160836 117836
rect 122800 117796 160836 117824
rect 122800 117784 122806 117796
rect 160830 117784 160836 117796
rect 160888 117784 160894 117836
rect 200393 117827 200451 117833
rect 200393 117793 200405 117827
rect 200439 117824 200451 117827
rect 234706 117824 234712 117836
rect 200439 117796 234712 117824
rect 200439 117793 200451 117796
rect 200393 117787 200451 117793
rect 234706 117784 234712 117796
rect 234764 117784 234770 117836
rect 238662 117784 238668 117836
rect 238720 117824 238726 117836
rect 256694 117824 256700 117836
rect 238720 117796 256700 117824
rect 238720 117784 238726 117796
rect 256694 117784 256700 117796
rect 256752 117784 256758 117836
rect 293052 117824 293080 117864
rect 293126 117852 293132 117904
rect 293184 117892 293190 117904
rect 293862 117892 293868 117904
rect 293184 117864 293868 117892
rect 293184 117852 293190 117864
rect 293862 117852 293868 117864
rect 293920 117852 293926 117904
rect 304810 117852 304816 117904
rect 304868 117892 304874 117904
rect 331306 117892 331312 117904
rect 304868 117864 331312 117892
rect 304868 117852 304874 117864
rect 331306 117852 331312 117864
rect 331364 117852 331370 117904
rect 359461 117895 359519 117901
rect 359461 117861 359473 117895
rect 359507 117892 359519 117895
rect 416774 117892 416780 117904
rect 359507 117864 416780 117892
rect 359507 117861 359519 117864
rect 359461 117855 359519 117861
rect 416774 117852 416780 117864
rect 416832 117852 416838 117904
rect 416869 117895 416927 117901
rect 416869 117861 416881 117895
rect 416915 117892 416927 117895
rect 420733 117895 420791 117901
rect 420733 117892 420745 117895
rect 416915 117864 420745 117892
rect 416915 117861 416927 117864
rect 416869 117855 416927 117861
rect 420733 117861 420745 117864
rect 420779 117861 420791 117895
rect 420733 117855 420791 117861
rect 420822 117852 420828 117904
rect 420880 117892 420886 117904
rect 500218 117892 500224 117904
rect 420880 117864 500224 117892
rect 420880 117852 420886 117864
rect 500218 117852 500224 117864
rect 500276 117852 500282 117904
rect 297358 117824 297364 117836
rect 293052 117796 297364 117824
rect 297358 117784 297364 117796
rect 297416 117784 297422 117836
rect 306650 117784 306656 117836
rect 306708 117824 306714 117836
rect 333974 117824 333980 117836
rect 306708 117796 333980 117824
rect 306708 117784 306714 117796
rect 333974 117784 333980 117796
rect 334032 117784 334038 117836
rect 344002 117784 344008 117836
rect 344060 117824 344066 117836
rect 344922 117824 344928 117836
rect 344060 117796 344928 117824
rect 344060 117784 344066 117796
rect 344922 117784 344928 117796
rect 344980 117784 344986 117836
rect 345842 117784 345848 117836
rect 345900 117824 345906 117836
rect 396718 117824 396724 117836
rect 345900 117796 396724 117824
rect 345900 117784 345906 117796
rect 396718 117784 396724 117796
rect 396776 117784 396782 117836
rect 422297 117827 422355 117833
rect 422297 117793 422309 117827
rect 422343 117824 422355 117827
rect 423033 117827 423091 117833
rect 423033 117824 423045 117827
rect 422343 117796 423045 117824
rect 422343 117793 422355 117796
rect 422297 117787 422355 117793
rect 423033 117793 423045 117796
rect 423079 117793 423091 117827
rect 423033 117787 423091 117793
rect 427725 117827 427783 117833
rect 427725 117793 427737 117827
rect 427771 117824 427783 117827
rect 480898 117824 480904 117836
rect 427771 117796 480904 117824
rect 427771 117793 427783 117796
rect 427725 117787 427783 117793
rect 480898 117784 480904 117796
rect 480956 117784 480962 117836
rect 89717 117759 89775 117765
rect 89717 117725 89729 117759
rect 89763 117756 89775 117759
rect 108945 117759 109003 117765
rect 108945 117756 108957 117759
rect 89763 117728 108957 117756
rect 89763 117725 89775 117728
rect 89717 117719 89775 117725
rect 108945 117725 108957 117728
rect 108991 117725 109003 117759
rect 108945 117719 109003 117725
rect 115937 117759 115995 117765
rect 115937 117725 115949 117759
rect 115983 117756 115995 117759
rect 123757 117759 123815 117765
rect 123757 117756 123769 117759
rect 115983 117728 123769 117756
rect 115983 117725 115995 117728
rect 115937 117719 115995 117725
rect 123757 117725 123769 117728
rect 123803 117725 123815 117759
rect 123757 117719 123815 117725
rect 125778 117716 125784 117768
rect 125836 117756 125842 117768
rect 162854 117756 162860 117768
rect 125836 117728 162860 117756
rect 125836 117716 125842 117728
rect 162854 117716 162860 117728
rect 162912 117716 162918 117768
rect 185578 117716 185584 117768
rect 185636 117756 185642 117768
rect 219989 117759 220047 117765
rect 219989 117756 220001 117759
rect 185636 117728 220001 117756
rect 185636 117716 185642 117728
rect 219989 117725 220001 117728
rect 220035 117725 220047 117759
rect 219989 117719 220047 117725
rect 220081 117759 220139 117765
rect 220081 117725 220093 117759
rect 220127 117756 220139 117759
rect 229833 117759 229891 117765
rect 229833 117756 229845 117759
rect 220127 117728 229845 117756
rect 220127 117725 220139 117728
rect 220081 117719 220139 117725
rect 229833 117725 229845 117728
rect 229879 117725 229891 117759
rect 229833 117719 229891 117725
rect 233878 117716 233884 117768
rect 233936 117756 233942 117768
rect 238846 117756 238852 117768
rect 233936 117728 238852 117756
rect 233936 117716 233942 117728
rect 238846 117716 238852 117728
rect 238904 117716 238910 117768
rect 243633 117759 243691 117765
rect 243633 117756 243645 117759
rect 239968 117728 243645 117756
rect 104986 117648 104992 117700
rect 105044 117688 105050 117700
rect 115198 117688 115204 117700
rect 105044 117660 115204 117688
rect 105044 117648 105050 117660
rect 115198 117648 115204 117660
rect 115256 117648 115262 117700
rect 129366 117648 129372 117700
rect 129424 117688 129430 117700
rect 135254 117688 135260 117700
rect 129424 117660 135260 117688
rect 129424 117648 129430 117660
rect 135254 117648 135260 117660
rect 135312 117648 135318 117700
rect 135349 117691 135407 117697
rect 135349 117657 135361 117691
rect 135395 117688 135407 117691
rect 166350 117688 166356 117700
rect 135395 117660 166356 117688
rect 135395 117657 135407 117660
rect 135349 117651 135407 117657
rect 166350 117648 166356 117660
rect 166408 117648 166414 117700
rect 175274 117648 175280 117700
rect 175332 117688 175338 117700
rect 175458 117688 175464 117700
rect 175332 117660 175464 117688
rect 175332 117648 175338 117660
rect 175458 117648 175464 117660
rect 175516 117688 175522 117700
rect 195974 117688 195980 117700
rect 175516 117660 195980 117688
rect 175516 117648 175522 117660
rect 195974 117648 195980 117660
rect 196032 117648 196038 117700
rect 197262 117648 197268 117700
rect 197320 117688 197326 117700
rect 197320 117660 226380 117688
rect 197320 117648 197326 117660
rect 128814 117580 128820 117632
rect 128872 117620 128878 117632
rect 130749 117623 130807 117629
rect 130749 117620 130761 117623
rect 128872 117592 130761 117620
rect 128872 117580 128878 117592
rect 130749 117589 130761 117592
rect 130795 117589 130807 117623
rect 158990 117620 158996 117632
rect 130749 117583 130807 117589
rect 130856 117592 158996 117620
rect 130856 117564 130884 117592
rect 158990 117580 158996 117592
rect 159048 117580 159054 117632
rect 195882 117580 195888 117632
rect 195940 117620 195946 117632
rect 200393 117623 200451 117629
rect 200393 117620 200405 117623
rect 195940 117592 200405 117620
rect 195940 117580 195946 117592
rect 200393 117589 200405 117592
rect 200439 117589 200451 117623
rect 226245 117623 226303 117629
rect 226245 117620 226257 117623
rect 200393 117583 200451 117589
rect 200500 117592 226257 117620
rect 120718 117512 120724 117564
rect 120776 117552 120782 117564
rect 125686 117552 125692 117564
rect 120776 117524 125692 117552
rect 120776 117512 120782 117524
rect 125686 117512 125692 117524
rect 125744 117512 125750 117564
rect 130378 117512 130384 117564
rect 130436 117552 130442 117564
rect 130838 117552 130844 117564
rect 130436 117524 130844 117552
rect 130436 117512 130442 117524
rect 130838 117512 130844 117524
rect 130896 117512 130902 117564
rect 130933 117555 130991 117561
rect 130933 117521 130945 117555
rect 130979 117552 130991 117555
rect 135165 117555 135223 117561
rect 135165 117552 135177 117555
rect 130979 117524 135177 117552
rect 130979 117521 130991 117524
rect 130933 117515 130991 117521
rect 135165 117521 135177 117524
rect 135211 117521 135223 117555
rect 135165 117515 135223 117521
rect 135254 117512 135260 117564
rect 135312 117552 135318 117564
rect 135438 117552 135444 117564
rect 135312 117524 135444 117552
rect 135312 117512 135318 117524
rect 135438 117512 135444 117524
rect 135496 117552 135502 117564
rect 142982 117552 142988 117564
rect 135496 117524 142988 117552
rect 135496 117512 135502 117524
rect 142982 117512 142988 117524
rect 143040 117512 143046 117564
rect 143718 117552 143724 117564
rect 143092 117524 143724 117552
rect 122098 117444 122104 117496
rect 122156 117484 122162 117496
rect 122742 117484 122748 117496
rect 122156 117456 122748 117484
rect 122156 117444 122162 117456
rect 122742 117444 122748 117456
rect 122800 117444 122806 117496
rect 123478 117444 123484 117496
rect 123536 117484 123542 117496
rect 124122 117484 124128 117496
rect 123536 117456 124128 117484
rect 123536 117444 123542 117456
rect 124122 117444 124128 117456
rect 124180 117444 124186 117496
rect 130562 117444 130568 117496
rect 130620 117484 130626 117496
rect 143092 117484 143120 117524
rect 143718 117512 143724 117524
rect 143776 117552 143782 117564
rect 157334 117552 157340 117564
rect 143776 117524 157340 117552
rect 143776 117512 143782 117524
rect 157334 117512 157340 117524
rect 157392 117512 157398 117564
rect 193858 117512 193864 117564
rect 193916 117552 193922 117564
rect 200500 117552 200528 117592
rect 226245 117589 226257 117592
rect 226291 117589 226303 117623
rect 226352 117620 226380 117660
rect 233142 117648 233148 117700
rect 233200 117688 233206 117700
rect 239968 117688 239996 117728
rect 243633 117725 243645 117728
rect 243679 117725 243691 117759
rect 243633 117719 243691 117725
rect 245470 117716 245476 117768
rect 245528 117756 245534 117768
rect 259454 117756 259460 117768
rect 245528 117728 259460 117756
rect 245528 117716 245534 117728
rect 259454 117716 259460 117728
rect 259512 117716 259518 117768
rect 302142 117716 302148 117768
rect 302200 117756 302206 117768
rect 325697 117759 325755 117765
rect 325697 117756 325709 117759
rect 302200 117728 325709 117756
rect 302200 117716 302206 117728
rect 325697 117725 325709 117728
rect 325743 117725 325755 117759
rect 325697 117719 325755 117725
rect 329282 117716 329288 117768
rect 329340 117756 329346 117768
rect 358170 117756 358176 117768
rect 329340 117728 358176 117756
rect 329340 117716 329346 117728
rect 358170 117716 358176 117728
rect 358228 117716 358234 117768
rect 364058 117716 364064 117768
rect 364116 117756 364122 117768
rect 391201 117759 391259 117765
rect 391201 117756 391213 117759
rect 364116 117728 391213 117756
rect 364116 117716 364122 117728
rect 391201 117725 391213 117728
rect 391247 117725 391259 117759
rect 391201 117719 391259 117725
rect 400858 117716 400864 117768
rect 400916 117756 400922 117768
rect 413189 117759 413247 117765
rect 413189 117756 413201 117759
rect 400916 117728 413201 117756
rect 400916 117716 400922 117728
rect 413189 117725 413201 117728
rect 413235 117725 413247 117759
rect 413189 117719 413247 117725
rect 415302 117716 415308 117768
rect 415360 117756 415366 117768
rect 418154 117756 418160 117768
rect 415360 117728 418160 117756
rect 415360 117716 415366 117728
rect 418154 117716 418160 117728
rect 418212 117716 418218 117768
rect 429654 117716 429660 117768
rect 429712 117756 429718 117768
rect 430482 117756 430488 117768
rect 429712 117728 430488 117756
rect 429712 117716 429718 117728
rect 430482 117716 430488 117728
rect 430540 117716 430546 117768
rect 430942 117716 430948 117768
rect 431000 117756 431006 117768
rect 431862 117756 431868 117768
rect 431000 117728 431868 117756
rect 431000 117716 431006 117728
rect 431862 117716 431868 117728
rect 431920 117716 431926 117768
rect 431957 117759 432015 117765
rect 431957 117725 431969 117759
rect 432003 117756 432015 117759
rect 502978 117756 502984 117768
rect 432003 117728 502984 117756
rect 432003 117725 432015 117728
rect 431957 117719 432015 117725
rect 502978 117716 502984 117728
rect 503036 117716 503042 117768
rect 233200 117660 239996 117688
rect 233200 117648 233206 117660
rect 240042 117648 240048 117700
rect 240100 117688 240106 117700
rect 256970 117688 256976 117700
rect 240100 117660 256976 117688
rect 240100 117648 240106 117660
rect 256970 117648 256976 117660
rect 257028 117648 257034 117700
rect 261478 117648 261484 117700
rect 261536 117688 261542 117700
rect 267734 117688 267740 117700
rect 261536 117660 267740 117688
rect 261536 117648 261542 117660
rect 267734 117648 267740 117660
rect 267792 117648 267798 117700
rect 304166 117648 304172 117700
rect 304224 117688 304230 117700
rect 329834 117688 329840 117700
rect 304224 117660 329840 117688
rect 304224 117648 304230 117660
rect 329834 117648 329840 117660
rect 329892 117648 329898 117700
rect 360470 117648 360476 117700
rect 360528 117688 360534 117700
rect 398098 117688 398104 117700
rect 360528 117660 398104 117688
rect 360528 117648 360534 117660
rect 398098 117648 398104 117660
rect 398156 117648 398162 117700
rect 411898 117648 411904 117700
rect 411956 117688 411962 117700
rect 416777 117691 416835 117697
rect 416777 117688 416789 117691
rect 411956 117660 416789 117688
rect 411956 117648 411962 117660
rect 416777 117657 416789 117660
rect 416823 117657 416835 117691
rect 416777 117651 416835 117657
rect 417418 117648 417424 117700
rect 417476 117688 417482 117700
rect 417476 117660 422800 117688
rect 417476 117648 417482 117660
rect 234982 117620 234988 117632
rect 226352 117592 234988 117620
rect 226245 117583 226303 117589
rect 234982 117580 234988 117592
rect 235040 117580 235046 117632
rect 236822 117620 236828 117632
rect 235092 117592 236828 117620
rect 193916 117524 200528 117552
rect 193916 117512 193922 117524
rect 201402 117512 201408 117564
rect 201460 117552 201466 117564
rect 235092 117552 235120 117592
rect 236822 117580 236828 117592
rect 236880 117580 236886 117632
rect 242250 117620 242256 117632
rect 239048 117592 242256 117620
rect 201460 117524 235120 117552
rect 201460 117512 201466 117524
rect 236638 117512 236644 117564
rect 236696 117552 236702 117564
rect 239048 117552 239076 117592
rect 242250 117580 242256 117592
rect 242308 117580 242314 117632
rect 244182 117580 244188 117632
rect 244240 117620 244246 117632
rect 258810 117620 258816 117632
rect 244240 117592 258816 117620
rect 244240 117580 244246 117592
rect 258810 117580 258816 117592
rect 258868 117580 258874 117632
rect 294966 117580 294972 117632
rect 295024 117620 295030 117632
rect 311894 117620 311900 117632
rect 295024 117592 311900 117620
rect 295024 117580 295030 117592
rect 311894 117580 311900 117592
rect 311952 117580 311958 117632
rect 314562 117580 314568 117632
rect 314620 117620 314626 117632
rect 320818 117620 320824 117632
rect 314620 117592 320824 117620
rect 314620 117580 314626 117592
rect 320818 117580 320824 117592
rect 320876 117580 320882 117632
rect 330478 117580 330484 117632
rect 330536 117620 330542 117632
rect 331030 117620 331036 117632
rect 330536 117592 331036 117620
rect 330536 117580 330542 117592
rect 331030 117580 331036 117592
rect 331088 117580 331094 117632
rect 356790 117580 356796 117632
rect 356848 117620 356854 117632
rect 356848 117592 384344 117620
rect 356848 117580 356854 117592
rect 236696 117524 239076 117552
rect 239140 117524 240640 117552
rect 236696 117512 236702 117524
rect 130620 117456 143120 117484
rect 147677 117487 147735 117493
rect 130620 117444 130626 117456
rect 147677 117453 147689 117487
rect 147723 117484 147735 117487
rect 150437 117487 150495 117493
rect 150437 117484 150449 117487
rect 147723 117456 150449 117484
rect 147723 117453 147735 117456
rect 147677 117447 147735 117453
rect 150437 117453 150449 117456
rect 150483 117453 150495 117487
rect 150437 117447 150495 117453
rect 154577 117487 154635 117493
rect 154577 117453 154589 117487
rect 154623 117484 154635 117487
rect 164145 117487 164203 117493
rect 164145 117484 164157 117487
rect 154623 117456 164157 117484
rect 154623 117453 154635 117456
rect 154577 117447 154635 117453
rect 164145 117453 164157 117456
rect 164191 117453 164203 117487
rect 164145 117447 164203 117453
rect 208302 117444 208308 117496
rect 208360 117484 208366 117496
rect 208360 117456 229784 117484
rect 208360 117444 208366 117456
rect 67542 117376 67548 117428
rect 67600 117416 67606 117428
rect 71038 117416 71044 117428
rect 67600 117388 71044 117416
rect 67600 117376 67606 117388
rect 71038 117376 71044 117388
rect 71096 117416 71102 117428
rect 168374 117416 168380 117428
rect 71096 117388 168380 117416
rect 71096 117376 71102 117388
rect 168374 117376 168380 117388
rect 168432 117376 168438 117428
rect 211062 117376 211068 117428
rect 211120 117416 211126 117428
rect 220081 117419 220139 117425
rect 220081 117416 220093 117419
rect 211120 117388 220093 117416
rect 211120 117376 211126 117388
rect 220081 117385 220093 117388
rect 220127 117385 220139 117419
rect 220081 117379 220139 117385
rect 225598 117376 225604 117428
rect 225656 117416 225662 117428
rect 229281 117419 229339 117425
rect 229281 117416 229293 117419
rect 225656 117388 229293 117416
rect 225656 117376 225662 117388
rect 229281 117385 229293 117388
rect 229327 117385 229339 117419
rect 229281 117379 229339 117385
rect 97258 117308 97264 117360
rect 97316 117348 97322 117360
rect 97902 117348 97908 117360
rect 97316 117320 97908 117348
rect 97316 117308 97322 117320
rect 97902 117308 97908 117320
rect 97960 117308 97966 117360
rect 111702 117308 111708 117360
rect 111760 117348 111766 117360
rect 148042 117348 148048 117360
rect 111760 117320 148048 117348
rect 111760 117308 111766 117320
rect 148042 117308 148048 117320
rect 148100 117308 148106 117360
rect 171778 117308 171784 117360
rect 171836 117348 171842 117360
rect 212902 117348 212908 117360
rect 171836 117320 212908 117348
rect 171836 117308 171842 117320
rect 212902 117308 212908 117320
rect 212960 117308 212966 117360
rect 214558 117308 214564 117360
rect 214616 117348 214622 117360
rect 226978 117348 226984 117360
rect 214616 117320 226984 117348
rect 214616 117308 214622 117320
rect 226978 117308 226984 117320
rect 227036 117308 227042 117360
rect 229756 117348 229784 117456
rect 230382 117444 230388 117496
rect 230440 117484 230446 117496
rect 237929 117487 237987 117493
rect 237929 117484 237941 117487
rect 230440 117456 237941 117484
rect 230440 117444 230446 117456
rect 237929 117453 237941 117456
rect 237975 117453 237987 117487
rect 237929 117447 237987 117453
rect 238018 117444 238024 117496
rect 238076 117484 238082 117496
rect 239140 117484 239168 117524
rect 240505 117487 240563 117493
rect 240505 117484 240517 117487
rect 238076 117456 239168 117484
rect 239232 117456 240517 117484
rect 238076 117444 238082 117456
rect 229833 117419 229891 117425
rect 229833 117385 229845 117419
rect 229879 117416 229891 117419
rect 239232 117416 239260 117456
rect 240505 117453 240517 117456
rect 240551 117453 240563 117487
rect 240505 117447 240563 117453
rect 240410 117416 240416 117428
rect 229879 117388 239260 117416
rect 239324 117388 240416 117416
rect 229879 117385 229891 117388
rect 229833 117379 229891 117385
rect 239324 117348 239352 117388
rect 240410 117376 240416 117388
rect 240468 117376 240474 117428
rect 240612 117416 240640 117524
rect 241422 117512 241428 117564
rect 241480 117552 241486 117564
rect 257614 117552 257620 117564
rect 241480 117524 257620 117552
rect 241480 117512 241486 117524
rect 257614 117512 257620 117524
rect 257672 117512 257678 117564
rect 266262 117512 266268 117564
rect 266320 117552 266326 117564
rect 270494 117552 270500 117564
rect 266320 117524 270500 117552
rect 266320 117512 266326 117524
rect 270494 117512 270500 117524
rect 270552 117512 270558 117564
rect 280062 117512 280068 117564
rect 280120 117552 280126 117564
rect 283006 117552 283012 117564
rect 280120 117524 283012 117552
rect 280120 117512 280126 117524
rect 283006 117512 283012 117524
rect 283064 117512 283070 117564
rect 299842 117512 299848 117564
rect 299900 117552 299906 117564
rect 315298 117552 315304 117564
rect 299900 117524 315304 117552
rect 299900 117512 299906 117524
rect 315298 117512 315304 117524
rect 315356 117512 315362 117564
rect 354950 117512 354956 117564
rect 355008 117552 355014 117564
rect 369210 117552 369216 117564
rect 355008 117524 369216 117552
rect 355008 117512 355014 117524
rect 369210 117512 369216 117524
rect 369268 117512 369274 117564
rect 240689 117487 240747 117493
rect 240689 117453 240701 117487
rect 240735 117484 240747 117487
rect 241698 117484 241704 117496
rect 240735 117456 241704 117484
rect 240735 117453 240747 117456
rect 240689 117447 240747 117453
rect 241698 117444 241704 117456
rect 241756 117444 241762 117496
rect 241808 117456 245516 117484
rect 241808 117416 241836 117456
rect 240612 117388 241836 117416
rect 243538 117376 243544 117428
rect 243596 117416 243602 117428
rect 245488 117416 245516 117456
rect 245562 117444 245568 117496
rect 245620 117484 245626 117496
rect 260006 117484 260012 117496
rect 245620 117456 260012 117484
rect 245620 117444 245626 117456
rect 260006 117444 260012 117456
rect 260064 117444 260070 117496
rect 267642 117444 267648 117496
rect 267700 117484 267706 117496
rect 271046 117484 271052 117496
rect 267700 117456 271052 117484
rect 267700 117444 267706 117456
rect 271046 117444 271052 117456
rect 271104 117444 271110 117496
rect 282730 117444 282736 117496
rect 282788 117484 282794 117496
rect 284938 117484 284944 117496
rect 282788 117456 284944 117484
rect 282788 117444 282794 117456
rect 284938 117444 284944 117456
rect 284996 117444 285002 117496
rect 320082 117444 320088 117496
rect 320140 117484 320146 117496
rect 324869 117487 324927 117493
rect 324869 117484 324881 117487
rect 320140 117456 324881 117484
rect 320140 117444 320146 117456
rect 324869 117453 324881 117456
rect 324915 117453 324927 117487
rect 324869 117447 324927 117453
rect 324958 117444 324964 117496
rect 325016 117484 325022 117496
rect 326338 117484 326344 117496
rect 325016 117456 326344 117484
rect 325016 117444 325022 117456
rect 326338 117444 326344 117456
rect 326396 117444 326402 117496
rect 328086 117444 328092 117496
rect 328144 117484 328150 117496
rect 328270 117484 328276 117496
rect 328144 117456 328276 117484
rect 328144 117444 328150 117456
rect 328270 117444 328276 117456
rect 328328 117444 328334 117496
rect 367830 117444 367836 117496
rect 367888 117484 367894 117496
rect 377398 117484 377404 117496
rect 367888 117456 377404 117484
rect 367888 117444 367894 117456
rect 377398 117444 377404 117456
rect 377456 117444 377462 117496
rect 384316 117484 384344 117592
rect 391106 117580 391112 117632
rect 391164 117620 391170 117632
rect 391750 117620 391756 117632
rect 391164 117592 391756 117620
rect 391164 117580 391170 117592
rect 391750 117580 391756 117592
rect 391808 117580 391814 117632
rect 404262 117580 404268 117632
rect 404320 117620 404326 117632
rect 422297 117623 422355 117629
rect 422297 117620 422309 117623
rect 404320 117592 422309 117620
rect 404320 117580 404326 117592
rect 422297 117589 422309 117592
rect 422343 117589 422355 117623
rect 422297 117583 422355 117589
rect 384390 117512 384396 117564
rect 384448 117552 384454 117564
rect 398745 117555 398803 117561
rect 398745 117552 398757 117555
rect 384448 117524 398757 117552
rect 384448 117512 384454 117524
rect 398745 117521 398757 117524
rect 398791 117521 398803 117555
rect 398745 117515 398803 117521
rect 398837 117555 398895 117561
rect 398837 117521 398849 117555
rect 398883 117552 398895 117555
rect 413278 117552 413284 117564
rect 398883 117524 413284 117552
rect 398883 117521 398895 117524
rect 398837 117515 398895 117521
rect 413278 117512 413284 117524
rect 413336 117512 413342 117564
rect 416869 117555 416927 117561
rect 416869 117552 416881 117555
rect 413388 117524 416881 117552
rect 393958 117484 393964 117496
rect 384316 117456 393964 117484
rect 393958 117444 393964 117456
rect 394016 117444 394022 117496
rect 399662 117444 399668 117496
rect 399720 117484 399726 117496
rect 400030 117484 400036 117496
rect 399720 117456 400036 117484
rect 399720 117444 399726 117456
rect 400030 117444 400036 117456
rect 400088 117444 400094 117496
rect 413189 117487 413247 117493
rect 413189 117453 413201 117487
rect 413235 117484 413247 117487
rect 413388 117484 413416 117524
rect 416869 117521 416881 117524
rect 416915 117521 416927 117555
rect 416869 117515 416927 117521
rect 419258 117512 419264 117564
rect 419316 117552 419322 117564
rect 420178 117552 420184 117564
rect 419316 117524 420184 117552
rect 419316 117512 419322 117524
rect 420178 117512 420184 117524
rect 420236 117512 420242 117564
rect 420733 117555 420791 117561
rect 420733 117521 420745 117555
rect 420779 117552 420791 117555
rect 422772 117552 422800 117660
rect 422938 117648 422944 117700
rect 422996 117688 423002 117700
rect 424318 117688 424324 117700
rect 422996 117660 424324 117688
rect 422996 117648 423002 117660
rect 424318 117648 424324 117660
rect 424376 117648 424382 117700
rect 424413 117691 424471 117697
rect 424413 117657 424425 117691
rect 424459 117688 424471 117691
rect 427633 117691 427691 117697
rect 427633 117688 427645 117691
rect 424459 117660 427645 117688
rect 424459 117657 424471 117660
rect 424413 117651 424471 117657
rect 427633 117657 427645 117660
rect 427679 117657 427691 117691
rect 427633 117651 427691 117657
rect 427722 117648 427728 117700
rect 427780 117688 427786 117700
rect 493318 117688 493324 117700
rect 427780 117660 493324 117688
rect 427780 117648 427786 117660
rect 493318 117648 493324 117660
rect 493376 117648 493382 117700
rect 423033 117623 423091 117629
rect 423033 117589 423045 117623
rect 423079 117620 423091 117623
rect 482278 117620 482284 117632
rect 423079 117592 482284 117620
rect 423079 117589 423091 117592
rect 423033 117583 423091 117589
rect 482278 117580 482284 117592
rect 482336 117580 482342 117632
rect 496078 117552 496084 117564
rect 420779 117524 422340 117552
rect 422772 117524 496084 117552
rect 420779 117521 420791 117524
rect 420733 117515 420791 117521
rect 413235 117456 413416 117484
rect 413235 117453 413247 117456
rect 413189 117447 413247 117453
rect 413738 117444 413744 117496
rect 413796 117484 413802 117496
rect 416038 117484 416044 117496
rect 413796 117456 416044 117484
rect 413796 117444 413802 117456
rect 416038 117444 416044 117456
rect 416096 117444 416102 117496
rect 418614 117444 418620 117496
rect 418672 117484 418678 117496
rect 419442 117484 419448 117496
rect 418672 117456 419448 117484
rect 418672 117444 418678 117456
rect 419442 117444 419448 117456
rect 419500 117444 419506 117496
rect 419902 117444 419908 117496
rect 419960 117484 419966 117496
rect 420822 117484 420828 117496
rect 419960 117456 420828 117484
rect 419960 117444 419966 117456
rect 420822 117444 420828 117456
rect 420880 117444 420886 117496
rect 421742 117444 421748 117496
rect 421800 117484 421806 117496
rect 422202 117484 422208 117496
rect 421800 117456 422208 117484
rect 421800 117444 421806 117456
rect 422202 117444 422208 117456
rect 422260 117444 422266 117496
rect 422312 117484 422340 117524
rect 496078 117512 496084 117524
rect 496136 117512 496142 117564
rect 424045 117487 424103 117493
rect 424045 117484 424057 117487
rect 422312 117456 424057 117484
rect 424045 117453 424057 117456
rect 424091 117453 424103 117487
rect 424045 117447 424103 117453
rect 424134 117444 424140 117496
rect 424192 117484 424198 117496
rect 424962 117484 424968 117496
rect 424192 117456 424968 117484
rect 424192 117444 424198 117456
rect 424962 117444 424968 117456
rect 425020 117444 425026 117496
rect 425422 117444 425428 117496
rect 425480 117484 425486 117496
rect 426342 117484 426348 117496
rect 425480 117456 426348 117484
rect 425480 117444 425486 117456
rect 426342 117444 426348 117456
rect 426400 117444 426406 117496
rect 427262 117444 427268 117496
rect 427320 117484 427326 117496
rect 427722 117484 427728 117496
rect 427320 117456 427728 117484
rect 427320 117444 427326 117456
rect 427722 117444 427728 117456
rect 427780 117444 427786 117496
rect 428458 117444 428464 117496
rect 428516 117484 428522 117496
rect 430209 117487 430267 117493
rect 430209 117484 430221 117487
rect 428516 117456 430221 117484
rect 428516 117444 428522 117456
rect 430209 117453 430221 117456
rect 430255 117453 430267 117487
rect 430209 117447 430267 117453
rect 430298 117444 430304 117496
rect 430356 117484 430362 117496
rect 431218 117484 431224 117496
rect 430356 117456 431224 117484
rect 430356 117444 430362 117456
rect 431218 117444 431224 117456
rect 431276 117444 431282 117496
rect 432782 117444 432788 117496
rect 432840 117484 432846 117496
rect 433242 117484 433248 117496
rect 432840 117456 433248 117484
rect 432840 117444 432846 117456
rect 433242 117444 433248 117456
rect 433300 117444 433306 117496
rect 433337 117487 433395 117493
rect 433337 117453 433349 117487
rect 433383 117484 433395 117487
rect 507118 117484 507124 117496
rect 433383 117456 507124 117484
rect 433383 117453 433395 117456
rect 433337 117447 433395 117453
rect 507118 117444 507124 117456
rect 507176 117444 507182 117496
rect 247218 117416 247224 117428
rect 243596 117388 245424 117416
rect 245488 117388 247224 117416
rect 243596 117376 243602 117388
rect 229756 117320 239352 117348
rect 239398 117308 239404 117360
rect 239456 117348 239462 117360
rect 244274 117348 244280 117360
rect 239456 117320 244280 117348
rect 239456 117308 239462 117320
rect 244274 117308 244280 117320
rect 244332 117308 244338 117360
rect 245396 117348 245424 117388
rect 247218 117376 247224 117388
rect 247276 117376 247282 117428
rect 247678 117376 247684 117428
rect 247736 117416 247742 117428
rect 251450 117416 251456 117428
rect 247736 117388 251456 117416
rect 247736 117376 247742 117388
rect 251450 117376 251456 117388
rect 251508 117376 251514 117428
rect 252462 117376 252468 117428
rect 252520 117416 252526 117428
rect 263134 117416 263140 117428
rect 252520 117388 263140 117416
rect 252520 117376 252526 117388
rect 263134 117376 263140 117388
rect 263192 117376 263198 117428
rect 269758 117376 269764 117428
rect 269816 117416 269822 117428
rect 271874 117416 271880 117428
rect 269816 117388 271880 117416
rect 269816 117376 269822 117388
rect 271874 117376 271880 117388
rect 271932 117376 271938 117428
rect 272518 117376 272524 117428
rect 272576 117416 272582 117428
rect 273530 117416 273536 117428
rect 272576 117388 273536 117416
rect 272576 117376 272582 117388
rect 273530 117376 273536 117388
rect 273588 117376 273594 117428
rect 278406 117376 278412 117428
rect 278464 117416 278470 117428
rect 279142 117416 279148 117428
rect 278464 117388 279148 117416
rect 278464 117376 278470 117388
rect 279142 117376 279148 117388
rect 279200 117376 279206 117428
rect 282086 117376 282092 117428
rect 282144 117416 282150 117428
rect 283558 117416 283564 117428
rect 282144 117388 283564 117416
rect 282144 117376 282150 117388
rect 283558 117376 283564 117388
rect 283616 117376 283622 117428
rect 289446 117376 289452 117428
rect 289504 117416 289510 117428
rect 294598 117416 294604 117428
rect 289504 117388 294604 117416
rect 289504 117376 289510 117388
rect 294598 117376 294604 117388
rect 294656 117376 294662 117428
rect 318242 117376 318248 117428
rect 318300 117416 318306 117428
rect 322198 117416 322204 117428
rect 318300 117388 322204 117416
rect 318300 117376 318306 117388
rect 322198 117376 322204 117388
rect 322256 117376 322262 117428
rect 332962 117376 332968 117428
rect 333020 117416 333026 117428
rect 333882 117416 333888 117428
rect 333020 117388 333888 117416
rect 333020 117376 333026 117388
rect 333882 117376 333888 117388
rect 333940 117376 333946 117428
rect 371510 117376 371516 117428
rect 371568 117416 371574 117428
rect 372522 117416 372528 117428
rect 371568 117388 372528 117416
rect 371568 117376 371574 117388
rect 372522 117376 372528 117388
rect 372580 117376 372586 117428
rect 391201 117419 391259 117425
rect 391201 117385 391213 117419
rect 391247 117416 391259 117419
rect 396077 117419 396135 117425
rect 396077 117416 396089 117419
rect 391247 117388 396089 117416
rect 391247 117385 391259 117388
rect 391201 117379 391259 117385
rect 396077 117385 396089 117388
rect 396123 117385 396135 117419
rect 396077 117379 396135 117385
rect 405182 117376 405188 117428
rect 405240 117416 405246 117428
rect 405642 117416 405648 117428
rect 405240 117388 405648 117416
rect 405240 117376 405246 117388
rect 405642 117376 405648 117388
rect 405700 117376 405706 117428
rect 408218 117376 408224 117428
rect 408276 117416 408282 117428
rect 486418 117416 486424 117428
rect 408276 117388 486424 117416
rect 408276 117376 408282 117388
rect 486418 117376 486424 117388
rect 486476 117376 486482 117428
rect 249061 117351 249119 117357
rect 249061 117348 249073 117351
rect 245396 117320 249073 117348
rect 249061 117317 249073 117320
rect 249107 117317 249119 117351
rect 249061 117311 249119 117317
rect 250438 117308 250444 117360
rect 250496 117348 250502 117360
rect 254578 117348 254584 117360
rect 250496 117320 254584 117348
rect 250496 117308 250502 117320
rect 254578 117308 254584 117320
rect 254636 117308 254642 117360
rect 259362 117308 259368 117360
rect 259420 117348 259426 117360
rect 266814 117348 266820 117360
rect 259420 117320 266820 117348
rect 259420 117308 259426 117320
rect 266814 117308 266820 117320
rect 266872 117308 266878 117360
rect 268378 117308 268384 117360
rect 268436 117348 268442 117360
rect 269850 117348 269856 117360
rect 268436 117320 269856 117348
rect 268436 117308 268442 117320
rect 269850 117308 269856 117320
rect 269908 117308 269914 117360
rect 273162 117308 273168 117360
rect 273220 117348 273226 117360
rect 274174 117348 274180 117360
rect 273220 117320 274180 117348
rect 273220 117308 273226 117320
rect 274174 117308 274180 117320
rect 274232 117308 274238 117360
rect 277854 117308 277860 117360
rect 277912 117348 277918 117360
rect 278866 117348 278872 117360
rect 277912 117320 278872 117348
rect 277912 117308 277918 117320
rect 278866 117308 278872 117320
rect 278924 117308 278930 117360
rect 279050 117308 279056 117360
rect 279108 117348 279114 117360
rect 280338 117348 280344 117360
rect 279108 117320 280344 117348
rect 279108 117308 279114 117320
rect 280338 117308 280344 117320
rect 280396 117308 280402 117360
rect 280890 117308 280896 117360
rect 280948 117348 280954 117360
rect 281350 117348 281356 117360
rect 280948 117320 281356 117348
rect 280948 117308 280954 117320
rect 281350 117308 281356 117320
rect 281408 117308 281414 117360
rect 283374 117308 283380 117360
rect 283432 117348 283438 117360
rect 284202 117348 284208 117360
rect 283432 117320 284208 117348
rect 283432 117308 283438 117320
rect 284202 117308 284208 117320
rect 284260 117308 284266 117360
rect 285214 117308 285220 117360
rect 285272 117348 285278 117360
rect 285582 117348 285588 117360
rect 285272 117320 285588 117348
rect 285272 117308 285278 117320
rect 285582 117308 285588 117320
rect 285640 117308 285646 117360
rect 286410 117308 286416 117360
rect 286468 117348 286474 117360
rect 286962 117348 286968 117360
rect 286468 117320 286968 117348
rect 286468 117308 286474 117320
rect 286962 117308 286968 117320
rect 287020 117308 287026 117360
rect 287606 117308 287612 117360
rect 287664 117348 287670 117360
rect 288342 117348 288348 117360
rect 287664 117320 288348 117348
rect 287664 117308 287670 117320
rect 288342 117308 288348 117320
rect 288400 117308 288406 117360
rect 289998 117308 290004 117360
rect 290056 117348 290062 117360
rect 291102 117348 291108 117360
rect 290056 117320 291108 117348
rect 290056 117308 290062 117320
rect 291102 117308 291108 117320
rect 291160 117308 291166 117360
rect 291930 117308 291936 117360
rect 291988 117348 291994 117360
rect 292482 117348 292488 117360
rect 291988 117320 292488 117348
rect 291988 117308 291994 117320
rect 292482 117308 292488 117320
rect 292540 117308 292546 117360
rect 301130 117308 301136 117360
rect 301188 117348 301194 117360
rect 302142 117348 302148 117360
rect 301188 117320 302148 117348
rect 301188 117308 301194 117320
rect 302142 117308 302148 117320
rect 302200 117308 302206 117360
rect 302970 117308 302976 117360
rect 303028 117348 303034 117360
rect 303522 117348 303528 117360
rect 303028 117320 303528 117348
rect 303028 117308 303034 117320
rect 303522 117308 303528 117320
rect 303580 117308 303586 117360
rect 305362 117308 305368 117360
rect 305420 117348 305426 117360
rect 306282 117348 306288 117360
rect 305420 117320 306288 117348
rect 305420 117308 305426 117320
rect 306282 117308 306288 117320
rect 306340 117308 306346 117360
rect 312722 117308 312728 117360
rect 312780 117348 312786 117360
rect 313182 117348 313188 117360
rect 312780 117320 313188 117348
rect 312780 117308 312786 117320
rect 313182 117308 313188 117320
rect 313240 117308 313246 117360
rect 313918 117308 313924 117360
rect 313976 117348 313982 117360
rect 314562 117348 314568 117360
rect 313976 117320 314568 117348
rect 313976 117308 313982 117320
rect 314562 117308 314568 117320
rect 314620 117308 314626 117360
rect 315206 117308 315212 117360
rect 315264 117348 315270 117360
rect 315850 117348 315856 117360
rect 315264 117320 315856 117348
rect 315264 117308 315270 117320
rect 315850 117308 315856 117320
rect 315908 117308 315914 117360
rect 316402 117308 316408 117360
rect 316460 117348 316466 117360
rect 317322 117348 317328 117360
rect 316460 117320 317328 117348
rect 316460 117308 316466 117320
rect 317322 117308 317328 117320
rect 317380 117308 317386 117360
rect 319438 117308 319444 117360
rect 319496 117348 319502 117360
rect 320082 117348 320088 117360
rect 319496 117320 320088 117348
rect 319496 117308 319502 117320
rect 320082 117308 320088 117320
rect 320140 117308 320146 117360
rect 320726 117308 320732 117360
rect 320784 117348 320790 117360
rect 321370 117348 321376 117360
rect 320784 117320 321376 117348
rect 320784 117308 320790 117320
rect 321370 117308 321376 117320
rect 321428 117308 321434 117360
rect 323762 117308 323768 117360
rect 323820 117348 323826 117360
rect 324222 117348 324228 117360
rect 323820 117320 324228 117348
rect 323820 117308 323826 117320
rect 324222 117308 324228 117320
rect 324280 117308 324286 117360
rect 326246 117308 326252 117360
rect 326304 117348 326310 117360
rect 326982 117348 326988 117360
rect 326304 117320 326988 117348
rect 326304 117308 326310 117320
rect 326982 117308 326988 117320
rect 327040 117308 327046 117360
rect 327442 117308 327448 117360
rect 327500 117348 327506 117360
rect 328362 117348 328368 117360
rect 327500 117320 328368 117348
rect 327500 117308 327506 117320
rect 328362 117308 328368 117320
rect 328420 117308 328426 117360
rect 331674 117308 331680 117360
rect 331732 117348 331738 117360
rect 332502 117348 332508 117360
rect 331732 117320 332508 117348
rect 331732 117308 331738 117320
rect 332502 117308 332508 117320
rect 332560 117308 332566 117360
rect 333514 117308 333520 117360
rect 333572 117348 333578 117360
rect 333790 117348 333796 117360
rect 333572 117320 333796 117348
rect 333572 117308 333578 117320
rect 333790 117308 333796 117320
rect 333848 117308 333854 117360
rect 334802 117308 334808 117360
rect 334860 117348 334866 117360
rect 335262 117348 335268 117360
rect 334860 117320 335268 117348
rect 334860 117308 334866 117320
rect 335262 117308 335268 117320
rect 335320 117308 335326 117360
rect 335998 117308 336004 117360
rect 336056 117348 336062 117360
rect 336642 117348 336648 117360
rect 336056 117320 336648 117348
rect 336056 117308 336062 117320
rect 336642 117308 336648 117320
rect 336700 117308 336706 117360
rect 337194 117308 337200 117360
rect 337252 117348 337258 117360
rect 338022 117348 338028 117360
rect 337252 117320 338028 117348
rect 337252 117308 337258 117320
rect 338022 117308 338028 117320
rect 338080 117308 338086 117360
rect 339034 117308 339040 117360
rect 339092 117348 339098 117360
rect 339402 117348 339408 117360
rect 339092 117320 339408 117348
rect 339092 117308 339098 117320
rect 339402 117308 339408 117320
rect 339460 117308 339466 117360
rect 340322 117308 340328 117360
rect 340380 117348 340386 117360
rect 340782 117348 340788 117360
rect 340380 117320 340788 117348
rect 340380 117308 340386 117320
rect 340782 117308 340788 117320
rect 340840 117308 340846 117360
rect 341518 117308 341524 117360
rect 341576 117348 341582 117360
rect 342162 117348 342168 117360
rect 341576 117320 342168 117348
rect 341576 117308 341582 117320
rect 342162 117308 342168 117320
rect 342220 117308 342226 117360
rect 342714 117308 342720 117360
rect 342772 117348 342778 117360
rect 343542 117348 343548 117360
rect 342772 117320 343548 117348
rect 342772 117308 342778 117320
rect 343542 117308 343548 117320
rect 343600 117308 343606 117360
rect 344554 117308 344560 117360
rect 344612 117348 344618 117360
rect 344830 117348 344836 117360
rect 344612 117320 344836 117348
rect 344612 117308 344618 117320
rect 344830 117308 344836 117320
rect 344888 117308 344894 117360
rect 347038 117308 347044 117360
rect 347096 117348 347102 117360
rect 347682 117348 347688 117360
rect 347096 117320 347688 117348
rect 347096 117308 347102 117320
rect 347682 117308 347688 117320
rect 347740 117308 347746 117360
rect 348234 117308 348240 117360
rect 348292 117348 348298 117360
rect 349062 117348 349068 117360
rect 348292 117320 349068 117348
rect 348292 117308 348298 117320
rect 349062 117308 349068 117320
rect 349120 117308 349126 117360
rect 350074 117308 350080 117360
rect 350132 117348 350138 117360
rect 350442 117348 350448 117360
rect 350132 117320 350448 117348
rect 350132 117308 350138 117320
rect 350442 117308 350448 117320
rect 350500 117308 350506 117360
rect 351270 117308 351276 117360
rect 351328 117348 351334 117360
rect 351822 117348 351828 117360
rect 351328 117320 351828 117348
rect 351328 117308 351334 117320
rect 351822 117308 351828 117320
rect 351880 117308 351886 117360
rect 352558 117308 352564 117360
rect 352616 117348 352622 117360
rect 353202 117348 353208 117360
rect 352616 117320 353208 117348
rect 352616 117308 352622 117320
rect 353202 117308 353208 117320
rect 353260 117308 353266 117360
rect 353754 117308 353760 117360
rect 353812 117348 353818 117360
rect 354582 117348 354588 117360
rect 353812 117320 354588 117348
rect 353812 117308 353818 117320
rect 354582 117308 354588 117320
rect 354640 117308 354646 117360
rect 355594 117308 355600 117360
rect 355652 117348 355658 117360
rect 355962 117348 355968 117360
rect 355652 117320 355968 117348
rect 355652 117308 355658 117320
rect 355962 117308 355968 117320
rect 356020 117308 356026 117360
rect 358078 117308 358084 117360
rect 358136 117348 358142 117360
rect 358630 117348 358636 117360
rect 358136 117320 358636 117348
rect 358136 117308 358142 117320
rect 358630 117308 358636 117320
rect 358688 117308 358694 117360
rect 359274 117308 359280 117360
rect 359332 117348 359338 117360
rect 360102 117348 360108 117360
rect 359332 117320 360108 117348
rect 359332 117308 359338 117320
rect 360102 117308 360108 117320
rect 360160 117308 360166 117360
rect 361114 117308 361120 117360
rect 361172 117348 361178 117360
rect 361482 117348 361488 117360
rect 361172 117320 361488 117348
rect 361172 117308 361178 117320
rect 361482 117308 361488 117320
rect 361540 117308 361546 117360
rect 363598 117308 363604 117360
rect 363656 117348 363662 117360
rect 364242 117348 364248 117360
rect 363656 117320 364248 117348
rect 363656 117308 363662 117320
rect 364242 117308 364248 117320
rect 364300 117308 364306 117360
rect 364794 117308 364800 117360
rect 364852 117348 364858 117360
rect 365622 117348 365628 117360
rect 364852 117320 365628 117348
rect 364852 117308 364858 117320
rect 365622 117308 365628 117320
rect 365680 117308 365686 117360
rect 366634 117308 366640 117360
rect 366692 117348 366698 117360
rect 367002 117348 367008 117360
rect 366692 117320 367008 117348
rect 366692 117308 366698 117320
rect 367002 117308 367008 117320
rect 367060 117308 367066 117360
rect 369026 117308 369032 117360
rect 369084 117348 369090 117360
rect 369762 117348 369768 117360
rect 369084 117320 369768 117348
rect 369084 117308 369090 117320
rect 369762 117308 369768 117320
rect 369820 117308 369826 117360
rect 370314 117308 370320 117360
rect 370372 117348 370378 117360
rect 371142 117348 371148 117360
rect 370372 117320 371148 117348
rect 370372 117308 370378 117320
rect 371142 117308 371148 117320
rect 371200 117308 371206 117360
rect 372154 117308 372160 117360
rect 372212 117348 372218 117360
rect 372430 117348 372436 117360
rect 372212 117320 372436 117348
rect 372212 117308 372218 117320
rect 372430 117308 372436 117320
rect 372488 117308 372494 117360
rect 374546 117308 374552 117360
rect 374604 117348 374610 117360
rect 375190 117348 375196 117360
rect 374604 117320 375196 117348
rect 374604 117308 374610 117320
rect 375190 117308 375196 117320
rect 375248 117308 375254 117360
rect 375834 117308 375840 117360
rect 375892 117348 375898 117360
rect 376662 117348 376668 117360
rect 375892 117320 376668 117348
rect 375892 117308 375898 117320
rect 376662 117308 376668 117320
rect 376720 117308 376726 117360
rect 377674 117308 377680 117360
rect 377732 117348 377738 117360
rect 378042 117348 378048 117360
rect 377732 117320 378048 117348
rect 377732 117308 377738 117320
rect 378042 117308 378048 117320
rect 378100 117308 378106 117360
rect 378870 117308 378876 117360
rect 378928 117348 378934 117360
rect 379422 117348 379428 117360
rect 378928 117320 379428 117348
rect 378928 117308 378934 117320
rect 379422 117308 379428 117320
rect 379480 117308 379486 117360
rect 380066 117308 380072 117360
rect 380124 117348 380130 117360
rect 380802 117348 380808 117360
rect 380124 117320 380808 117348
rect 380124 117308 380130 117320
rect 380802 117308 380808 117320
rect 380860 117308 380866 117360
rect 381354 117308 381360 117360
rect 381412 117348 381418 117360
rect 382182 117348 382188 117360
rect 381412 117320 382188 117348
rect 381412 117308 381418 117320
rect 382182 117308 382188 117320
rect 382240 117308 382246 117360
rect 382550 117308 382556 117360
rect 382608 117348 382614 117360
rect 383562 117348 383568 117360
rect 382608 117320 383568 117348
rect 382608 117308 382614 117320
rect 383562 117308 383568 117320
rect 383620 117308 383626 117360
rect 385586 117308 385592 117360
rect 385644 117348 385650 117360
rect 386322 117348 386328 117360
rect 385644 117320 386328 117348
rect 385644 117308 385650 117320
rect 386322 117308 386328 117320
rect 386380 117308 386386 117360
rect 386782 117308 386788 117360
rect 386840 117348 386846 117360
rect 387610 117348 387616 117360
rect 386840 117320 387616 117348
rect 386840 117308 386846 117320
rect 387610 117308 387616 117320
rect 387668 117308 387674 117360
rect 388070 117308 388076 117360
rect 388128 117348 388134 117360
rect 389082 117348 389088 117360
rect 388128 117320 389088 117348
rect 388128 117308 388134 117320
rect 389082 117308 389088 117320
rect 389140 117308 389146 117360
rect 392302 117308 392308 117360
rect 392360 117348 392366 117360
rect 393130 117348 393136 117360
rect 392360 117320 393136 117348
rect 392360 117308 392366 117320
rect 393130 117308 393136 117320
rect 393188 117308 393194 117360
rect 396626 117308 396632 117360
rect 396684 117348 396690 117360
rect 397362 117348 397368 117360
rect 396684 117320 397368 117348
rect 396684 117308 396690 117320
rect 397362 117308 397368 117320
rect 397420 117308 397426 117360
rect 397822 117308 397828 117360
rect 397880 117348 397886 117360
rect 398742 117348 398748 117360
rect 397880 117320 398748 117348
rect 397880 117308 397886 117320
rect 398742 117308 398748 117320
rect 398800 117308 398806 117360
rect 399110 117308 399116 117360
rect 399168 117348 399174 117360
rect 400122 117348 400128 117360
rect 399168 117320 400128 117348
rect 399168 117308 399174 117320
rect 400122 117308 400128 117320
rect 400180 117308 400186 117360
rect 402146 117308 402152 117360
rect 402204 117348 402210 117360
rect 402790 117348 402796 117360
rect 402204 117320 402796 117348
rect 402204 117308 402210 117320
rect 402790 117308 402796 117320
rect 402848 117308 402854 117360
rect 403342 117308 403348 117360
rect 403400 117348 403406 117360
rect 404262 117348 404268 117360
rect 403400 117320 404268 117348
rect 403400 117308 403406 117320
rect 404262 117308 404268 117320
rect 404320 117308 404326 117360
rect 406378 117308 406384 117360
rect 406436 117348 406442 117360
rect 407022 117348 407028 117360
rect 406436 117320 407028 117348
rect 406436 117308 406442 117320
rect 407022 117308 407028 117320
rect 407080 117308 407086 117360
rect 407666 117308 407672 117360
rect 407724 117348 407730 117360
rect 408402 117348 408408 117360
rect 407724 117320 408408 117348
rect 407724 117308 407730 117320
rect 408402 117308 408408 117320
rect 408460 117308 408466 117360
rect 408862 117308 408868 117360
rect 408920 117348 408926 117360
rect 409690 117348 409696 117360
rect 408920 117320 409696 117348
rect 408920 117308 408926 117320
rect 409690 117308 409696 117320
rect 409748 117308 409754 117360
rect 410702 117308 410708 117360
rect 410760 117348 410766 117360
rect 411162 117348 411168 117360
rect 410760 117320 411168 117348
rect 410760 117308 410766 117320
rect 411162 117308 411168 117320
rect 411220 117308 411226 117360
rect 413186 117308 413192 117360
rect 413244 117348 413250 117360
rect 413922 117348 413928 117360
rect 413244 117320 413928 117348
rect 413244 117308 413250 117320
rect 413922 117308 413928 117320
rect 413980 117308 413986 117360
rect 414382 117308 414388 117360
rect 414440 117348 414446 117360
rect 415302 117348 415308 117360
rect 414440 117320 415308 117348
rect 414440 117308 414446 117320
rect 415302 117308 415308 117320
rect 415360 117308 415366 117360
rect 416222 117308 416228 117360
rect 416280 117348 416286 117360
rect 416682 117348 416688 117360
rect 416280 117320 416688 117348
rect 416280 117308 416286 117320
rect 416682 117308 416688 117320
rect 416740 117308 416746 117360
rect 416777 117351 416835 117357
rect 416777 117317 416789 117351
rect 416823 117348 416835 117351
rect 489178 117348 489184 117360
rect 416823 117320 489184 117348
rect 416823 117317 416835 117320
rect 416777 117311 416835 117317
rect 489178 117308 489184 117320
rect 489236 117308 489242 117360
rect 122834 117240 122840 117292
rect 122892 117280 122898 117292
rect 133782 117280 133788 117292
rect 122892 117252 133788 117280
rect 122892 117240 122898 117252
rect 133782 117240 133788 117252
rect 133840 117240 133846 117292
rect 137925 117283 137983 117289
rect 137925 117249 137937 117283
rect 137971 117280 137983 117283
rect 138017 117283 138075 117289
rect 138017 117280 138029 117283
rect 137971 117252 138029 117280
rect 137971 117249 137983 117252
rect 137925 117243 137983 117249
rect 138017 117249 138029 117252
rect 138063 117249 138075 117283
rect 138017 117243 138075 117249
rect 396077 117283 396135 117289
rect 396077 117249 396089 117283
rect 396123 117280 396135 117283
rect 402238 117280 402244 117292
rect 396123 117252 402244 117280
rect 396123 117249 396135 117252
rect 396077 117243 396135 117249
rect 402238 117240 402244 117252
rect 402296 117240 402302 117292
rect 430209 117283 430267 117289
rect 430209 117249 430221 117283
rect 430255 117280 430267 117283
rect 433337 117283 433395 117289
rect 433337 117280 433349 117283
rect 430255 117252 433349 117280
rect 430255 117249 430267 117252
rect 430209 117243 430267 117249
rect 433337 117249 433349 117252
rect 433383 117249 433395 117283
rect 433337 117243 433395 117249
rect 198734 116560 198740 116612
rect 198792 116600 198798 116612
rect 199470 116600 199476 116612
rect 198792 116572 199476 116600
rect 198792 116560 198798 116572
rect 199470 116560 199476 116572
rect 199528 116560 199534 116612
rect 200114 116560 200120 116612
rect 200172 116600 200178 116612
rect 200666 116600 200672 116612
rect 200172 116572 200672 116600
rect 200172 116560 200178 116572
rect 200666 116560 200672 116572
rect 200724 116560 200730 116612
rect 201494 116560 201500 116612
rect 201552 116600 201558 116612
rect 201862 116600 201868 116612
rect 201552 116572 201868 116600
rect 201552 116560 201558 116572
rect 201862 116560 201868 116572
rect 201920 116560 201926 116612
rect 202966 116560 202972 116612
rect 203024 116600 203030 116612
rect 203702 116600 203708 116612
rect 203024 116572 203708 116600
rect 203024 116560 203030 116572
rect 203702 116560 203708 116572
rect 203760 116560 203766 116612
rect 204254 116560 204260 116612
rect 204312 116600 204318 116612
rect 204898 116600 204904 116612
rect 204312 116572 204904 116600
rect 204312 116560 204318 116572
rect 204898 116560 204904 116572
rect 204956 116560 204962 116612
rect 190730 115948 190736 116000
rect 190788 115988 190794 116000
rect 191006 115988 191012 116000
rect 190788 115960 191012 115988
rect 190788 115948 190794 115960
rect 191006 115948 191012 115960
rect 191064 115948 191070 116000
rect 272242 115948 272248 116000
rect 272300 115988 272306 116000
rect 272426 115988 272432 116000
rect 272300 115960 272432 115988
rect 272300 115948 272306 115960
rect 272426 115948 272432 115960
rect 272484 115948 272490 116000
rect 322382 115948 322388 116000
rect 322440 115988 322446 116000
rect 322566 115988 322572 116000
rect 322440 115960 322572 115988
rect 322440 115948 322446 115960
rect 322566 115948 322572 115960
rect 322624 115948 322630 116000
rect 382918 115948 382924 116000
rect 382976 115988 382982 116000
rect 383102 115988 383108 116000
rect 382976 115960 383108 115988
rect 382976 115948 382982 115960
rect 383102 115948 383108 115960
rect 383160 115948 383166 116000
rect 133782 115880 133788 115932
rect 133840 115920 133846 115932
rect 134518 115920 134524 115932
rect 133840 115892 134524 115920
rect 133840 115880 133846 115892
rect 134518 115880 134524 115892
rect 134576 115880 134582 115932
rect 150802 115880 150808 115932
rect 150860 115920 150866 115932
rect 151354 115920 151360 115932
rect 150860 115892 151360 115920
rect 150860 115880 150866 115892
rect 151354 115880 151360 115892
rect 151412 115880 151418 115932
rect 173986 115880 173992 115932
rect 174044 115920 174050 115932
rect 174354 115920 174360 115932
rect 174044 115892 174360 115920
rect 174044 115880 174050 115892
rect 174354 115880 174360 115892
rect 174412 115880 174418 115932
rect 248322 115880 248328 115932
rect 248380 115920 248386 115932
rect 248414 115920 248420 115932
rect 248380 115892 248420 115920
rect 248380 115880 248386 115892
rect 248414 115880 248420 115892
rect 248472 115880 248478 115932
rect 276014 115880 276020 115932
rect 276072 115920 276078 115932
rect 276106 115920 276112 115932
rect 276072 115892 276112 115920
rect 276072 115880 276078 115892
rect 276106 115880 276112 115892
rect 276164 115880 276170 115932
rect 301682 115880 301688 115932
rect 301740 115920 301746 115932
rect 301958 115920 301964 115932
rect 301740 115892 301964 115920
rect 301740 115880 301746 115892
rect 301958 115880 301964 115892
rect 302016 115880 302022 115932
rect 388714 115880 388720 115932
rect 388772 115920 388778 115932
rect 388898 115920 388904 115932
rect 388772 115892 388904 115920
rect 388772 115880 388778 115892
rect 388898 115880 388904 115892
rect 388956 115880 388962 115932
rect 403897 115923 403955 115929
rect 403897 115889 403909 115923
rect 403943 115920 403955 115923
rect 404078 115920 404084 115932
rect 403943 115892 404084 115920
rect 403943 115889 403955 115892
rect 403897 115883 403955 115889
rect 404078 115880 404084 115892
rect 404136 115880 404142 115932
rect 414842 115880 414848 115932
rect 414900 115920 414906 115932
rect 414934 115920 414940 115932
rect 414900 115892 414940 115920
rect 414900 115880 414906 115892
rect 414934 115880 414940 115892
rect 414992 115880 414998 115932
rect 420546 115920 420552 115932
rect 420507 115892 420552 115920
rect 420546 115880 420552 115892
rect 420604 115880 420610 115932
rect 426066 115880 426072 115932
rect 426124 115920 426130 115932
rect 426250 115920 426256 115932
rect 426124 115892 426256 115920
rect 426124 115880 426130 115892
rect 426250 115880 426256 115892
rect 426308 115880 426314 115932
rect 431494 115920 431500 115932
rect 431455 115892 431500 115920
rect 431494 115880 431500 115892
rect 431552 115880 431558 115932
rect 202874 114520 202880 114572
rect 202932 114560 202938 114572
rect 203150 114560 203156 114572
rect 202932 114532 203156 114560
rect 202932 114520 202938 114532
rect 203150 114520 203156 114532
rect 203208 114520 203214 114572
rect 215386 114520 215392 114572
rect 215444 114560 215450 114572
rect 215938 114560 215944 114572
rect 215444 114532 215944 114560
rect 215444 114520 215450 114532
rect 215938 114520 215944 114532
rect 215996 114520 216002 114572
rect 232222 114520 232228 114572
rect 232280 114560 232286 114572
rect 232590 114560 232596 114572
rect 232280 114532 232596 114560
rect 232280 114520 232286 114532
rect 232590 114520 232596 114532
rect 232648 114520 232654 114572
rect 325694 114560 325700 114572
rect 325655 114532 325700 114560
rect 325694 114520 325700 114532
rect 325752 114520 325758 114572
rect 174173 114495 174231 114501
rect 174173 114461 174185 114495
rect 174219 114492 174231 114495
rect 174354 114492 174360 114504
rect 174219 114464 174360 114492
rect 174219 114461 174231 114464
rect 174173 114455 174231 114461
rect 174354 114452 174360 114464
rect 174412 114452 174418 114504
rect 230382 114492 230388 114504
rect 230343 114464 230388 114492
rect 230382 114452 230388 114464
rect 230440 114452 230446 114504
rect 248325 114495 248383 114501
rect 248325 114461 248337 114495
rect 248371 114492 248383 114495
rect 248414 114492 248420 114504
rect 248371 114464 248420 114492
rect 248371 114461 248383 114464
rect 248325 114455 248383 114461
rect 248414 114452 248420 114464
rect 248472 114452 248478 114504
rect 135254 113840 135260 113892
rect 135312 113880 135318 113892
rect 135714 113880 135720 113892
rect 135312 113852 135720 113880
rect 135312 113840 135318 113852
rect 135714 113840 135720 113852
rect 135772 113840 135778 113892
rect 139394 113840 139400 113892
rect 139452 113880 139458 113892
rect 140038 113880 140044 113892
rect 139452 113852 140044 113880
rect 139452 113840 139458 113852
rect 140038 113840 140044 113852
rect 140096 113840 140102 113892
rect 151814 113840 151820 113892
rect 151872 113880 151878 113892
rect 152274 113880 152280 113892
rect 151872 113852 152280 113880
rect 151872 113840 151878 113852
rect 152274 113840 152280 113852
rect 152332 113840 152338 113892
rect 153194 113840 153200 113892
rect 153252 113880 153258 113892
rect 154114 113880 154120 113892
rect 153252 113852 154120 113880
rect 153252 113840 153258 113852
rect 154114 113840 154120 113852
rect 154172 113840 154178 113892
rect 155954 113840 155960 113892
rect 156012 113880 156018 113892
rect 156598 113880 156604 113892
rect 156012 113852 156604 113880
rect 156012 113840 156018 113852
rect 156598 113840 156604 113852
rect 156656 113840 156662 113892
rect 166994 113840 167000 113892
rect 167052 113880 167058 113892
rect 167638 113880 167644 113892
rect 167052 113852 167644 113880
rect 167052 113840 167058 113852
rect 167638 113840 167644 113852
rect 167696 113840 167702 113892
rect 169846 113840 169852 113892
rect 169904 113880 169910 113892
rect 170674 113880 170680 113892
rect 169904 113852 170680 113880
rect 169904 113840 169910 113852
rect 170674 113840 170680 113852
rect 170732 113840 170738 113892
rect 172514 113840 172520 113892
rect 172572 113880 172578 113892
rect 173066 113880 173072 113892
rect 172572 113852 173072 113880
rect 172572 113840 172578 113852
rect 173066 113840 173072 113852
rect 173124 113840 173130 113892
rect 175366 113840 175372 113892
rect 175424 113880 175430 113892
rect 176194 113880 176200 113892
rect 175424 113852 176200 113880
rect 175424 113840 175430 113852
rect 176194 113840 176200 113852
rect 176252 113840 176258 113892
rect 178034 113840 178040 113892
rect 178092 113880 178098 113892
rect 178586 113880 178592 113892
rect 178092 113852 178592 113880
rect 178092 113840 178098 113852
rect 178586 113840 178592 113852
rect 178644 113840 178650 113892
rect 186406 113840 186412 113892
rect 186464 113880 186470 113892
rect 186590 113880 186596 113892
rect 186464 113852 186596 113880
rect 186464 113840 186470 113852
rect 186590 113840 186596 113852
rect 186648 113840 186654 113892
rect 191926 113840 191932 113892
rect 191984 113880 191990 113892
rect 192662 113880 192668 113892
rect 191984 113852 192668 113880
rect 191984 113840 191990 113852
rect 192662 113840 192668 113852
rect 192720 113840 192726 113892
rect 194686 113840 194692 113892
rect 194744 113880 194750 113892
rect 195146 113880 195152 113892
rect 194744 113852 195152 113880
rect 194744 113840 194750 113852
rect 195146 113840 195152 113852
rect 195204 113840 195210 113892
rect 205634 113840 205640 113892
rect 205692 113880 205698 113892
rect 206186 113880 206192 113892
rect 205692 113852 206192 113880
rect 205692 113840 205698 113852
rect 206186 113840 206192 113852
rect 206244 113840 206250 113892
rect 208486 113840 208492 113892
rect 208544 113880 208550 113892
rect 209222 113880 209228 113892
rect 208544 113852 209228 113880
rect 208544 113840 208550 113852
rect 209222 113840 209228 113852
rect 209280 113840 209286 113892
rect 209866 113840 209872 113892
rect 209924 113880 209930 113892
rect 210418 113880 210424 113892
rect 209924 113852 210424 113880
rect 209924 113840 209930 113852
rect 210418 113840 210424 113852
rect 210476 113840 210482 113892
rect 211154 113840 211160 113892
rect 211212 113880 211218 113892
rect 211706 113880 211712 113892
rect 211212 113852 211712 113880
rect 211212 113840 211218 113852
rect 211706 113840 211712 113852
rect 211764 113840 211770 113892
rect 219526 113840 219532 113892
rect 219584 113880 219590 113892
rect 219710 113880 219716 113892
rect 219584 113852 219716 113880
rect 219584 113840 219590 113852
rect 219710 113840 219716 113852
rect 219768 113840 219774 113892
rect 229186 113840 229192 113892
rect 229244 113880 229250 113892
rect 230014 113880 230020 113892
rect 229244 113852 230020 113880
rect 229244 113840 229250 113852
rect 230014 113840 230020 113852
rect 230072 113840 230078 113892
rect 223666 113092 223672 113144
rect 223724 113132 223730 113144
rect 224494 113132 224500 113144
rect 223724 113104 224500 113132
rect 223724 113092 223730 113104
rect 224494 113092 224500 113104
rect 224552 113092 224558 113144
rect 229186 113092 229192 113144
rect 229244 113132 229250 113144
rect 229281 113135 229339 113141
rect 229281 113132 229293 113135
rect 229244 113104 229293 113132
rect 229244 113092 229250 113104
rect 229281 113101 229293 113104
rect 229327 113101 229339 113135
rect 229281 113095 229339 113101
rect 136726 112480 136732 112532
rect 136784 112520 136790 112532
rect 137554 112520 137560 112532
rect 136784 112492 137560 112520
rect 136784 112480 136790 112492
rect 137554 112480 137560 112492
rect 137612 112480 137618 112532
rect 140774 111868 140780 111920
rect 140832 111908 140838 111920
rect 141234 111908 141240 111920
rect 140832 111880 141240 111908
rect 140832 111868 140838 111880
rect 141234 111868 141240 111880
rect 141292 111868 141298 111920
rect 436922 111732 436928 111784
rect 436980 111772 436986 111784
rect 579798 111772 579804 111784
rect 436980 111744 579804 111772
rect 436980 111732 436986 111744
rect 579798 111732 579804 111744
rect 579856 111732 579862 111784
rect 189074 111528 189080 111580
rect 189132 111568 189138 111580
rect 189626 111568 189632 111580
rect 189132 111540 189632 111568
rect 189132 111528 189138 111540
rect 189626 111528 189632 111540
rect 189684 111528 189690 111580
rect 244458 109080 244464 109132
rect 244516 109080 244522 109132
rect 143626 109012 143632 109064
rect 143684 109052 143690 109064
rect 144178 109052 144184 109064
rect 143684 109024 144184 109052
rect 143684 109012 143690 109024
rect 144178 109012 144184 109024
rect 144236 109012 144242 109064
rect 192018 109012 192024 109064
rect 192076 109012 192082 109064
rect 192036 108984 192064 109012
rect 244476 108996 244504 109080
rect 387518 109012 387524 109064
rect 387576 109052 387582 109064
rect 387702 109052 387708 109064
rect 387576 109024 387708 109052
rect 387576 109012 387582 109024
rect 387702 109012 387708 109024
rect 387760 109012 387766 109064
rect 393038 109012 393044 109064
rect 393096 109052 393102 109064
rect 393222 109052 393228 109064
rect 393096 109024 393228 109052
rect 393096 109012 393102 109024
rect 393222 109012 393228 109024
rect 393280 109012 393286 109064
rect 192202 108984 192208 108996
rect 192036 108956 192208 108984
rect 192202 108944 192208 108956
rect 192260 108944 192266 108996
rect 244458 108944 244464 108996
rect 244516 108944 244522 108996
rect 420546 108984 420552 108996
rect 420507 108956 420552 108984
rect 420546 108944 420552 108956
rect 420604 108944 420610 108996
rect 431497 108987 431555 108993
rect 431497 108953 431509 108987
rect 431543 108984 431555 108987
rect 431678 108984 431684 108996
rect 431543 108956 431684 108984
rect 431543 108953 431555 108956
rect 431497 108947 431555 108953
rect 431678 108944 431684 108956
rect 431736 108944 431742 108996
rect 186130 106292 186136 106344
rect 186188 106292 186194 106344
rect 403894 106332 403900 106344
rect 403855 106304 403900 106332
rect 403894 106292 403900 106304
rect 403952 106292 403958 106344
rect 128906 106264 128912 106276
rect 128867 106236 128912 106264
rect 128906 106224 128912 106236
rect 128964 106224 128970 106276
rect 133966 106224 133972 106276
rect 134024 106224 134030 106276
rect 157518 106264 157524 106276
rect 157479 106236 157524 106264
rect 157518 106224 157524 106236
rect 157576 106224 157582 106276
rect 179506 106264 179512 106276
rect 179467 106236 179512 106264
rect 179506 106224 179512 106236
rect 179564 106224 179570 106276
rect 133984 106140 134012 106224
rect 186148 106196 186176 106292
rect 220998 106264 221004 106276
rect 220959 106236 221004 106264
rect 220998 106224 221004 106236
rect 221056 106224 221062 106276
rect 244458 106224 244464 106276
rect 244516 106264 244522 106276
rect 244550 106264 244556 106276
rect 244516 106236 244556 106264
rect 244516 106224 244522 106236
rect 244550 106224 244556 106236
rect 244608 106224 244614 106276
rect 301958 106264 301964 106276
rect 301919 106236 301964 106264
rect 301958 106224 301964 106236
rect 302016 106224 302022 106276
rect 322658 106264 322664 106276
rect 322619 106236 322664 106264
rect 322658 106224 322664 106236
rect 322716 106224 322722 106276
rect 388714 106224 388720 106276
rect 388772 106264 388778 106276
rect 388806 106264 388812 106276
rect 388772 106236 388812 106264
rect 388772 106224 388778 106236
rect 388806 106224 388812 106236
rect 388864 106224 388870 106276
rect 394418 106264 394424 106276
rect 394379 106236 394424 106264
rect 394418 106224 394424 106236
rect 394476 106224 394482 106276
rect 420546 106224 420552 106276
rect 420604 106264 420610 106276
rect 420638 106264 420644 106276
rect 420604 106236 420644 106264
rect 420604 106224 420610 106236
rect 420638 106224 420644 106236
rect 420696 106224 420702 106276
rect 431586 106224 431592 106276
rect 431644 106264 431650 106276
rect 431678 106264 431684 106276
rect 431644 106236 431684 106264
rect 431644 106224 431650 106236
rect 431678 106224 431684 106236
rect 431736 106224 431742 106276
rect 186222 106196 186228 106208
rect 186148 106168 186228 106196
rect 186222 106156 186228 106168
rect 186280 106156 186286 106208
rect 133966 106088 133972 106140
rect 134024 106088 134030 106140
rect 227898 104972 227904 104984
rect 227824 104944 227904 104972
rect 227824 104916 227852 104944
rect 227898 104932 227904 104944
rect 227956 104932 227962 104984
rect 174170 104904 174176 104916
rect 174131 104876 174176 104904
rect 174170 104864 174176 104876
rect 174228 104864 174234 104916
rect 227806 104864 227812 104916
rect 227864 104864 227870 104916
rect 248322 104904 248328 104916
rect 248283 104876 248328 104904
rect 248322 104864 248328 104876
rect 248380 104864 248386 104916
rect 215386 104836 215392 104848
rect 215347 104808 215392 104836
rect 215386 104796 215392 104808
rect 215444 104796 215450 104848
rect 276106 104836 276112 104848
rect 276067 104808 276112 104836
rect 276106 104796 276112 104808
rect 276164 104796 276170 104848
rect 325694 104836 325700 104848
rect 325655 104808 325700 104836
rect 325694 104796 325700 104808
rect 325752 104796 325758 104848
rect 415026 104836 415032 104848
rect 414987 104808 415032 104836
rect 415026 104796 415032 104808
rect 415084 104796 415090 104848
rect 426250 104836 426256 104848
rect 426211 104808 426256 104836
rect 426250 104796 426256 104808
rect 426308 104796 426314 104848
rect 431586 104836 431592 104848
rect 431547 104808 431592 104836
rect 431586 104796 431592 104808
rect 431644 104796 431650 104848
rect 229186 103504 229192 103556
rect 229244 103544 229250 103556
rect 229281 103547 229339 103553
rect 229281 103544 229293 103547
rect 229244 103516 229293 103544
rect 229244 103504 229250 103516
rect 229281 103513 229293 103516
rect 229327 103513 229339 103547
rect 230382 103544 230388 103556
rect 230343 103516 230388 103544
rect 229281 103507 229339 103513
rect 230382 103504 230388 103516
rect 230440 103504 230446 103556
rect 186222 103476 186228 103488
rect 186183 103448 186228 103476
rect 186222 103436 186228 103448
rect 186280 103436 186286 103488
rect 233326 103476 233332 103488
rect 233287 103448 233332 103476
rect 233326 103436 233332 103448
rect 233384 103436 233390 103488
rect 279697 103479 279755 103485
rect 279697 103445 279709 103479
rect 279743 103476 279755 103479
rect 279786 103476 279792 103488
rect 279743 103448 279792 103476
rect 279743 103445 279755 103448
rect 279697 103439 279755 103445
rect 279786 103436 279792 103448
rect 279844 103436 279850 103488
rect 223666 102116 223672 102128
rect 223627 102088 223672 102116
rect 223666 102076 223672 102088
rect 223724 102076 223730 102128
rect 161382 101396 161388 101448
rect 161440 101436 161446 101448
rect 161750 101436 161756 101448
rect 161440 101408 161756 101436
rect 161440 101396 161446 101408
rect 161750 101396 161756 101408
rect 161808 101396 161814 101448
rect 222286 100688 222292 100700
rect 222247 100660 222292 100688
rect 222286 100648 222292 100660
rect 222344 100648 222350 100700
rect 240226 100076 240232 100088
rect 240187 100048 240232 100076
rect 240226 100036 240232 100048
rect 240284 100036 240290 100088
rect 248325 100079 248383 100085
rect 248325 100045 248337 100079
rect 248371 100076 248383 100079
rect 248414 100076 248420 100088
rect 248371 100048 248420 100076
rect 248371 100045 248383 100048
rect 248325 100039 248383 100045
rect 248414 100036 248420 100048
rect 248472 100036 248478 100088
rect 140958 99464 140964 99476
rect 140884 99436 140964 99464
rect 140884 99408 140912 99436
rect 140958 99424 140964 99436
rect 141016 99424 141022 99476
rect 208762 99464 208768 99476
rect 208596 99436 208768 99464
rect 208596 99408 208624 99436
rect 208762 99424 208768 99436
rect 208820 99424 208826 99476
rect 214190 99464 214196 99476
rect 214116 99436 214196 99464
rect 214116 99408 214144 99436
rect 214190 99424 214196 99436
rect 214248 99424 214254 99476
rect 232222 99464 232228 99476
rect 232148 99436 232228 99464
rect 232148 99408 232176 99436
rect 232222 99424 232228 99436
rect 232280 99424 232286 99476
rect 383286 99464 383292 99476
rect 383212 99436 383292 99464
rect 140866 99356 140872 99408
rect 140924 99356 140930 99408
rect 208578 99356 208584 99408
rect 208636 99356 208642 99408
rect 214098 99356 214104 99408
rect 214156 99356 214162 99408
rect 227806 99356 227812 99408
rect 227864 99356 227870 99408
rect 232130 99356 232136 99408
rect 232188 99356 232194 99408
rect 248506 99356 248512 99408
rect 248564 99356 248570 99408
rect 128906 99328 128912 99340
rect 128867 99300 128912 99328
rect 128906 99288 128912 99300
rect 128964 99288 128970 99340
rect 157521 99331 157579 99337
rect 157521 99297 157533 99331
rect 157567 99328 157579 99331
rect 157610 99328 157616 99340
rect 157567 99300 157616 99328
rect 157567 99297 157579 99300
rect 157521 99291 157579 99297
rect 157610 99288 157616 99300
rect 157668 99288 157674 99340
rect 179506 99328 179512 99340
rect 179467 99300 179512 99328
rect 179506 99288 179512 99300
rect 179564 99288 179570 99340
rect 227824 99328 227852 99356
rect 227898 99328 227904 99340
rect 227824 99300 227904 99328
rect 227898 99288 227904 99300
rect 227956 99288 227962 99340
rect 248414 99288 248420 99340
rect 248472 99328 248478 99340
rect 248524 99328 248552 99356
rect 383212 99340 383240 99436
rect 383286 99424 383292 99436
rect 383344 99424 383350 99476
rect 403894 99356 403900 99408
rect 403952 99356 403958 99408
rect 301958 99328 301964 99340
rect 248472 99300 248552 99328
rect 301919 99300 301964 99328
rect 248472 99288 248478 99300
rect 301958 99288 301964 99300
rect 302016 99288 302022 99340
rect 322658 99328 322664 99340
rect 322619 99300 322664 99328
rect 322658 99288 322664 99300
rect 322716 99288 322722 99340
rect 383194 99288 383200 99340
rect 383252 99288 383258 99340
rect 394418 99328 394424 99340
rect 394379 99300 394424 99328
rect 394418 99288 394424 99300
rect 394476 99288 394482 99340
rect 403912 99328 403940 99356
rect 403986 99328 403992 99340
rect 403912 99300 403992 99328
rect 403986 99288 403992 99300
rect 404044 99288 404050 99340
rect 173897 97223 173955 97229
rect 173897 97189 173909 97223
rect 173943 97220 173955 97223
rect 174170 97220 174176 97232
rect 173943 97192 174176 97220
rect 173943 97189 173955 97192
rect 173897 97183 173955 97189
rect 174170 97180 174176 97192
rect 174228 97180 174234 97232
rect 145006 96676 145012 96688
rect 144967 96648 145012 96676
rect 145006 96636 145012 96648
rect 145064 96636 145070 96688
rect 162946 96676 162952 96688
rect 162872 96648 162952 96676
rect 162872 96620 162900 96648
rect 162946 96636 162952 96648
rect 163004 96636 163010 96688
rect 220998 96676 221004 96688
rect 220959 96648 221004 96676
rect 220998 96636 221004 96648
rect 221056 96636 221062 96688
rect 128906 96568 128912 96620
rect 128964 96608 128970 96620
rect 128998 96608 129004 96620
rect 128964 96580 129004 96608
rect 128964 96568 128970 96580
rect 128998 96568 129004 96580
rect 129056 96568 129062 96620
rect 138014 96608 138020 96620
rect 137975 96580 138020 96608
rect 138014 96568 138020 96580
rect 138072 96568 138078 96620
rect 162854 96568 162860 96620
rect 162912 96568 162918 96620
rect 214098 96568 214104 96620
rect 214156 96608 214162 96620
rect 214282 96608 214288 96620
rect 214156 96580 214288 96608
rect 214156 96568 214162 96580
rect 214282 96568 214288 96580
rect 214340 96568 214346 96620
rect 216766 96608 216772 96620
rect 216727 96580 216772 96608
rect 216766 96568 216772 96580
rect 216824 96568 216830 96620
rect 290550 96608 290556 96620
rect 290511 96580 290556 96608
rect 290550 96568 290556 96580
rect 290608 96568 290614 96620
rect 341058 96568 341064 96620
rect 341116 96608 341122 96620
rect 341334 96608 341340 96620
rect 341116 96580 341340 96608
rect 341116 96568 341122 96580
rect 341334 96568 341340 96580
rect 341392 96568 341398 96620
rect 383105 96611 383163 96617
rect 383105 96577 383117 96611
rect 383151 96608 383163 96611
rect 383194 96608 383200 96620
rect 383151 96580 383200 96608
rect 383151 96577 383163 96580
rect 383105 96571 383163 96577
rect 383194 96568 383200 96580
rect 383252 96568 383258 96620
rect 388625 96611 388683 96617
rect 388625 96577 388637 96611
rect 388671 96608 388683 96611
rect 388714 96608 388720 96620
rect 388671 96580 388720 96608
rect 388671 96577 388683 96580
rect 388625 96571 388683 96577
rect 388714 96568 388720 96580
rect 388772 96568 388778 96620
rect 403897 96611 403955 96617
rect 403897 96577 403909 96611
rect 403943 96608 403955 96611
rect 403986 96608 403992 96620
rect 403943 96580 403992 96608
rect 403943 96577 403955 96580
rect 403897 96571 403955 96577
rect 403986 96568 403992 96580
rect 404044 96568 404050 96620
rect 420641 96611 420699 96617
rect 420641 96577 420653 96611
rect 420687 96608 420699 96611
rect 420730 96608 420736 96620
rect 420687 96580 420736 96608
rect 420687 96577 420699 96580
rect 420641 96571 420699 96577
rect 420730 96568 420736 96580
rect 420788 96568 420794 96620
rect 150618 95344 150624 95396
rect 150676 95384 150682 95396
rect 150802 95384 150808 95396
rect 150676 95356 150808 95384
rect 150676 95344 150682 95356
rect 150802 95344 150808 95356
rect 150860 95344 150866 95396
rect 426250 95316 426256 95328
rect 426211 95288 426256 95316
rect 426250 95276 426256 95288
rect 426308 95276 426314 95328
rect 173894 95248 173900 95260
rect 173855 95220 173900 95248
rect 173894 95208 173900 95220
rect 173952 95208 173958 95260
rect 215386 95248 215392 95260
rect 215347 95220 215392 95248
rect 215386 95208 215392 95220
rect 215444 95208 215450 95260
rect 240229 95251 240287 95257
rect 240229 95217 240241 95251
rect 240275 95248 240287 95251
rect 240318 95248 240324 95260
rect 240275 95220 240324 95248
rect 240275 95217 240287 95220
rect 240229 95211 240287 95217
rect 240318 95208 240324 95220
rect 240376 95208 240382 95260
rect 248322 95248 248328 95260
rect 248283 95220 248328 95248
rect 248322 95208 248328 95220
rect 248380 95208 248386 95260
rect 276106 95248 276112 95260
rect 276067 95220 276112 95248
rect 276106 95208 276112 95220
rect 276164 95208 276170 95260
rect 325694 95248 325700 95260
rect 325655 95220 325700 95248
rect 325694 95208 325700 95220
rect 325752 95208 325758 95260
rect 415029 95251 415087 95257
rect 415029 95217 415041 95251
rect 415075 95248 415087 95251
rect 415210 95248 415216 95260
rect 415075 95220 415216 95248
rect 415075 95217 415087 95220
rect 415029 95211 415087 95217
rect 415210 95208 415216 95220
rect 415268 95208 415274 95260
rect 140866 95180 140872 95192
rect 140827 95152 140872 95180
rect 140866 95140 140872 95152
rect 140924 95140 140930 95192
rect 150618 95180 150624 95192
rect 150579 95152 150624 95180
rect 150618 95140 150624 95152
rect 150676 95140 150682 95192
rect 162854 95140 162860 95192
rect 162912 95180 162918 95192
rect 271966 95180 271972 95192
rect 162912 95152 162957 95180
rect 271927 95152 271972 95180
rect 162912 95140 162918 95152
rect 271966 95140 271972 95152
rect 272024 95140 272030 95192
rect 229186 93916 229192 93968
rect 229244 93916 229250 93968
rect 186225 93891 186283 93897
rect 186225 93857 186237 93891
rect 186271 93888 186283 93891
rect 186314 93888 186320 93900
rect 186271 93860 186320 93888
rect 186271 93857 186283 93860
rect 186225 93851 186283 93857
rect 186314 93848 186320 93860
rect 186372 93848 186378 93900
rect 229204 93888 229232 93916
rect 229278 93888 229284 93900
rect 229204 93860 229284 93888
rect 229278 93848 229284 93860
rect 229336 93848 229342 93900
rect 233329 93891 233387 93897
rect 233329 93857 233341 93891
rect 233375 93888 233387 93891
rect 233418 93888 233424 93900
rect 233375 93860 233424 93888
rect 233375 93857 233387 93860
rect 233329 93851 233387 93857
rect 233418 93848 233424 93860
rect 233476 93848 233482 93900
rect 279694 93888 279700 93900
rect 279655 93860 279700 93888
rect 279694 93848 279700 93860
rect 279752 93848 279758 93900
rect 2774 93304 2780 93356
rect 2832 93344 2838 93356
rect 5350 93344 5356 93356
rect 2832 93316 5356 93344
rect 2832 93304 2838 93316
rect 5350 93304 5356 93316
rect 5408 93304 5414 93356
rect 161382 92964 161388 93016
rect 161440 93004 161446 93016
rect 161658 93004 161664 93016
rect 161440 92976 161664 93004
rect 161440 92964 161446 92976
rect 161658 92964 161664 92976
rect 161716 92964 161722 93016
rect 223669 92531 223727 92537
rect 223669 92497 223681 92531
rect 223715 92528 223727 92531
rect 223758 92528 223764 92540
rect 223715 92500 223764 92528
rect 223715 92497 223727 92500
rect 223669 92491 223727 92497
rect 223758 92488 223764 92500
rect 223816 92488 223822 92540
rect 227898 92460 227904 92472
rect 227859 92432 227904 92460
rect 227898 92420 227904 92432
rect 227956 92420 227962 92472
rect 207198 89768 207204 89820
rect 207256 89768 207262 89820
rect 415210 89808 415216 89820
rect 415136 89780 415216 89808
rect 126054 89700 126060 89752
rect 126112 89740 126118 89752
rect 126238 89740 126244 89752
rect 126112 89712 126244 89740
rect 126112 89700 126118 89712
rect 126238 89700 126244 89712
rect 126296 89700 126302 89752
rect 179414 89700 179420 89752
rect 179472 89740 179478 89752
rect 179598 89740 179604 89752
rect 179472 89712 179604 89740
rect 179472 89700 179478 89712
rect 179598 89700 179604 89712
rect 179656 89700 179662 89752
rect 183646 89700 183652 89752
rect 183704 89700 183710 89752
rect 190638 89700 190644 89752
rect 190696 89700 190702 89752
rect 192294 89700 192300 89752
rect 192352 89700 192358 89752
rect 138017 89675 138075 89681
rect 138017 89641 138029 89675
rect 138063 89672 138075 89675
rect 138106 89672 138112 89684
rect 138063 89644 138112 89672
rect 138063 89641 138075 89644
rect 138017 89635 138075 89641
rect 138106 89632 138112 89644
rect 138164 89632 138170 89684
rect 183664 89604 183692 89700
rect 183738 89604 183744 89616
rect 183664 89576 183744 89604
rect 183738 89564 183744 89576
rect 183796 89564 183802 89616
rect 190656 89604 190684 89700
rect 190730 89604 190736 89616
rect 190656 89576 190736 89604
rect 190730 89564 190736 89576
rect 190788 89564 190794 89616
rect 192312 89604 192340 89700
rect 207216 89684 207244 89768
rect 322566 89700 322572 89752
rect 322624 89740 322630 89752
rect 322750 89740 322756 89752
rect 322624 89712 322756 89740
rect 322624 89700 322630 89712
rect 322750 89700 322756 89712
rect 322808 89700 322814 89752
rect 394326 89700 394332 89752
rect 394384 89740 394390 89752
rect 394510 89740 394516 89752
rect 394384 89712 394516 89740
rect 394384 89700 394390 89712
rect 394510 89700 394516 89712
rect 394568 89700 394574 89752
rect 415136 89684 415164 89780
rect 415210 89768 415216 89780
rect 415268 89768 415274 89820
rect 207198 89632 207204 89684
rect 207256 89632 207262 89684
rect 415118 89632 415124 89684
rect 415176 89632 415182 89684
rect 192386 89604 192392 89616
rect 192312 89576 192392 89604
rect 192386 89564 192392 89576
rect 192444 89564 192450 89616
rect 234798 89564 234804 89616
rect 234856 89564 234862 89616
rect 216769 89539 216827 89545
rect 216769 89505 216781 89539
rect 216815 89536 216827 89539
rect 216858 89536 216864 89548
rect 216815 89508 216864 89536
rect 216815 89505 216827 89508
rect 216769 89499 216827 89505
rect 216858 89496 216864 89508
rect 216916 89496 216922 89548
rect 234816 89480 234844 89564
rect 234798 89428 234804 89480
rect 234856 89428 234862 89480
rect 290550 89400 290556 89412
rect 290511 89372 290556 89400
rect 290550 89360 290556 89372
rect 290608 89360 290614 89412
rect 131206 88272 131212 88324
rect 131264 88312 131270 88324
rect 580166 88312 580172 88324
rect 131264 88284 580172 88312
rect 131264 88272 131270 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 248598 86980 248604 87032
rect 248656 86980 248662 87032
rect 383102 87020 383108 87032
rect 383063 86992 383108 87020
rect 383102 86980 383108 86992
rect 383160 86980 383166 87032
rect 388622 87020 388628 87032
rect 388583 86992 388628 87020
rect 388622 86980 388628 86992
rect 388680 86980 388686 87032
rect 403894 87020 403900 87032
rect 403855 86992 403900 87020
rect 403894 86980 403900 86992
rect 403952 86980 403958 87032
rect 420638 87020 420644 87032
rect 420599 86992 420644 87020
rect 420638 86980 420644 86992
rect 420696 86980 420702 87032
rect 426161 87023 426219 87029
rect 426161 86989 426173 87023
rect 426207 87020 426219 87023
rect 426250 87020 426256 87032
rect 426207 86992 426256 87020
rect 426207 86989 426219 86992
rect 426161 86983 426219 86989
rect 426250 86980 426256 86992
rect 426308 86980 426314 87032
rect 431586 87020 431592 87032
rect 431547 86992 431592 87020
rect 431586 86980 431592 86992
rect 431644 86980 431650 87032
rect 128722 86912 128728 86964
rect 128780 86952 128786 86964
rect 128906 86952 128912 86964
rect 128780 86924 128912 86952
rect 128780 86912 128786 86924
rect 128906 86912 128912 86924
rect 128964 86912 128970 86964
rect 140869 86887 140927 86893
rect 140869 86853 140881 86887
rect 140915 86884 140927 86887
rect 140958 86884 140964 86896
rect 140915 86856 140964 86884
rect 140915 86853 140927 86856
rect 140869 86847 140927 86853
rect 140958 86844 140964 86856
rect 141016 86844 141022 86896
rect 162857 86887 162915 86893
rect 162857 86853 162869 86887
rect 162903 86884 162915 86887
rect 162946 86884 162952 86896
rect 162903 86856 162952 86884
rect 162903 86853 162915 86856
rect 162857 86847 162915 86853
rect 162946 86844 162952 86856
rect 163004 86844 163010 86896
rect 248616 86884 248644 86980
rect 290550 86952 290556 86964
rect 290511 86924 290556 86952
rect 290550 86912 290556 86924
rect 290608 86912 290614 86964
rect 322658 86952 322664 86964
rect 322619 86924 322664 86952
rect 322658 86912 322664 86924
rect 322716 86912 322722 86964
rect 394418 86952 394424 86964
rect 394379 86924 394424 86952
rect 394418 86912 394424 86924
rect 394476 86912 394482 86964
rect 248782 86884 248788 86896
rect 248616 86856 248788 86884
rect 248782 86844 248788 86856
rect 248840 86844 248846 86896
rect 150621 85595 150679 85601
rect 150621 85561 150633 85595
rect 150667 85592 150679 85595
rect 150710 85592 150716 85604
rect 150667 85564 150716 85592
rect 150667 85561 150679 85564
rect 150621 85555 150679 85561
rect 150710 85552 150716 85564
rect 150768 85552 150774 85604
rect 233326 85552 233332 85604
rect 233384 85592 233390 85604
rect 233510 85592 233516 85604
rect 233384 85564 233516 85592
rect 233384 85552 233390 85564
rect 233510 85552 233516 85564
rect 233568 85552 233574 85604
rect 271969 85595 272027 85601
rect 271969 85561 271981 85595
rect 272015 85592 272027 85595
rect 272058 85592 272064 85604
rect 272015 85564 272064 85592
rect 272015 85561 272027 85564
rect 271969 85555 272027 85561
rect 272058 85552 272064 85564
rect 272116 85552 272122 85604
rect 426158 85592 426164 85604
rect 426119 85564 426164 85592
rect 426158 85552 426164 85564
rect 426216 85552 426222 85604
rect 128633 85527 128691 85533
rect 128633 85493 128645 85527
rect 128679 85524 128691 85527
rect 128722 85524 128728 85536
rect 128679 85496 128728 85524
rect 128679 85493 128691 85496
rect 128633 85487 128691 85493
rect 128722 85484 128728 85496
rect 128780 85484 128786 85536
rect 147953 85527 148011 85533
rect 147953 85493 147965 85527
rect 147999 85524 148011 85527
rect 148134 85524 148140 85536
rect 147999 85496 148140 85524
rect 147999 85493 148011 85496
rect 147953 85487 148011 85493
rect 148134 85484 148140 85496
rect 148192 85484 148198 85536
rect 161658 85484 161664 85536
rect 161716 85524 161722 85536
rect 161750 85524 161756 85536
rect 161716 85496 161756 85524
rect 161716 85484 161722 85496
rect 161750 85484 161756 85496
rect 161808 85484 161814 85536
rect 214098 85524 214104 85536
rect 214059 85496 214104 85524
rect 214098 85484 214104 85496
rect 214156 85484 214162 85536
rect 325694 85524 325700 85536
rect 325655 85496 325700 85524
rect 325694 85484 325700 85496
rect 325752 85484 325758 85536
rect 140958 84164 140964 84176
rect 140919 84136 140964 84164
rect 140958 84124 140964 84136
rect 141016 84124 141022 84176
rect 192205 84167 192263 84173
rect 192205 84133 192217 84167
rect 192251 84164 192263 84167
rect 192386 84164 192392 84176
rect 192251 84136 192392 84164
rect 192251 84133 192263 84136
rect 192205 84127 192263 84133
rect 192386 84124 192392 84136
rect 192444 84124 192450 84176
rect 230382 84164 230388 84176
rect 230343 84136 230388 84164
rect 230382 84124 230388 84136
rect 230440 84124 230446 84176
rect 248417 84167 248475 84173
rect 248417 84133 248429 84167
rect 248463 84164 248475 84167
rect 248782 84164 248788 84176
rect 248463 84136 248788 84164
rect 248463 84133 248475 84136
rect 248417 84127 248475 84133
rect 248782 84124 248788 84136
rect 248840 84124 248846 84176
rect 279694 84164 279700 84176
rect 279655 84136 279700 84164
rect 279694 84124 279700 84136
rect 279752 84124 279758 84176
rect 426069 84167 426127 84173
rect 426069 84133 426081 84167
rect 426115 84164 426127 84167
rect 426158 84164 426164 84176
rect 426115 84136 426164 84164
rect 426115 84133 426127 84136
rect 426069 84127 426127 84133
rect 426158 84124 426164 84136
rect 426216 84124 426222 84176
rect 222289 82875 222347 82881
rect 222289 82841 222301 82875
rect 222335 82872 222347 82875
rect 222562 82872 222568 82884
rect 222335 82844 222568 82872
rect 222335 82841 222347 82844
rect 222289 82835 222347 82841
rect 222562 82832 222568 82844
rect 222620 82832 222626 82884
rect 227901 82875 227959 82881
rect 227901 82841 227913 82875
rect 227947 82872 227959 82875
rect 228082 82872 228088 82884
rect 227947 82844 228088 82872
rect 227947 82841 227959 82844
rect 227901 82835 227959 82841
rect 228082 82832 228088 82844
rect 228140 82832 228146 82884
rect 420270 82084 420276 82136
rect 420328 82124 420334 82136
rect 420638 82124 420644 82136
rect 420328 82096 420644 82124
rect 420328 82084 420334 82096
rect 420638 82084 420644 82096
rect 420696 82084 420702 82136
rect 207290 80832 207296 80844
rect 207251 80804 207296 80832
rect 207290 80792 207296 80804
rect 207348 80792 207354 80844
rect 271874 80724 271880 80776
rect 271932 80764 271938 80776
rect 272150 80764 272156 80776
rect 271932 80736 272156 80764
rect 271932 80724 271938 80736
rect 272150 80724 272156 80736
rect 272208 80724 272214 80776
rect 216858 80152 216864 80164
rect 216819 80124 216864 80152
rect 216858 80112 216864 80124
rect 216916 80112 216922 80164
rect 223669 80155 223727 80161
rect 223669 80121 223681 80155
rect 223715 80152 223727 80155
rect 223758 80152 223764 80164
rect 223715 80124 223764 80152
rect 223715 80121 223727 80124
rect 223669 80115 223727 80121
rect 223758 80112 223764 80124
rect 223816 80112 223822 80164
rect 229189 80155 229247 80161
rect 229189 80121 229201 80155
rect 229235 80152 229247 80155
rect 229278 80152 229284 80164
rect 229235 80124 229284 80152
rect 229235 80121 229247 80124
rect 229189 80115 229247 80121
rect 229278 80112 229284 80124
rect 229336 80112 229342 80164
rect 232130 80152 232136 80164
rect 232091 80124 232136 80152
rect 232130 80112 232136 80124
rect 232188 80112 232194 80164
rect 234798 80152 234804 80164
rect 234724 80124 234804 80152
rect 234724 80096 234752 80124
rect 234798 80112 234804 80124
rect 234856 80112 234862 80164
rect 240318 80152 240324 80164
rect 240244 80124 240324 80152
rect 240244 80096 240272 80124
rect 240318 80112 240324 80124
rect 240376 80112 240382 80164
rect 150526 80044 150532 80096
rect 150584 80084 150590 80096
rect 150710 80084 150716 80096
rect 150584 80056 150716 80084
rect 150584 80044 150590 80056
rect 150710 80044 150716 80056
rect 150768 80044 150774 80096
rect 234706 80044 234712 80096
rect 234764 80044 234770 80096
rect 240226 80044 240232 80096
rect 240284 80044 240290 80096
rect 431586 80044 431592 80096
rect 431644 80084 431650 80096
rect 431770 80084 431776 80096
rect 431644 80056 431776 80084
rect 431644 80044 431650 80056
rect 431770 80044 431776 80056
rect 431828 80044 431834 80096
rect 3234 79976 3240 80028
rect 3292 80016 3298 80028
rect 434990 80016 434996 80028
rect 3292 79988 434996 80016
rect 3292 79976 3298 79988
rect 434990 79976 434996 79988
rect 435048 79976 435054 80028
rect 216858 79948 216864 79960
rect 216819 79920 216864 79948
rect 216858 79908 216864 79920
rect 216916 79908 216922 79960
rect 232130 79948 232136 79960
rect 232091 79920 232136 79948
rect 232130 79908 232136 79920
rect 232188 79908 232194 79960
rect 290550 79948 290556 79960
rect 290511 79920 290556 79948
rect 290550 79908 290556 79920
rect 290608 79908 290614 79960
rect 301866 77324 301872 77376
rect 301924 77364 301930 77376
rect 302050 77364 302056 77376
rect 301924 77336 302056 77364
rect 301924 77324 301930 77336
rect 302050 77324 302056 77336
rect 302108 77324 302114 77376
rect 126238 77256 126244 77308
rect 126296 77296 126302 77308
rect 126330 77296 126336 77308
rect 126296 77268 126336 77296
rect 126296 77256 126302 77268
rect 126330 77256 126336 77268
rect 126388 77256 126394 77308
rect 207290 77296 207296 77308
rect 207251 77268 207296 77296
rect 207290 77256 207296 77268
rect 207348 77256 207354 77308
rect 245746 77256 245752 77308
rect 245804 77296 245810 77308
rect 245930 77296 245936 77308
rect 245804 77268 245936 77296
rect 245804 77256 245810 77268
rect 245930 77256 245936 77268
rect 245988 77256 245994 77308
rect 322661 77299 322719 77305
rect 322661 77265 322673 77299
rect 322707 77296 322719 77299
rect 322750 77296 322756 77308
rect 322707 77268 322756 77296
rect 322707 77265 322719 77268
rect 322661 77259 322719 77265
rect 322750 77256 322756 77268
rect 322808 77256 322814 77308
rect 394421 77299 394479 77305
rect 394421 77265 394433 77299
rect 394467 77296 394479 77299
rect 394510 77296 394516 77308
rect 394467 77268 394516 77296
rect 394467 77265 394479 77268
rect 394421 77259 394479 77265
rect 394510 77256 394516 77268
rect 394568 77256 394574 77308
rect 132126 77188 132132 77240
rect 132184 77228 132190 77240
rect 580166 77228 580172 77240
rect 132184 77200 580172 77228
rect 132184 77188 132190 77200
rect 580166 77188 580172 77200
rect 580224 77188 580230 77240
rect 301961 77163 302019 77169
rect 301961 77129 301973 77163
rect 302007 77160 302019 77163
rect 302050 77160 302056 77172
rect 302007 77132 302056 77160
rect 302007 77129 302019 77132
rect 301961 77123 302019 77129
rect 302050 77120 302056 77132
rect 302108 77120 302114 77172
rect 341334 77160 341340 77172
rect 341295 77132 341340 77160
rect 341334 77120 341340 77132
rect 341392 77120 341398 77172
rect 383194 77160 383200 77172
rect 383155 77132 383200 77160
rect 383194 77120 383200 77132
rect 383252 77120 383258 77172
rect 388714 77160 388720 77172
rect 388675 77132 388720 77160
rect 388714 77120 388720 77132
rect 388772 77120 388778 77172
rect 403986 77160 403992 77172
rect 403947 77132 403992 77160
rect 403986 77120 403992 77132
rect 404044 77120 404050 77172
rect 128630 75936 128636 75948
rect 128591 75908 128636 75936
rect 128630 75896 128636 75908
rect 128688 75896 128694 75948
rect 147950 75936 147956 75948
rect 147911 75908 147956 75936
rect 147950 75896 147956 75908
rect 148008 75896 148014 75948
rect 157334 75896 157340 75948
rect 157392 75936 157398 75948
rect 157702 75936 157708 75948
rect 157392 75908 157708 75936
rect 157392 75896 157398 75908
rect 157702 75896 157708 75908
rect 157760 75896 157766 75948
rect 183738 75896 183744 75948
rect 183796 75936 183802 75948
rect 183830 75936 183836 75948
rect 183796 75908 183836 75936
rect 183796 75896 183802 75908
rect 183830 75896 183836 75908
rect 183888 75896 183894 75948
rect 186222 75896 186228 75948
rect 186280 75936 186286 75948
rect 186314 75936 186320 75948
rect 186280 75908 186320 75936
rect 186280 75896 186286 75908
rect 186314 75896 186320 75908
rect 186372 75896 186378 75948
rect 190546 75896 190552 75948
rect 190604 75936 190610 75948
rect 190638 75936 190644 75948
rect 190604 75908 190644 75936
rect 190604 75896 190610 75908
rect 190638 75896 190644 75908
rect 190696 75896 190702 75948
rect 214098 75936 214104 75948
rect 214059 75908 214104 75936
rect 214098 75896 214104 75908
rect 214156 75896 214162 75948
rect 325694 75936 325700 75948
rect 325655 75908 325700 75936
rect 325694 75896 325700 75908
rect 325752 75896 325758 75948
rect 415026 75896 415032 75948
rect 415084 75936 415090 75948
rect 415118 75936 415124 75948
rect 415084 75908 415124 75936
rect 415084 75896 415090 75908
rect 415118 75896 415124 75908
rect 415176 75896 415182 75948
rect 244274 75868 244280 75880
rect 244235 75840 244280 75868
rect 244274 75828 244280 75840
rect 244332 75828 244338 75880
rect 245746 75868 245752 75880
rect 245707 75840 245752 75868
rect 245746 75828 245752 75840
rect 245804 75828 245810 75880
rect 271874 75868 271880 75880
rect 271835 75840 271880 75868
rect 271874 75828 271880 75840
rect 271932 75828 271938 75880
rect 431586 75868 431592 75880
rect 431547 75840 431592 75868
rect 431586 75828 431592 75840
rect 431644 75828 431650 75880
rect 140961 74579 141019 74585
rect 140961 74545 140973 74579
rect 141007 74576 141019 74579
rect 141050 74576 141056 74588
rect 141007 74548 141056 74576
rect 141007 74545 141019 74548
rect 140961 74539 141019 74545
rect 141050 74536 141056 74548
rect 141108 74536 141114 74588
rect 192202 74576 192208 74588
rect 192163 74548 192208 74576
rect 192202 74536 192208 74548
rect 192260 74536 192266 74588
rect 223666 74576 223672 74588
rect 223627 74548 223672 74576
rect 223666 74536 223672 74548
rect 223724 74536 223730 74588
rect 229186 74576 229192 74588
rect 229147 74548 229192 74576
rect 229186 74536 229192 74548
rect 229244 74536 229250 74588
rect 230382 74576 230388 74588
rect 230343 74548 230388 74576
rect 230382 74536 230388 74548
rect 230440 74536 230446 74588
rect 248414 74536 248420 74588
rect 248472 74576 248478 74588
rect 248472 74548 248517 74576
rect 248472 74536 248478 74548
rect 222378 73176 222384 73228
rect 222436 73216 222442 73228
rect 222470 73216 222476 73228
rect 222436 73188 222476 73216
rect 222436 73176 222442 73188
rect 222470 73176 222476 73188
rect 222528 73176 222534 73228
rect 227898 73176 227904 73228
rect 227956 73216 227962 73228
rect 227990 73216 227996 73228
rect 227956 73188 227996 73216
rect 227956 73176 227962 73188
rect 227990 73176 227996 73188
rect 228048 73176 228054 73228
rect 150710 70496 150716 70508
rect 150636 70468 150716 70496
rect 150636 70372 150664 70468
rect 150710 70456 150716 70468
rect 150768 70456 150774 70508
rect 179690 70496 179696 70508
rect 179616 70468 179696 70496
rect 179616 70372 179644 70468
rect 179690 70456 179696 70468
rect 179748 70456 179754 70508
rect 192202 70496 192208 70508
rect 192128 70468 192208 70496
rect 192128 70372 192156 70468
rect 192202 70456 192208 70468
rect 192260 70456 192266 70508
rect 150618 70320 150624 70372
rect 150676 70320 150682 70372
rect 179598 70320 179604 70372
rect 179656 70320 179662 70372
rect 192110 70320 192116 70372
rect 192168 70320 192174 70372
rect 245749 70363 245807 70369
rect 245749 70329 245761 70363
rect 245795 70360 245807 70363
rect 245838 70360 245844 70372
rect 245795 70332 245844 70360
rect 245795 70329 245807 70332
rect 245749 70323 245807 70329
rect 245838 70320 245844 70332
rect 245896 70320 245902 70372
rect 161750 70252 161756 70304
rect 161808 70252 161814 70304
rect 244277 70295 244335 70301
rect 244277 70261 244289 70295
rect 244323 70292 244335 70295
rect 244366 70292 244372 70304
rect 244323 70264 244372 70292
rect 244323 70261 244335 70264
rect 244277 70255 244335 70261
rect 244366 70252 244372 70264
rect 244424 70252 244430 70304
rect 161768 70168 161796 70252
rect 161750 70116 161756 70168
rect 161808 70116 161814 70168
rect 426066 69680 426072 69692
rect 426027 69652 426072 69680
rect 426066 69640 426072 69652
rect 426124 69640 426130 69692
rect 162946 67736 162952 67788
rect 163004 67736 163010 67788
rect 162964 67652 162992 67736
rect 145006 67600 145012 67652
rect 145064 67640 145070 67652
rect 145098 67640 145104 67652
rect 145064 67612 145104 67640
rect 145064 67600 145070 67612
rect 145098 67600 145104 67612
rect 145156 67600 145162 67652
rect 147950 67600 147956 67652
rect 148008 67640 148014 67652
rect 148042 67640 148048 67652
rect 148008 67612 148048 67640
rect 148008 67600 148014 67612
rect 148042 67600 148048 67612
rect 148100 67600 148106 67652
rect 162946 67600 162952 67652
rect 163004 67600 163010 67652
rect 173986 67600 173992 67652
rect 174044 67600 174050 67652
rect 301958 67640 301964 67652
rect 301919 67612 301964 67640
rect 301958 67600 301964 67612
rect 302016 67600 302022 67652
rect 341337 67643 341395 67649
rect 341337 67609 341349 67643
rect 341383 67640 341395 67643
rect 341426 67640 341432 67652
rect 341383 67612 341432 67640
rect 341383 67609 341395 67612
rect 341337 67603 341395 67609
rect 341426 67600 341432 67612
rect 341484 67600 341490 67652
rect 383197 67643 383255 67649
rect 383197 67609 383209 67643
rect 383243 67640 383255 67643
rect 383286 67640 383292 67652
rect 383243 67612 383292 67640
rect 383243 67609 383255 67612
rect 383197 67603 383255 67609
rect 383286 67600 383292 67612
rect 383344 67600 383350 67652
rect 388717 67643 388775 67649
rect 388717 67609 388729 67643
rect 388763 67640 388775 67643
rect 388806 67640 388812 67652
rect 388763 67612 388812 67640
rect 388763 67609 388775 67612
rect 388717 67603 388775 67609
rect 388806 67600 388812 67612
rect 388864 67600 388870 67652
rect 394418 67600 394424 67652
rect 394476 67640 394482 67652
rect 394510 67640 394516 67652
rect 394476 67612 394516 67640
rect 394476 67600 394482 67612
rect 394510 67600 394516 67612
rect 394568 67600 394574 67652
rect 403989 67643 404047 67649
rect 403989 67609 404001 67643
rect 404035 67640 404047 67643
rect 404078 67640 404084 67652
rect 404035 67612 404084 67640
rect 404035 67609 404047 67612
rect 403989 67603 404047 67609
rect 404078 67600 404084 67612
rect 404136 67600 404142 67652
rect 174004 67504 174032 67600
rect 216858 67572 216864 67584
rect 216819 67544 216864 67572
rect 216858 67532 216864 67544
rect 216916 67532 216922 67584
rect 238938 67572 238944 67584
rect 238899 67544 238944 67572
rect 238938 67532 238944 67544
rect 238996 67532 239002 67584
rect 174078 67504 174084 67516
rect 174004 67476 174084 67504
rect 174078 67464 174084 67476
rect 174136 67464 174142 67516
rect 271877 66283 271935 66289
rect 271877 66249 271889 66283
rect 271923 66280 271935 66283
rect 271966 66280 271972 66292
rect 271923 66252 271972 66280
rect 271923 66249 271935 66252
rect 271877 66243 271935 66249
rect 271966 66240 271972 66252
rect 272024 66240 272030 66292
rect 279697 66283 279755 66289
rect 279697 66249 279709 66283
rect 279743 66280 279755 66283
rect 279786 66280 279792 66292
rect 279743 66252 279792 66280
rect 279743 66249 279755 66252
rect 279697 66243 279755 66249
rect 279786 66240 279792 66252
rect 279844 66240 279850 66292
rect 322658 66240 322664 66292
rect 322716 66280 322722 66292
rect 322750 66280 322756 66292
rect 322716 66252 322756 66280
rect 322716 66240 322722 66252
rect 322750 66240 322756 66252
rect 322808 66240 322814 66292
rect 420454 66240 420460 66292
rect 420512 66280 420518 66292
rect 420546 66280 420552 66292
rect 420512 66252 420552 66280
rect 420512 66240 420518 66252
rect 420546 66240 420552 66252
rect 420604 66240 420610 66292
rect 431586 66280 431592 66292
rect 431547 66252 431592 66280
rect 431586 66240 431592 66252
rect 431644 66240 431650 66292
rect 128814 66212 128820 66224
rect 128775 66184 128820 66212
rect 128814 66172 128820 66184
rect 128872 66172 128878 66224
rect 162946 66212 162952 66224
rect 162907 66184 162952 66212
rect 162946 66172 162952 66184
rect 163004 66172 163010 66224
rect 214098 66172 214104 66224
rect 214156 66212 214162 66224
rect 214193 66215 214251 66221
rect 214193 66212 214205 66215
rect 214156 66184 214205 66212
rect 214156 66172 214162 66184
rect 214193 66181 214205 66184
rect 214239 66181 214251 66215
rect 214193 66175 214251 66181
rect 276106 66172 276112 66224
rect 276164 66212 276170 66224
rect 276290 66212 276296 66224
rect 276164 66184 276296 66212
rect 276164 66172 276170 66184
rect 276290 66172 276296 66184
rect 276348 66172 276354 66224
rect 325513 66215 325571 66221
rect 325513 66181 325525 66215
rect 325559 66212 325571 66215
rect 325694 66212 325700 66224
rect 325559 66184 325700 66212
rect 325559 66181 325571 66184
rect 325513 66175 325571 66181
rect 325694 66172 325700 66184
rect 325752 66172 325758 66224
rect 415026 66212 415032 66224
rect 414987 66184 415032 66212
rect 415026 66172 415032 66184
rect 415084 66172 415090 66224
rect 420454 66104 420460 66156
rect 420512 66144 420518 66156
rect 420638 66144 420644 66156
rect 420512 66116 420644 66144
rect 420512 66104 420518 66116
rect 420638 66104 420644 66116
rect 420696 66104 420702 66156
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 131666 64852 131672 64864
rect 3384 64824 131672 64852
rect 3384 64812 3390 64824
rect 131666 64812 131672 64824
rect 131724 64812 131730 64864
rect 144917 64855 144975 64861
rect 144917 64821 144929 64855
rect 144963 64852 144975 64855
rect 145006 64852 145012 64864
rect 144963 64824 145012 64852
rect 144963 64821 144975 64824
rect 144917 64815 144975 64821
rect 145006 64812 145012 64824
rect 145064 64812 145070 64864
rect 157334 64852 157340 64864
rect 157295 64824 157340 64852
rect 157334 64812 157340 64824
rect 157392 64812 157398 64864
rect 174078 64812 174084 64864
rect 174136 64852 174142 64864
rect 174262 64852 174268 64864
rect 174136 64824 174268 64852
rect 174136 64812 174142 64824
rect 174262 64812 174268 64824
rect 174320 64812 174326 64864
rect 290458 64852 290464 64864
rect 290419 64824 290464 64852
rect 290458 64812 290464 64824
rect 290516 64812 290522 64864
rect 436830 64812 436836 64864
rect 436888 64852 436894 64864
rect 579798 64852 579804 64864
rect 436888 64824 579804 64852
rect 436888 64812 436894 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 216858 61044 216864 61056
rect 216819 61016 216864 61044
rect 216858 61004 216864 61016
rect 216916 61004 216922 61056
rect 192110 60800 192116 60852
rect 192168 60800 192174 60852
rect 383286 60840 383292 60852
rect 383212 60812 383292 60840
rect 192128 60716 192156 60800
rect 383212 60716 383240 60812
rect 383286 60800 383292 60812
rect 383344 60800 383350 60852
rect 388806 60840 388812 60852
rect 388732 60812 388812 60840
rect 388732 60716 388760 60812
rect 388806 60800 388812 60812
rect 388864 60800 388870 60852
rect 404078 60840 404084 60852
rect 404004 60812 404084 60840
rect 404004 60716 404032 60812
rect 404078 60800 404084 60812
rect 404136 60800 404142 60852
rect 150526 60664 150532 60716
rect 150584 60704 150590 60716
rect 150710 60704 150716 60716
rect 150584 60676 150716 60704
rect 150584 60664 150590 60676
rect 150710 60664 150716 60676
rect 150768 60664 150774 60716
rect 161566 60664 161572 60716
rect 161624 60704 161630 60716
rect 161750 60704 161756 60716
rect 161624 60676 161756 60704
rect 161624 60664 161630 60676
rect 161750 60664 161756 60676
rect 161808 60664 161814 60716
rect 183646 60664 183652 60716
rect 183704 60704 183710 60716
rect 183830 60704 183836 60716
rect 183704 60676 183836 60704
rect 183704 60664 183710 60676
rect 183830 60664 183836 60676
rect 183888 60664 183894 60716
rect 190638 60664 190644 60716
rect 190696 60704 190702 60716
rect 190822 60704 190828 60716
rect 190696 60676 190828 60704
rect 190696 60664 190702 60676
rect 190822 60664 190828 60676
rect 190880 60664 190886 60716
rect 192110 60664 192116 60716
rect 192168 60664 192174 60716
rect 244366 60664 244372 60716
rect 244424 60704 244430 60716
rect 244550 60704 244556 60716
rect 244424 60676 244556 60704
rect 244424 60664 244430 60676
rect 244550 60664 244556 60676
rect 244608 60664 244614 60716
rect 245838 60664 245844 60716
rect 245896 60704 245902 60716
rect 246022 60704 246028 60716
rect 245896 60676 246028 60704
rect 245896 60664 245902 60676
rect 246022 60664 246028 60676
rect 246080 60664 246086 60716
rect 248414 60664 248420 60716
rect 248472 60704 248478 60716
rect 248598 60704 248604 60716
rect 248472 60676 248604 60704
rect 248472 60664 248478 60676
rect 248598 60664 248604 60676
rect 248656 60664 248662 60716
rect 271966 60664 271972 60716
rect 272024 60704 272030 60716
rect 272150 60704 272156 60716
rect 272024 60676 272156 60704
rect 272024 60664 272030 60676
rect 272150 60664 272156 60676
rect 272208 60664 272214 60716
rect 279878 60664 279884 60716
rect 279936 60704 279942 60716
rect 280062 60704 280068 60716
rect 279936 60676 280068 60704
rect 279936 60664 279942 60676
rect 280062 60664 280068 60676
rect 280120 60664 280126 60716
rect 383194 60664 383200 60716
rect 383252 60664 383258 60716
rect 388714 60664 388720 60716
rect 388772 60664 388778 60716
rect 403986 60664 403992 60716
rect 404044 60664 404050 60716
rect 220722 58624 220728 58676
rect 220780 58664 220786 58676
rect 220998 58664 221004 58676
rect 220780 58636 221004 58664
rect 220780 58624 220786 58636
rect 220998 58624 221004 58636
rect 221056 58624 221062 58676
rect 140866 57944 140872 57996
rect 140924 57984 140930 57996
rect 141050 57984 141056 57996
rect 140924 57956 141056 57984
rect 140924 57944 140930 57956
rect 141050 57944 141056 57956
rect 141108 57944 141114 57996
rect 186222 57944 186228 57996
rect 186280 57944 186286 57996
rect 238938 57984 238944 57996
rect 238899 57956 238944 57984
rect 238938 57944 238944 57956
rect 238996 57944 239002 57996
rect 186240 57916 186268 57944
rect 186314 57916 186320 57928
rect 186240 57888 186320 57916
rect 186314 57876 186320 57888
rect 186372 57876 186378 57928
rect 248230 57876 248236 57928
rect 248288 57916 248294 57928
rect 248322 57916 248328 57928
rect 248288 57888 248328 57916
rect 248288 57876 248294 57888
rect 248322 57876 248328 57888
rect 248380 57876 248386 57928
rect 280062 57916 280068 57928
rect 280023 57888 280068 57916
rect 280062 57876 280068 57888
rect 280120 57876 280126 57928
rect 301774 57916 301780 57928
rect 301735 57888 301780 57916
rect 301774 57876 301780 57888
rect 301832 57876 301838 57928
rect 322661 57919 322719 57925
rect 322661 57885 322673 57919
rect 322707 57916 322719 57919
rect 322750 57916 322756 57928
rect 322707 57888 322756 57916
rect 322707 57885 322719 57888
rect 322661 57879 322719 57885
rect 322750 57876 322756 57888
rect 322808 57876 322814 57928
rect 383194 57916 383200 57928
rect 383155 57888 383200 57916
rect 383194 57876 383200 57888
rect 383252 57876 383258 57928
rect 388714 57916 388720 57928
rect 388675 57888 388720 57916
rect 388714 57876 388720 57888
rect 388772 57876 388778 57928
rect 403986 57916 403992 57928
rect 403947 57888 403992 57916
rect 403986 57876 403992 57888
rect 404044 57876 404050 57928
rect 140866 57848 140872 57860
rect 140827 57820 140872 57848
rect 140866 57808 140872 57820
rect 140924 57808 140930 57860
rect 126238 56692 126244 56704
rect 125980 56664 126244 56692
rect 125980 56636 126008 56664
rect 126238 56652 126244 56664
rect 126296 56652 126302 56704
rect 125962 56584 125968 56636
rect 126020 56584 126026 56636
rect 128817 56627 128875 56633
rect 128817 56593 128829 56627
rect 128863 56624 128875 56627
rect 128906 56624 128912 56636
rect 128863 56596 128912 56624
rect 128863 56593 128875 56596
rect 128817 56587 128875 56593
rect 128906 56584 128912 56596
rect 128964 56584 128970 56636
rect 162946 56624 162952 56636
rect 162907 56596 162952 56624
rect 162946 56584 162952 56596
rect 163004 56584 163010 56636
rect 214098 56584 214104 56636
rect 214156 56624 214162 56636
rect 214193 56627 214251 56633
rect 214193 56624 214205 56627
rect 214156 56596 214205 56624
rect 214156 56584 214162 56596
rect 214193 56593 214205 56596
rect 214239 56593 214251 56627
rect 325510 56624 325516 56636
rect 325471 56596 325516 56624
rect 214193 56587 214251 56593
rect 325510 56584 325516 56596
rect 325568 56584 325574 56636
rect 415026 56624 415032 56636
rect 414987 56596 415032 56624
rect 415026 56584 415032 56596
rect 415084 56584 415090 56636
rect 179414 56556 179420 56568
rect 179375 56528 179420 56556
rect 179414 56516 179420 56528
rect 179472 56516 179478 56568
rect 192110 56556 192116 56568
rect 192071 56528 192116 56556
rect 192110 56516 192116 56528
rect 192168 56516 192174 56568
rect 207198 56516 207204 56568
rect 207256 56556 207262 56568
rect 207477 56559 207535 56565
rect 207477 56556 207489 56559
rect 207256 56528 207489 56556
rect 207256 56516 207262 56528
rect 207477 56525 207489 56528
rect 207523 56525 207535 56559
rect 207477 56519 207535 56525
rect 431586 56516 431592 56568
rect 431644 56556 431650 56568
rect 431770 56556 431776 56568
rect 431644 56528 431776 56556
rect 431644 56516 431650 56528
rect 431770 56516 431776 56528
rect 431828 56516 431834 56568
rect 144914 55264 144920 55276
rect 144875 55236 144920 55264
rect 144914 55224 144920 55236
rect 144972 55224 144978 55276
rect 157337 55267 157395 55273
rect 157337 55233 157349 55267
rect 157383 55264 157395 55267
rect 157426 55264 157432 55276
rect 157383 55236 157432 55264
rect 157383 55233 157395 55236
rect 157337 55227 157395 55233
rect 157426 55224 157432 55236
rect 157484 55224 157490 55276
rect 290461 55267 290519 55273
rect 290461 55233 290473 55267
rect 290507 55264 290519 55267
rect 290550 55264 290556 55276
rect 290507 55236 290556 55264
rect 290507 55233 290519 55236
rect 290461 55227 290519 55233
rect 290550 55224 290556 55236
rect 290608 55224 290614 55276
rect 186225 55199 186283 55205
rect 186225 55165 186237 55199
rect 186271 55196 186283 55199
rect 186314 55196 186320 55208
rect 186271 55168 186320 55196
rect 186271 55165 186283 55168
rect 186225 55159 186283 55165
rect 186314 55156 186320 55168
rect 186372 55156 186378 55208
rect 426066 53116 426072 53168
rect 426124 53156 426130 53168
rect 426250 53156 426256 53168
rect 426124 53128 426256 53156
rect 426124 53116 426130 53128
rect 426250 53116 426256 53128
rect 426308 53116 426314 53168
rect 157426 51756 157432 51808
rect 157484 51796 157490 51808
rect 157613 51799 157671 51805
rect 157613 51796 157625 51799
rect 157484 51768 157625 51796
rect 157484 51756 157490 51768
rect 157613 51765 157625 51768
rect 157659 51765 157671 51799
rect 157613 51759 157671 51765
rect 415026 51280 415032 51332
rect 415084 51320 415090 51332
rect 415210 51320 415216 51332
rect 415084 51292 415216 51320
rect 415084 51280 415090 51292
rect 415210 51280 415216 51292
rect 415268 51280 415274 51332
rect 223666 51144 223672 51196
rect 223724 51144 223730 51196
rect 229186 51144 229192 51196
rect 229244 51144 229250 51196
rect 290369 51187 290427 51193
rect 290369 51153 290381 51187
rect 290415 51184 290427 51187
rect 290550 51184 290556 51196
rect 290415 51156 290556 51184
rect 290415 51153 290427 51156
rect 290369 51147 290427 51153
rect 290550 51144 290556 51156
rect 290608 51144 290614 51196
rect 341518 51184 341524 51196
rect 341479 51156 341524 51184
rect 341518 51144 341524 51156
rect 341576 51144 341582 51196
rect 125962 51116 125968 51128
rect 125923 51088 125968 51116
rect 125962 51076 125968 51088
rect 126020 51076 126026 51128
rect 148042 51116 148048 51128
rect 147968 51088 148048 51116
rect 147968 51060 147996 51088
rect 148042 51076 148048 51088
rect 148100 51076 148106 51128
rect 161750 51076 161756 51128
rect 161808 51076 161814 51128
rect 128906 51008 128912 51060
rect 128964 51008 128970 51060
rect 147950 51008 147956 51060
rect 148008 51008 148014 51060
rect 128924 50980 128952 51008
rect 128998 50980 129004 50992
rect 128924 50952 129004 50980
rect 128998 50940 129004 50952
rect 129056 50940 129062 50992
rect 161768 50924 161796 51076
rect 223684 51060 223712 51144
rect 229204 51060 229232 51144
rect 272150 51116 272156 51128
rect 272076 51088 272156 51116
rect 272076 51060 272104 51088
rect 272150 51076 272156 51088
rect 272208 51076 272214 51128
rect 223666 51008 223672 51060
rect 223724 51008 223730 51060
rect 229186 51008 229192 51060
rect 229244 51008 229250 51060
rect 272058 51008 272064 51060
rect 272116 51008 272122 51060
rect 280062 51048 280068 51060
rect 280023 51020 280068 51048
rect 280062 51008 280068 51020
rect 280120 51008 280126 51060
rect 161750 50872 161756 50924
rect 161808 50872 161814 50924
rect 140869 48331 140927 48337
rect 140869 48297 140881 48331
rect 140915 48328 140927 48331
rect 140958 48328 140964 48340
rect 140915 48300 140964 48328
rect 140915 48297 140927 48300
rect 140869 48291 140927 48297
rect 140958 48288 140964 48300
rect 141016 48288 141022 48340
rect 162854 48288 162860 48340
rect 162912 48328 162918 48340
rect 162946 48328 162952 48340
rect 162912 48300 162952 48328
rect 162912 48288 162918 48300
rect 162946 48288 162952 48300
rect 163004 48288 163010 48340
rect 183830 48288 183836 48340
rect 183888 48328 183894 48340
rect 183922 48328 183928 48340
rect 183888 48300 183928 48328
rect 183888 48288 183894 48300
rect 183922 48288 183928 48300
rect 183980 48288 183986 48340
rect 301777 48331 301835 48337
rect 301777 48297 301789 48331
rect 301823 48328 301835 48331
rect 301866 48328 301872 48340
rect 301823 48300 301872 48328
rect 301823 48297 301835 48300
rect 301777 48291 301835 48297
rect 301866 48288 301872 48300
rect 301924 48288 301930 48340
rect 322658 48328 322664 48340
rect 322619 48300 322664 48328
rect 322658 48288 322664 48300
rect 322716 48288 322722 48340
rect 383197 48331 383255 48337
rect 383197 48297 383209 48331
rect 383243 48328 383255 48331
rect 383286 48328 383292 48340
rect 383243 48300 383292 48328
rect 383243 48297 383255 48300
rect 383197 48291 383255 48297
rect 383286 48288 383292 48300
rect 383344 48288 383350 48340
rect 388717 48331 388775 48337
rect 388717 48297 388729 48331
rect 388763 48328 388775 48331
rect 388806 48328 388812 48340
rect 388763 48300 388812 48328
rect 388763 48297 388775 48300
rect 388717 48291 388775 48297
rect 388806 48288 388812 48300
rect 388864 48288 388870 48340
rect 394418 48288 394424 48340
rect 394476 48328 394482 48340
rect 394510 48328 394516 48340
rect 394476 48300 394516 48328
rect 394476 48288 394482 48300
rect 394510 48288 394516 48300
rect 394568 48288 394574 48340
rect 403989 48331 404047 48337
rect 403989 48297 404001 48331
rect 404035 48328 404047 48331
rect 404078 48328 404084 48340
rect 404035 48300 404084 48328
rect 404035 48297 404047 48300
rect 403989 48291 404047 48297
rect 404078 48288 404084 48300
rect 404136 48288 404142 48340
rect 271877 48195 271935 48201
rect 271877 48161 271889 48195
rect 271923 48192 271935 48195
rect 272058 48192 272064 48204
rect 271923 48164 272064 48192
rect 271923 48161 271935 48164
rect 271877 48155 271935 48161
rect 272058 48152 272064 48164
rect 272116 48152 272122 48204
rect 290366 47036 290372 47048
rect 290327 47008 290372 47036
rect 290366 46996 290372 47008
rect 290424 46996 290430 47048
rect 125962 46968 125968 46980
rect 125923 46940 125968 46968
rect 125962 46928 125968 46940
rect 126020 46928 126026 46980
rect 179417 46971 179475 46977
rect 179417 46937 179429 46971
rect 179463 46968 179475 46971
rect 179506 46968 179512 46980
rect 179463 46940 179512 46968
rect 179463 46937 179475 46940
rect 179417 46931 179475 46937
rect 179506 46928 179512 46940
rect 179564 46928 179570 46980
rect 192110 46968 192116 46980
rect 192071 46940 192116 46968
rect 192110 46928 192116 46940
rect 192168 46928 192174 46980
rect 133322 46900 133328 46912
rect 133283 46872 133328 46900
rect 133322 46860 133328 46872
rect 133380 46860 133386 46912
rect 145006 46900 145012 46912
rect 144932 46872 145012 46900
rect 144932 46844 144960 46872
rect 145006 46860 145012 46872
rect 145064 46860 145070 46912
rect 147950 46900 147956 46912
rect 147876 46872 147956 46900
rect 147876 46844 147904 46872
rect 147950 46860 147956 46872
rect 148008 46860 148014 46912
rect 150621 46903 150679 46909
rect 150621 46869 150633 46903
rect 150667 46900 150679 46903
rect 150802 46900 150808 46912
rect 150667 46872 150808 46900
rect 150667 46869 150679 46872
rect 150621 46863 150679 46869
rect 150802 46860 150808 46872
rect 150860 46860 150866 46912
rect 162946 46900 162952 46912
rect 162907 46872 162952 46900
rect 162946 46860 162952 46872
rect 163004 46860 163010 46912
rect 214098 46900 214104 46912
rect 214059 46872 214104 46900
rect 214098 46860 214104 46872
rect 214156 46860 214162 46912
rect 215386 46900 215392 46912
rect 215347 46872 215392 46900
rect 215386 46860 215392 46872
rect 215444 46860 215450 46912
rect 248322 46900 248328 46912
rect 248283 46872 248328 46900
rect 248322 46860 248328 46872
rect 248380 46860 248386 46912
rect 276106 46860 276112 46912
rect 276164 46860 276170 46912
rect 290366 46860 290372 46912
rect 290424 46900 290430 46912
rect 290645 46903 290703 46909
rect 290645 46900 290657 46903
rect 290424 46872 290657 46900
rect 290424 46860 290430 46872
rect 290645 46869 290657 46872
rect 290691 46869 290703 46903
rect 325694 46900 325700 46912
rect 325655 46872 325700 46900
rect 290645 46863 290703 46869
rect 325694 46860 325700 46872
rect 325752 46860 325758 46912
rect 420454 46860 420460 46912
rect 420512 46900 420518 46912
rect 420638 46900 420644 46912
rect 420512 46872 420644 46900
rect 420512 46860 420518 46872
rect 420638 46860 420644 46872
rect 420696 46860 420702 46912
rect 425974 46900 425980 46912
rect 425935 46872 425980 46900
rect 425974 46860 425980 46872
rect 426032 46860 426038 46912
rect 431494 46860 431500 46912
rect 431552 46900 431558 46912
rect 431586 46900 431592 46912
rect 431552 46872 431592 46900
rect 431552 46860 431558 46872
rect 431586 46860 431592 46872
rect 431644 46860 431650 46912
rect 125962 46792 125968 46844
rect 126020 46832 126026 46844
rect 126146 46832 126152 46844
rect 126020 46804 126152 46832
rect 126020 46792 126026 46804
rect 126146 46792 126152 46804
rect 126204 46792 126210 46844
rect 144914 46792 144920 46844
rect 144972 46792 144978 46844
rect 147858 46792 147864 46844
rect 147916 46792 147922 46844
rect 276124 46773 276152 46860
rect 276109 46767 276167 46773
rect 276109 46733 276121 46767
rect 276155 46733 276167 46767
rect 276109 46727 276167 46733
rect 192110 45880 192116 45892
rect 192071 45852 192116 45880
rect 192110 45840 192116 45852
rect 192168 45840 192174 45892
rect 173986 45568 173992 45620
rect 174044 45608 174050 45620
rect 174262 45608 174268 45620
rect 174044 45580 174268 45608
rect 174044 45568 174050 45580
rect 174262 45568 174268 45580
rect 174320 45568 174326 45620
rect 186222 45608 186228 45620
rect 186183 45580 186228 45608
rect 186222 45568 186228 45580
rect 186280 45568 186286 45620
rect 341518 45608 341524 45620
rect 341479 45580 341524 45608
rect 341518 45568 341524 45580
rect 341576 45568 341582 45620
rect 183741 45543 183799 45549
rect 183741 45509 183753 45543
rect 183787 45540 183799 45543
rect 183922 45540 183928 45552
rect 183787 45512 183928 45540
rect 183787 45509 183799 45512
rect 183741 45503 183799 45509
rect 183922 45500 183928 45512
rect 183980 45500 183986 45552
rect 190641 45543 190699 45549
rect 190641 45509 190653 45543
rect 190687 45540 190699 45543
rect 190730 45540 190736 45552
rect 190687 45512 190736 45540
rect 190687 45509 190699 45512
rect 190641 45503 190699 45509
rect 190730 45500 190736 45512
rect 190788 45500 190794 45552
rect 414934 45540 414940 45552
rect 414895 45512 414940 45540
rect 414934 45500 414940 45512
rect 414992 45500 414998 45552
rect 341429 45475 341487 45481
rect 341429 45441 341441 45475
rect 341475 45472 341487 45475
rect 341518 45472 341524 45484
rect 341475 45444 341524 45472
rect 341475 45441 341487 45444
rect 341429 45435 341487 45441
rect 341518 45432 341524 45444
rect 341576 45432 341582 45484
rect 220998 44140 221004 44192
rect 221056 44180 221062 44192
rect 221182 44180 221188 44192
rect 221056 44152 221188 44180
rect 221056 44140 221062 44152
rect 221182 44140 221188 44152
rect 221240 44140 221246 44192
rect 248690 42032 248696 42084
rect 248748 42072 248754 42084
rect 248874 42072 248880 42084
rect 248748 42044 248880 42072
rect 248748 42032 248754 42044
rect 248874 42032 248880 42044
rect 248932 42032 248938 42084
rect 133598 41352 133604 41404
rect 133656 41392 133662 41404
rect 580166 41392 580172 41404
rect 133656 41364 580172 41392
rect 133656 41352 133662 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 192113 41327 192171 41333
rect 192113 41293 192125 41327
rect 192159 41324 192171 41327
rect 192202 41324 192208 41336
rect 192159 41296 192208 41324
rect 192159 41293 192171 41296
rect 192113 41287 192171 41293
rect 192202 41284 192208 41296
rect 192260 41284 192266 41336
rect 227898 41284 227904 41336
rect 227956 41324 227962 41336
rect 228174 41324 228180 41336
rect 227956 41296 228180 41324
rect 227956 41284 227962 41296
rect 228174 41284 228180 41296
rect 228232 41284 228238 41336
rect 271874 41324 271880 41336
rect 271835 41296 271880 41324
rect 271874 41284 271880 41296
rect 271932 41284 271938 41336
rect 173986 40712 173992 40724
rect 173947 40684 173992 40712
rect 173986 40672 173992 40684
rect 174044 40672 174050 40724
rect 186225 40715 186283 40721
rect 186225 40681 186237 40715
rect 186271 40712 186283 40715
rect 186314 40712 186320 40724
rect 186271 40684 186320 40712
rect 186271 40681 186283 40684
rect 186225 40675 186283 40681
rect 186314 40672 186320 40684
rect 186372 40672 186378 40724
rect 190638 40712 190644 40724
rect 190599 40684 190644 40712
rect 190638 40672 190644 40684
rect 190696 40672 190702 40724
rect 140866 38632 140872 38684
rect 140924 38672 140930 38684
rect 141050 38672 141056 38684
rect 140924 38644 141056 38672
rect 140924 38632 140930 38644
rect 141050 38632 141056 38644
rect 141108 38632 141114 38684
rect 157610 38672 157616 38684
rect 157571 38644 157616 38672
rect 157610 38632 157616 38644
rect 157668 38632 157674 38684
rect 207474 38672 207480 38684
rect 207435 38644 207480 38672
rect 207474 38632 207480 38644
rect 207532 38632 207538 38684
rect 244274 38632 244280 38684
rect 244332 38672 244338 38684
rect 244550 38672 244556 38684
rect 244332 38644 244556 38672
rect 244332 38632 244338 38644
rect 244550 38632 244556 38644
rect 244608 38632 244614 38684
rect 245746 38632 245752 38684
rect 245804 38672 245810 38684
rect 246022 38672 246028 38684
rect 245804 38644 246028 38672
rect 245804 38632 245810 38644
rect 246022 38632 246028 38644
rect 246080 38632 246086 38684
rect 279878 38632 279884 38684
rect 279936 38672 279942 38684
rect 280062 38672 280068 38684
rect 279936 38644 280068 38672
rect 279936 38632 279942 38644
rect 280062 38632 280068 38644
rect 280120 38632 280126 38684
rect 271874 38604 271880 38616
rect 271835 38576 271880 38604
rect 271874 38564 271880 38576
rect 271932 38564 271938 38616
rect 322661 38607 322719 38613
rect 322661 38573 322673 38607
rect 322707 38604 322719 38607
rect 322750 38604 322756 38616
rect 322707 38576 322756 38604
rect 322707 38573 322719 38576
rect 322661 38567 322719 38573
rect 322750 38564 322756 38576
rect 322808 38564 322814 38616
rect 383194 38604 383200 38616
rect 383155 38576 383200 38604
rect 383194 38564 383200 38576
rect 383252 38564 383258 38616
rect 403986 38604 403992 38616
rect 403947 38576 403992 38604
rect 403986 38564 403992 38576
rect 404044 38564 404050 38616
rect 290642 38536 290648 38548
rect 290603 38508 290648 38536
rect 290642 38496 290648 38508
rect 290700 38496 290706 38548
rect 341426 38264 341432 38276
rect 341387 38236 341432 38264
rect 341426 38224 341432 38236
rect 341484 38224 341490 38276
rect 133325 37315 133383 37321
rect 133325 37281 133337 37315
rect 133371 37312 133383 37315
rect 133506 37312 133512 37324
rect 133371 37284 133512 37312
rect 133371 37281 133383 37284
rect 133325 37275 133383 37281
rect 133506 37272 133512 37284
rect 133564 37272 133570 37324
rect 150618 37312 150624 37324
rect 150579 37284 150624 37312
rect 150618 37272 150624 37284
rect 150676 37272 150682 37324
rect 162946 37312 162952 37324
rect 162907 37284 162952 37312
rect 162946 37272 162952 37284
rect 163004 37272 163010 37324
rect 214098 37312 214104 37324
rect 214059 37284 214104 37312
rect 214098 37272 214104 37284
rect 214156 37272 214162 37324
rect 215386 37312 215392 37324
rect 215347 37284 215392 37312
rect 215386 37272 215392 37284
rect 215444 37272 215450 37324
rect 248322 37312 248328 37324
rect 248283 37284 248328 37312
rect 248322 37272 248328 37284
rect 248380 37272 248386 37324
rect 425977 37315 426035 37321
rect 425977 37281 425989 37315
rect 426023 37312 426035 37315
rect 426066 37312 426072 37324
rect 426023 37284 426072 37312
rect 426023 37281 426035 37284
rect 425977 37275 426035 37281
rect 426066 37272 426072 37284
rect 426124 37272 426130 37324
rect 179414 37244 179420 37256
rect 179375 37216 179420 37244
rect 179414 37204 179420 37216
rect 179472 37204 179478 37256
rect 244274 37244 244280 37256
rect 244235 37216 244280 37244
rect 244274 37204 244280 37216
rect 244332 37204 244338 37256
rect 245746 37244 245752 37256
rect 245707 37216 245752 37244
rect 245746 37204 245752 37216
rect 245804 37204 245810 37256
rect 431586 37244 431592 37256
rect 431547 37216 431592 37244
rect 431586 37204 431592 37216
rect 431644 37204 431650 37256
rect 414937 35955 414995 35961
rect 414937 35921 414949 35955
rect 414983 35952 414995 35955
rect 415026 35952 415032 35964
rect 414983 35924 415032 35952
rect 414983 35921 414995 35924
rect 414937 35915 414995 35921
rect 415026 35912 415032 35924
rect 415084 35912 415090 35964
rect 3418 35844 3424 35896
rect 3476 35884 3482 35896
rect 436186 35884 436192 35896
rect 3476 35856 436192 35884
rect 3476 35844 3482 35856
rect 436186 35844 436192 35856
rect 436244 35844 436250 35896
rect 227898 34416 227904 34468
rect 227956 34456 227962 34468
rect 227990 34456 227996 34468
rect 227956 34428 227996 34456
rect 227956 34416 227962 34428
rect 227990 34416 227996 34428
rect 228048 34416 228054 34468
rect 150618 33804 150624 33856
rect 150676 33844 150682 33856
rect 150802 33844 150808 33856
rect 150676 33816 150808 33844
rect 150676 33804 150682 33816
rect 150802 33804 150808 33816
rect 150860 33804 150866 33856
rect 223666 31872 223672 31884
rect 223592 31844 223672 31872
rect 128998 31804 129004 31816
rect 128924 31776 129004 31804
rect 128924 31748 128952 31776
rect 128998 31764 129004 31776
rect 129056 31764 129062 31816
rect 223592 31748 223620 31844
rect 223666 31832 223672 31844
rect 223724 31832 223730 31884
rect 301958 31832 301964 31884
rect 302016 31832 302022 31884
rect 290642 31764 290648 31816
rect 290700 31764 290706 31816
rect 128906 31696 128912 31748
rect 128964 31696 128970 31748
rect 192202 31736 192208 31748
rect 192163 31708 192208 31736
rect 192202 31696 192208 31708
rect 192260 31696 192266 31748
rect 223574 31696 223580 31748
rect 223632 31696 223638 31748
rect 279878 31696 279884 31748
rect 279936 31736 279942 31748
rect 280062 31736 280068 31748
rect 279936 31708 280068 31736
rect 279936 31696 279942 31708
rect 280062 31696 280068 31708
rect 280120 31696 280126 31748
rect 290660 31680 290688 31764
rect 301976 31736 302004 31832
rect 302050 31736 302056 31748
rect 301976 31708 302056 31736
rect 302050 31696 302056 31708
rect 302108 31696 302114 31748
rect 388714 31696 388720 31748
rect 388772 31736 388778 31748
rect 388898 31736 388904 31748
rect 388772 31708 388904 31736
rect 388772 31696 388778 31708
rect 388898 31696 388904 31708
rect 388956 31696 388962 31748
rect 244277 31671 244335 31677
rect 244277 31637 244289 31671
rect 244323 31668 244335 31671
rect 244366 31668 244372 31680
rect 244323 31640 244372 31668
rect 244323 31637 244335 31640
rect 244277 31631 244335 31637
rect 244366 31628 244372 31640
rect 244424 31628 244430 31680
rect 245749 31671 245807 31677
rect 245749 31637 245761 31671
rect 245795 31668 245807 31671
rect 245838 31668 245844 31680
rect 245795 31640 245844 31668
rect 245795 31637 245807 31640
rect 245749 31631 245807 31637
rect 245838 31628 245844 31640
rect 245896 31628 245902 31680
rect 290642 31628 290648 31680
rect 290700 31628 290706 31680
rect 341426 31628 341432 31680
rect 341484 31668 341490 31680
rect 341518 31668 341524 31680
rect 341484 31640 341524 31668
rect 341484 31628 341490 31640
rect 341518 31628 341524 31640
rect 341576 31628 341582 31680
rect 431589 31671 431647 31677
rect 431589 31637 431601 31671
rect 431635 31668 431647 31671
rect 431678 31668 431684 31680
rect 431635 31640 431684 31668
rect 431635 31637 431647 31640
rect 431589 31631 431647 31637
rect 431678 31628 431684 31640
rect 431736 31628 431742 31680
rect 132402 30268 132408 30320
rect 132460 30308 132466 30320
rect 580166 30308 580172 30320
rect 132460 30280 580172 30308
rect 132460 30268 132466 30280
rect 580166 30268 580172 30280
rect 580224 30268 580230 30320
rect 276106 29084 276112 29096
rect 276067 29056 276112 29084
rect 276106 29044 276112 29056
rect 276164 29044 276170 29096
rect 325694 29084 325700 29096
rect 325655 29056 325700 29084
rect 325694 29044 325700 29056
rect 325752 29044 325758 29096
rect 133322 28976 133328 29028
rect 133380 29016 133386 29028
rect 133506 29016 133512 29028
rect 133380 28988 133512 29016
rect 133380 28976 133386 28988
rect 133506 28976 133512 28988
rect 133564 28976 133570 29028
rect 161750 28976 161756 29028
rect 161808 29016 161814 29028
rect 161842 29016 161848 29028
rect 161808 28988 161848 29016
rect 161808 28976 161814 28988
rect 161842 28976 161848 28988
rect 161900 28976 161906 29028
rect 271877 29019 271935 29025
rect 271877 28985 271889 29019
rect 271923 29016 271935 29019
rect 271966 29016 271972 29028
rect 271923 28988 271972 29016
rect 271923 28985 271935 28988
rect 271877 28979 271935 28985
rect 271966 28976 271972 28988
rect 272024 28976 272030 29028
rect 322658 29016 322664 29028
rect 322619 28988 322664 29016
rect 322658 28976 322664 28988
rect 322716 28976 322722 29028
rect 383197 29019 383255 29025
rect 383197 28985 383209 29019
rect 383243 29016 383255 29019
rect 383286 29016 383292 29028
rect 383243 28988 383292 29016
rect 383243 28985 383255 28988
rect 383197 28979 383255 28985
rect 383286 28976 383292 28988
rect 383344 28976 383350 29028
rect 394418 28976 394424 29028
rect 394476 29016 394482 29028
rect 394510 29016 394516 29028
rect 394476 28988 394516 29016
rect 394476 28976 394482 28988
rect 394510 28976 394516 28988
rect 394568 28976 394574 29028
rect 403989 29019 404047 29025
rect 403989 28985 404001 29019
rect 404035 29016 404047 29019
rect 404078 29016 404084 29028
rect 404035 28988 404084 29016
rect 404035 28985 404047 28988
rect 403989 28979 404047 28985
rect 404078 28976 404084 28988
rect 404136 28976 404142 29028
rect 128906 28908 128912 28960
rect 128964 28908 128970 28960
rect 140869 28951 140927 28957
rect 140869 28917 140881 28951
rect 140915 28948 140927 28951
rect 140958 28948 140964 28960
rect 140915 28920 140964 28948
rect 140915 28917 140927 28920
rect 140869 28911 140927 28917
rect 140958 28908 140964 28920
rect 141016 28908 141022 28960
rect 207474 28948 207480 28960
rect 207435 28920 207480 28948
rect 207474 28908 207480 28920
rect 207532 28908 207538 28960
rect 279973 28951 280031 28957
rect 279973 28917 279985 28951
rect 280019 28948 280031 28951
rect 280062 28948 280068 28960
rect 280019 28920 280068 28948
rect 280019 28917 280031 28920
rect 279973 28911 280031 28917
rect 280062 28908 280068 28920
rect 280120 28908 280126 28960
rect 128924 28880 128952 28908
rect 128998 28880 129004 28892
rect 128924 28852 129004 28880
rect 128998 28840 129004 28852
rect 129056 28840 129062 28892
rect 179417 27659 179475 27665
rect 179417 27625 179429 27659
rect 179463 27656 179475 27659
rect 179506 27656 179512 27668
rect 179463 27628 179512 27656
rect 179463 27625 179475 27628
rect 179417 27619 179475 27625
rect 179506 27616 179512 27628
rect 179564 27616 179570 27668
rect 183738 27656 183744 27668
rect 183699 27628 183744 27656
rect 183738 27616 183744 27628
rect 183796 27616 183802 27668
rect 248506 27616 248512 27668
rect 248564 27656 248570 27668
rect 248690 27656 248696 27668
rect 248564 27628 248696 27656
rect 248564 27616 248570 27628
rect 248690 27616 248696 27628
rect 248748 27616 248754 27668
rect 125965 27591 126023 27597
rect 125965 27557 125977 27591
rect 126011 27588 126023 27591
rect 126054 27588 126060 27600
rect 126011 27560 126060 27588
rect 126011 27557 126023 27560
rect 125965 27551 126023 27557
rect 126054 27548 126060 27560
rect 126112 27548 126118 27600
rect 133322 27588 133328 27600
rect 133283 27560 133328 27588
rect 133322 27548 133328 27560
rect 133380 27548 133386 27600
rect 162946 27588 162952 27600
rect 162907 27560 162952 27588
rect 162946 27548 162952 27560
rect 163004 27548 163010 27600
rect 190457 27591 190515 27597
rect 190457 27557 190469 27591
rect 190503 27588 190515 27591
rect 190638 27588 190644 27600
rect 190503 27560 190644 27588
rect 190503 27557 190515 27560
rect 190457 27551 190515 27557
rect 190638 27548 190644 27560
rect 190696 27548 190702 27600
rect 192202 27588 192208 27600
rect 192163 27560 192208 27588
rect 192202 27548 192208 27560
rect 192260 27548 192266 27600
rect 214098 27588 214104 27600
rect 214059 27560 214104 27588
rect 214098 27548 214104 27560
rect 214156 27548 214162 27600
rect 215386 27588 215392 27600
rect 215347 27560 215392 27588
rect 215386 27548 215392 27560
rect 215444 27548 215450 27600
rect 276106 27588 276112 27600
rect 276067 27560 276112 27588
rect 276106 27548 276112 27560
rect 276164 27548 276170 27600
rect 325694 27588 325700 27600
rect 325655 27560 325700 27588
rect 325694 27548 325700 27560
rect 325752 27548 325758 27600
rect 420454 27588 420460 27600
rect 420415 27560 420460 27588
rect 420454 27548 420460 27560
rect 420512 27548 420518 27600
rect 186222 27112 186228 27124
rect 186183 27084 186228 27112
rect 186222 27072 186228 27084
rect 186280 27072 186286 27124
rect 173989 26299 174047 26305
rect 173989 26265 174001 26299
rect 174035 26296 174047 26299
rect 174078 26296 174084 26308
rect 174035 26268 174084 26296
rect 174035 26265 174047 26268
rect 173989 26259 174047 26265
rect 174078 26256 174084 26268
rect 174136 26256 174142 26308
rect 183738 26228 183744 26240
rect 183699 26200 183744 26228
rect 183738 26188 183744 26200
rect 183796 26188 183802 26240
rect 192202 26188 192208 26240
rect 192260 26228 192266 26240
rect 301866 26228 301872 26240
rect 192260 26200 192305 26228
rect 301827 26200 301872 26228
rect 192260 26188 192266 26200
rect 301866 26188 301872 26200
rect 301924 26188 301930 26240
rect 415026 26228 415032 26240
rect 414987 26200 415032 26228
rect 415026 26188 415032 26200
rect 415084 26188 415090 26240
rect 431497 26231 431555 26237
rect 431497 26197 431509 26231
rect 431543 26228 431555 26231
rect 431678 26228 431684 26240
rect 431543 26200 431684 26228
rect 431543 26197 431555 26200
rect 431497 26191 431555 26197
rect 431678 26188 431684 26200
rect 431736 26188 431742 26240
rect 383378 25276 383384 25288
rect 383339 25248 383384 25276
rect 383378 25236 383384 25248
rect 383436 25236 383442 25288
rect 222289 24939 222347 24945
rect 222289 24905 222301 24939
rect 222335 24936 222347 24939
rect 222378 24936 222384 24948
rect 222335 24908 222384 24936
rect 222335 24905 222347 24908
rect 222289 24899 222347 24905
rect 222378 24896 222384 24908
rect 222436 24896 222442 24948
rect 220998 24828 221004 24880
rect 221056 24868 221062 24880
rect 221182 24868 221188 24880
rect 221056 24840 221188 24868
rect 221056 24828 221062 24840
rect 221182 24828 221188 24840
rect 221240 24828 221246 24880
rect 230109 24803 230167 24809
rect 230109 24769 230121 24803
rect 230155 24800 230167 24803
rect 230382 24800 230388 24812
rect 230155 24772 230388 24800
rect 230155 24769 230167 24772
rect 230109 24763 230167 24769
rect 230382 24760 230388 24772
rect 230440 24760 230446 24812
rect 147858 24148 147864 24200
rect 147916 24188 147922 24200
rect 148042 24188 148048 24200
rect 147916 24160 148048 24188
rect 147916 24148 147922 24160
rect 148042 24148 148048 24160
rect 148100 24148 148106 24200
rect 388714 24148 388720 24200
rect 388772 24188 388778 24200
rect 388898 24188 388904 24200
rect 388772 24160 388904 24188
rect 388772 24148 388778 24160
rect 388898 24148 388904 24160
rect 388956 24148 388962 24200
rect 222286 23508 222292 23520
rect 222247 23480 222292 23508
rect 222286 23468 222292 23480
rect 222344 23468 222350 23520
rect 161750 22760 161756 22772
rect 161711 22732 161756 22760
rect 161750 22720 161756 22732
rect 161808 22720 161814 22772
rect 238938 22216 238944 22228
rect 238899 22188 238944 22216
rect 238938 22176 238944 22188
rect 238996 22176 239002 22228
rect 174078 22108 174084 22160
rect 174136 22108 174142 22160
rect 404078 22148 404084 22160
rect 404004 22120 404084 22148
rect 3142 22040 3148 22092
rect 3200 22080 3206 22092
rect 132218 22080 132224 22092
rect 3200 22052 132224 22080
rect 3200 22040 3206 22052
rect 132218 22040 132224 22052
rect 132276 22040 132282 22092
rect 144914 22040 144920 22092
rect 144972 22080 144978 22092
rect 145098 22080 145104 22092
rect 144972 22052 145104 22080
rect 144972 22040 144978 22052
rect 145098 22040 145104 22052
rect 145156 22040 145162 22092
rect 174096 22024 174124 22108
rect 404004 22092 404032 22120
rect 404078 22108 404084 22120
rect 404136 22108 404142 22160
rect 244366 22040 244372 22092
rect 244424 22080 244430 22092
rect 244550 22080 244556 22092
rect 244424 22052 244556 22080
rect 244424 22040 244430 22052
rect 244550 22040 244556 22052
rect 244608 22040 244614 22092
rect 245838 22040 245844 22092
rect 245896 22080 245902 22092
rect 246022 22080 246028 22092
rect 245896 22052 246028 22080
rect 245896 22040 245902 22052
rect 246022 22040 246028 22052
rect 246080 22040 246086 22092
rect 248414 22040 248420 22092
rect 248472 22080 248478 22092
rect 248598 22080 248604 22092
rect 248472 22052 248604 22080
rect 248472 22040 248478 22052
rect 248598 22040 248604 22052
rect 248656 22040 248662 22092
rect 290734 22040 290740 22092
rect 290792 22080 290798 22092
rect 290918 22080 290924 22092
rect 290792 22052 290924 22080
rect 290792 22040 290798 22052
rect 290918 22040 290924 22052
rect 290976 22040 290982 22092
rect 403986 22040 403992 22092
rect 404044 22040 404050 22092
rect 174078 21972 174084 22024
rect 174136 21972 174142 22024
rect 220998 20068 221004 20120
rect 221056 20068 221062 20120
rect 221016 19984 221044 20068
rect 227809 20043 227867 20049
rect 227809 20009 227821 20043
rect 227855 20040 227867 20043
rect 227990 20040 227996 20052
rect 227855 20012 227996 20040
rect 227855 20009 227867 20012
rect 227809 20003 227867 20009
rect 227990 20000 227996 20012
rect 228048 20000 228054 20052
rect 220998 19932 221004 19984
rect 221056 19932 221062 19984
rect 140866 19428 140872 19440
rect 140827 19400 140872 19428
rect 140866 19388 140872 19400
rect 140924 19388 140930 19440
rect 207198 19388 207204 19440
rect 207256 19428 207262 19440
rect 207477 19431 207535 19437
rect 207477 19428 207489 19431
rect 207256 19400 207489 19428
rect 207256 19388 207262 19400
rect 207477 19397 207489 19400
rect 207523 19397 207535 19431
rect 207477 19391 207535 19397
rect 150618 19320 150624 19372
rect 150676 19360 150682 19372
rect 150710 19360 150716 19372
rect 150676 19332 150716 19360
rect 150676 19320 150682 19332
rect 150710 19320 150716 19332
rect 150768 19320 150774 19372
rect 238938 19360 238944 19372
rect 238899 19332 238944 19360
rect 238938 19320 238944 19332
rect 238996 19320 239002 19372
rect 279970 19360 279976 19372
rect 279931 19332 279976 19360
rect 279970 19320 279976 19332
rect 280028 19320 280034 19372
rect 383378 19360 383384 19372
rect 383339 19332 383384 19360
rect 383378 19320 383384 19332
rect 383436 19320 383442 19372
rect 133322 19292 133328 19304
rect 133283 19264 133328 19292
rect 133322 19252 133328 19264
rect 133380 19252 133386 19304
rect 140866 19292 140872 19304
rect 140827 19264 140872 19292
rect 140866 19252 140872 19264
rect 140924 19252 140930 19304
rect 179690 19292 179696 19304
rect 179651 19264 179696 19292
rect 179690 19252 179696 19264
rect 179748 19252 179754 19304
rect 207201 19295 207259 19301
rect 207201 19261 207213 19295
rect 207247 19292 207259 19295
rect 207290 19292 207296 19304
rect 207247 19264 207296 19292
rect 207247 19261 207259 19264
rect 207201 19255 207259 19261
rect 207290 19252 207296 19264
rect 207348 19252 207354 19304
rect 238389 19295 238447 19301
rect 238389 19261 238401 19295
rect 238435 19292 238447 19295
rect 238662 19292 238668 19304
rect 238435 19264 238668 19292
rect 238435 19261 238447 19264
rect 238389 19255 238447 19261
rect 238662 19252 238668 19264
rect 238720 19252 238726 19304
rect 290918 19292 290924 19304
rect 290879 19264 290924 19292
rect 290918 19252 290924 19264
rect 290976 19252 290982 19304
rect 425974 19252 425980 19304
rect 426032 19292 426038 19304
rect 426066 19292 426072 19304
rect 426032 19264 426072 19292
rect 426032 19252 426038 19264
rect 426066 19252 426072 19264
rect 426124 19252 426130 19304
rect 162946 18000 162952 18012
rect 162907 17972 162952 18000
rect 162946 17960 162952 17972
rect 163004 17960 163010 18012
rect 190454 18000 190460 18012
rect 190415 17972 190460 18000
rect 190454 17960 190460 17972
rect 190512 17960 190518 18012
rect 276106 18000 276112 18012
rect 276067 17972 276112 18000
rect 276106 17960 276112 17972
rect 276164 17960 276170 18012
rect 420457 18003 420515 18009
rect 420457 17969 420469 18003
rect 420503 18000 420515 18003
rect 420546 18000 420552 18012
rect 420503 17972 420552 18000
rect 420503 17969 420515 17972
rect 420457 17963 420515 17969
rect 420546 17960 420552 17972
rect 420604 17960 420610 18012
rect 436738 17892 436744 17944
rect 436796 17932 436802 17944
rect 579798 17932 579804 17944
rect 436796 17904 579804 17932
rect 436796 17892 436802 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 183741 16643 183799 16649
rect 183741 16609 183753 16643
rect 183787 16640 183799 16643
rect 183830 16640 183836 16652
rect 183787 16612 183836 16640
rect 183787 16609 183799 16612
rect 183741 16603 183799 16609
rect 183830 16600 183836 16612
rect 183888 16600 183894 16652
rect 192202 16640 192208 16652
rect 192163 16612 192208 16640
rect 192202 16600 192208 16612
rect 192260 16600 192266 16652
rect 415026 16640 415032 16652
rect 414987 16612 415032 16640
rect 415026 16600 415032 16612
rect 415084 16600 415090 16652
rect 431494 16640 431500 16652
rect 431455 16612 431500 16640
rect 431494 16600 431500 16612
rect 431552 16600 431558 16652
rect 274818 15892 274824 15904
rect 274779 15864 274824 15892
rect 274818 15852 274824 15864
rect 274876 15852 274882 15904
rect 222286 15172 222292 15224
rect 222344 15172 222350 15224
rect 222304 15144 222332 15172
rect 222378 15144 222384 15156
rect 222304 15116 222384 15144
rect 222378 15104 222384 15116
rect 222436 15104 222442 15156
rect 237282 12560 237288 12572
rect 237116 12532 237288 12560
rect 162946 12492 162952 12504
rect 162872 12464 162952 12492
rect 162872 12436 162900 12464
rect 162946 12452 162952 12464
rect 163004 12452 163010 12504
rect 168377 12495 168435 12501
rect 168377 12461 168389 12495
rect 168423 12492 168435 12495
rect 168466 12492 168472 12504
rect 168423 12464 168472 12492
rect 168423 12461 168435 12464
rect 168377 12455 168435 12461
rect 168466 12452 168472 12464
rect 168524 12452 168530 12504
rect 186222 12492 186228 12504
rect 186056 12464 186228 12492
rect 186056 12436 186084 12464
rect 186222 12452 186228 12464
rect 186280 12452 186286 12504
rect 208394 12452 208400 12504
rect 208452 12492 208458 12504
rect 208578 12492 208584 12504
rect 208452 12464 208584 12492
rect 208452 12452 208458 12464
rect 208578 12452 208584 12464
rect 208636 12452 208642 12504
rect 237116 12436 237144 12532
rect 237282 12520 237288 12532
rect 237340 12520 237346 12572
rect 383286 12560 383292 12572
rect 383247 12532 383292 12560
rect 383286 12520 383292 12532
rect 383344 12520 383350 12572
rect 237190 12452 237196 12504
rect 237248 12452 237254 12504
rect 248322 12492 248328 12504
rect 247972 12464 248328 12492
rect 162854 12384 162860 12436
rect 162912 12384 162918 12436
rect 186038 12384 186044 12436
rect 186096 12384 186102 12436
rect 237098 12384 237104 12436
rect 237156 12384 237162 12436
rect 237208 12368 237236 12452
rect 247972 12436 248000 12464
rect 248322 12452 248328 12464
rect 248380 12452 248386 12504
rect 276106 12452 276112 12504
rect 276164 12452 276170 12504
rect 394326 12452 394332 12504
rect 394384 12452 394390 12504
rect 415026 12492 415032 12504
rect 414952 12464 415032 12492
rect 247954 12384 247960 12436
rect 248012 12384 248018 12436
rect 237190 12316 237196 12368
rect 237248 12316 237254 12368
rect 276124 12356 276152 12452
rect 321738 12384 321744 12436
rect 321796 12384 321802 12436
rect 276474 12356 276480 12368
rect 276124 12328 276480 12356
rect 276474 12316 276480 12328
rect 276532 12316 276538 12368
rect 321756 12356 321784 12384
rect 322750 12356 322756 12368
rect 321756 12328 322756 12356
rect 322750 12316 322756 12328
rect 322808 12316 322814 12368
rect 394344 12356 394372 12452
rect 414952 12436 414980 12464
rect 415026 12452 415032 12464
rect 415084 12452 415090 12504
rect 420546 12492 420552 12504
rect 420472 12464 420552 12492
rect 420472 12436 420500 12464
rect 420546 12452 420552 12464
rect 420604 12452 420610 12504
rect 414934 12384 414940 12436
rect 414992 12384 414998 12436
rect 420454 12384 420460 12436
rect 420512 12384 420518 12436
rect 463694 12384 463700 12436
rect 463752 12424 463758 12436
rect 464338 12424 464344 12436
rect 463752 12396 464344 12424
rect 463752 12384 463758 12396
rect 464338 12384 464344 12396
rect 464396 12384 464402 12436
rect 394418 12356 394424 12368
rect 394344 12328 394424 12356
rect 394418 12316 394424 12328
rect 394476 12316 394482 12368
rect 161750 11880 161756 11892
rect 161711 11852 161756 11880
rect 161750 11840 161756 11852
rect 161808 11840 161814 11892
rect 371050 10684 371056 10736
rect 371108 10724 371114 10736
rect 459646 10724 459652 10736
rect 371108 10696 459652 10724
rect 371108 10684 371114 10696
rect 459646 10684 459652 10696
rect 459704 10684 459710 10736
rect 372338 10616 372344 10668
rect 372396 10656 372402 10668
rect 463234 10656 463240 10668
rect 372396 10628 463240 10656
rect 372396 10616 372402 10628
rect 463234 10616 463240 10628
rect 463292 10616 463298 10668
rect 375190 10548 375196 10600
rect 375248 10588 375254 10600
rect 466822 10588 466828 10600
rect 375248 10560 466828 10588
rect 375248 10548 375254 10560
rect 466822 10548 466828 10560
rect 466880 10548 466886 10600
rect 376570 10480 376576 10532
rect 376628 10520 376634 10532
rect 470318 10520 470324 10532
rect 376628 10492 470324 10520
rect 376628 10480 376634 10492
rect 470318 10480 470324 10492
rect 470376 10480 470382 10532
rect 377950 10412 377956 10464
rect 378008 10452 378014 10464
rect 473354 10452 473360 10464
rect 378008 10424 473360 10452
rect 378008 10412 378014 10424
rect 473354 10412 473360 10424
rect 473412 10412 473418 10464
rect 380802 10344 380808 10396
rect 380860 10384 380866 10396
rect 477678 10384 477684 10396
rect 380860 10356 477684 10384
rect 380860 10344 380866 10356
rect 477678 10344 477684 10356
rect 477736 10344 477742 10396
rect 382090 10276 382096 10328
rect 382148 10316 382154 10328
rect 481082 10316 481088 10328
rect 382148 10288 481088 10316
rect 382148 10276 382154 10288
rect 481082 10276 481088 10288
rect 481140 10276 481146 10328
rect 125962 9704 125968 9716
rect 125923 9676 125968 9704
rect 125962 9664 125968 9676
rect 126020 9664 126026 9716
rect 133138 9664 133144 9716
rect 133196 9704 133202 9716
rect 133322 9704 133328 9716
rect 133196 9676 133328 9704
rect 133196 9664 133202 9676
rect 133322 9664 133328 9676
rect 133380 9664 133386 9716
rect 140869 9707 140927 9713
rect 140869 9673 140881 9707
rect 140915 9704 140927 9707
rect 141050 9704 141056 9716
rect 140915 9676 141056 9704
rect 140915 9673 140927 9676
rect 140869 9667 140927 9673
rect 141050 9664 141056 9676
rect 141108 9664 141114 9716
rect 168374 9704 168380 9716
rect 168335 9676 168380 9704
rect 168374 9664 168380 9676
rect 168432 9664 168438 9716
rect 179693 9707 179751 9713
rect 179693 9673 179705 9707
rect 179739 9704 179751 9707
rect 179782 9704 179788 9716
rect 179739 9676 179788 9704
rect 179739 9673 179751 9676
rect 179693 9667 179751 9673
rect 179782 9664 179788 9676
rect 179840 9664 179846 9716
rect 207198 9704 207204 9716
rect 207159 9676 207204 9704
rect 207198 9664 207204 9676
rect 207256 9664 207262 9716
rect 214101 9707 214159 9713
rect 214101 9673 214113 9707
rect 214147 9704 214159 9707
rect 214190 9704 214196 9716
rect 214147 9676 214196 9704
rect 214147 9673 214159 9676
rect 214101 9667 214159 9673
rect 214190 9664 214196 9676
rect 214248 9664 214254 9716
rect 215389 9707 215447 9713
rect 215389 9673 215401 9707
rect 215435 9704 215447 9707
rect 215478 9704 215484 9716
rect 215435 9676 215484 9704
rect 215435 9673 215447 9676
rect 215389 9667 215447 9673
rect 215478 9664 215484 9676
rect 215536 9664 215542 9716
rect 238386 9704 238392 9716
rect 238347 9676 238392 9704
rect 238386 9664 238392 9676
rect 238444 9664 238450 9716
rect 274821 9707 274879 9713
rect 274821 9673 274833 9707
rect 274867 9704 274879 9707
rect 275278 9704 275284 9716
rect 274867 9676 275284 9704
rect 274867 9673 274879 9676
rect 274821 9667 274879 9673
rect 275278 9664 275284 9676
rect 275336 9664 275342 9716
rect 280430 9664 280436 9716
rect 280488 9704 280494 9716
rect 281258 9704 281264 9716
rect 280488 9676 281264 9704
rect 280488 9664 280494 9676
rect 281258 9664 281264 9676
rect 281316 9664 281322 9716
rect 282914 9664 282920 9716
rect 282972 9704 282978 9716
rect 283374 9704 283380 9716
rect 282972 9676 283380 9704
rect 282972 9664 282978 9676
rect 283374 9664 283380 9676
rect 283432 9664 283438 9716
rect 290918 9704 290924 9716
rect 290879 9676 290924 9704
rect 290918 9664 290924 9676
rect 290976 9664 290982 9716
rect 325697 9707 325755 9713
rect 325697 9673 325709 9707
rect 325743 9704 325755 9707
rect 326246 9704 326252 9716
rect 325743 9676 326252 9704
rect 325743 9673 325755 9676
rect 325697 9667 325755 9673
rect 326246 9664 326252 9676
rect 326304 9664 326310 9716
rect 383286 9704 383292 9716
rect 383247 9676 383292 9704
rect 383286 9664 383292 9676
rect 383344 9664 383350 9716
rect 57606 9596 57612 9648
rect 57664 9636 57670 9648
rect 162854 9636 162860 9648
rect 57664 9608 162860 9636
rect 57664 9596 57670 9608
rect 162854 9596 162860 9608
rect 162912 9596 162918 9648
rect 368382 9596 368388 9648
rect 368440 9636 368446 9648
rect 454862 9636 454868 9648
rect 368440 9608 454868 9636
rect 368440 9596 368446 9608
rect 454862 9596 454868 9608
rect 454920 9596 454926 9648
rect 58802 9528 58808 9580
rect 58860 9568 58866 9580
rect 164326 9568 164332 9580
rect 58860 9540 164332 9568
rect 58860 9528 58866 9540
rect 164326 9528 164332 9540
rect 164384 9528 164390 9580
rect 371142 9528 371148 9580
rect 371200 9568 371206 9580
rect 458450 9568 458456 9580
rect 371200 9540 458456 9568
rect 371200 9528 371206 9540
rect 458450 9528 458456 9540
rect 458508 9528 458514 9580
rect 55214 9460 55220 9512
rect 55272 9500 55278 9512
rect 161750 9500 161756 9512
rect 55272 9472 161756 9500
rect 55272 9460 55278 9472
rect 161750 9460 161756 9472
rect 161808 9460 161814 9512
rect 372430 9460 372436 9512
rect 372488 9500 372494 9512
rect 462038 9500 462044 9512
rect 372488 9472 462044 9500
rect 372488 9460 372494 9472
rect 462038 9460 462044 9472
rect 462096 9460 462102 9512
rect 51626 9392 51632 9444
rect 51684 9432 51690 9444
rect 160186 9432 160192 9444
rect 51684 9404 160192 9432
rect 51684 9392 51690 9404
rect 160186 9392 160192 9404
rect 160244 9392 160250 9444
rect 419442 9392 419448 9444
rect 419500 9432 419506 9444
rect 552382 9432 552388 9444
rect 419500 9404 552388 9432
rect 419500 9392 419506 9404
rect 552382 9392 552388 9404
rect 552440 9392 552446 9444
rect 43346 9324 43352 9376
rect 43404 9364 43410 9376
rect 156046 9364 156052 9376
rect 43404 9336 156052 9364
rect 43404 9324 43410 9336
rect 156046 9324 156052 9336
rect 156104 9324 156110 9376
rect 420454 9324 420460 9376
rect 420512 9364 420518 9376
rect 555970 9364 555976 9376
rect 420512 9336 555976 9364
rect 420512 9324 420518 9336
rect 555970 9324 555976 9336
rect 556028 9324 556034 9376
rect 40954 9256 40960 9308
rect 41012 9296 41018 9308
rect 154666 9296 154672 9308
rect 41012 9268 154672 9296
rect 41012 9256 41018 9268
rect 154666 9256 154672 9268
rect 154724 9256 154730 9308
rect 422110 9256 422116 9308
rect 422168 9296 422174 9308
rect 559558 9296 559564 9308
rect 422168 9268 559564 9296
rect 422168 9256 422174 9268
rect 559558 9256 559564 9268
rect 559616 9256 559622 9308
rect 36170 9188 36176 9240
rect 36228 9228 36234 9240
rect 151814 9228 151820 9240
rect 36228 9200 151820 9228
rect 36228 9188 36234 9200
rect 151814 9188 151820 9200
rect 151872 9188 151878 9240
rect 409506 9188 409512 9240
rect 409564 9228 409570 9240
rect 409782 9228 409788 9240
rect 409564 9200 409788 9228
rect 409564 9188 409570 9200
rect 409782 9188 409788 9200
rect 409840 9188 409846 9240
rect 424962 9188 424968 9240
rect 425020 9228 425026 9240
rect 563146 9228 563152 9240
rect 425020 9200 563152 9228
rect 425020 9188 425026 9200
rect 563146 9188 563152 9200
rect 563204 9188 563210 9240
rect 18322 9120 18328 9172
rect 18380 9160 18386 9172
rect 135438 9160 135444 9172
rect 18380 9132 135444 9160
rect 18380 9120 18386 9132
rect 135438 9120 135444 9132
rect 135496 9120 135502 9172
rect 350350 9120 350356 9172
rect 350408 9160 350414 9172
rect 420362 9160 420368 9172
rect 350408 9132 420368 9160
rect 350408 9120 350414 9132
rect 420362 9120 420368 9132
rect 420420 9120 420426 9172
rect 425974 9120 425980 9172
rect 426032 9160 426038 9172
rect 566734 9160 566740 9172
rect 426032 9132 566740 9160
rect 426032 9120 426038 9132
rect 566734 9120 566740 9132
rect 566792 9120 566798 9172
rect 20714 9052 20720 9104
rect 20772 9092 20778 9104
rect 143626 9092 143632 9104
rect 20772 9064 143632 9092
rect 20772 9052 20778 9064
rect 143626 9052 143632 9064
rect 143684 9052 143690 9104
rect 353202 9052 353208 9104
rect 353260 9092 353266 9104
rect 423950 9092 423956 9104
rect 353260 9064 423956 9092
rect 353260 9052 353266 9064
rect 423950 9052 423956 9064
rect 424008 9052 424014 9104
rect 427630 9052 427636 9104
rect 427688 9092 427694 9104
rect 570230 9092 570236 9104
rect 427688 9064 570236 9092
rect 427688 9052 427694 9064
rect 570230 9052 570236 9064
rect 570288 9052 570294 9104
rect 11238 8984 11244 9036
rect 11296 9024 11302 9036
rect 139486 9024 139492 9036
rect 11296 8996 139492 9024
rect 11296 8984 11302 8996
rect 139486 8984 139492 8996
rect 139544 8984 139550 9036
rect 354490 8984 354496 9036
rect 354548 9024 354554 9036
rect 427538 9024 427544 9036
rect 354548 8996 427544 9024
rect 354548 8984 354554 8996
rect 427538 8984 427544 8996
rect 427596 8984 427602 9036
rect 431494 8984 431500 9036
rect 431552 9024 431558 9036
rect 577406 9024 577412 9036
rect 431552 8996 577412 9024
rect 431552 8984 431558 8996
rect 577406 8984 577412 8996
rect 577464 8984 577470 9036
rect 5258 8916 5264 8968
rect 5316 8956 5322 8968
rect 136818 8956 136824 8968
rect 5316 8928 136824 8956
rect 5316 8916 5322 8928
rect 136818 8916 136824 8928
rect 136876 8916 136882 8968
rect 143258 8916 143264 8968
rect 143316 8956 143322 8968
rect 207198 8956 207204 8968
rect 143316 8928 207204 8956
rect 143316 8916 143322 8928
rect 207198 8916 207204 8928
rect 207256 8916 207262 8968
rect 355870 8916 355876 8968
rect 355928 8956 355934 8968
rect 431126 8956 431132 8968
rect 355928 8928 431132 8956
rect 355928 8916 355934 8928
rect 431126 8916 431132 8928
rect 431184 8916 431190 8968
rect 433150 8916 433156 8968
rect 433208 8956 433214 8968
rect 580994 8956 581000 8968
rect 433208 8928 581000 8956
rect 433208 8916 433214 8928
rect 580994 8916 581000 8928
rect 581052 8916 581058 8968
rect 64782 8848 64788 8900
rect 64840 8888 64846 8900
rect 167086 8888 167092 8900
rect 64840 8860 167092 8888
rect 64840 8848 64846 8860
rect 167086 8848 167092 8860
rect 167144 8848 167150 8900
rect 369762 8848 369768 8900
rect 369820 8888 369826 8900
rect 456058 8888 456064 8900
rect 369820 8860 456064 8888
rect 369820 8848 369826 8860
rect 456058 8848 456064 8860
rect 456116 8848 456122 8900
rect 71866 8780 71872 8832
rect 71924 8820 71930 8832
rect 169846 8820 169852 8832
rect 71924 8792 169852 8820
rect 71924 8780 71930 8792
rect 169846 8780 169852 8792
rect 169904 8780 169910 8832
rect 366910 8780 366916 8832
rect 366968 8820 366974 8832
rect 452470 8820 452476 8832
rect 366968 8792 452476 8820
rect 366968 8780 366974 8792
rect 452470 8780 452476 8792
rect 452528 8780 452534 8832
rect 79042 8712 79048 8764
rect 79100 8752 79106 8764
rect 173986 8752 173992 8764
rect 79100 8724 173992 8752
rect 79100 8712 79106 8724
rect 173986 8712 173992 8724
rect 174044 8712 174050 8764
rect 365530 8712 365536 8764
rect 365588 8752 365594 8764
rect 448974 8752 448980 8764
rect 365588 8724 448980 8752
rect 365588 8712 365594 8724
rect 448974 8712 448980 8724
rect 449032 8712 449038 8764
rect 120626 8644 120632 8696
rect 120684 8684 120690 8696
rect 175458 8684 175464 8696
rect 120684 8656 175464 8684
rect 120684 8644 120690 8656
rect 175458 8644 175464 8656
rect 175516 8644 175522 8696
rect 361390 8644 361396 8696
rect 361448 8684 361454 8696
rect 441798 8684 441804 8696
rect 361448 8656 441804 8684
rect 361448 8644 361454 8656
rect 441798 8644 441804 8656
rect 441856 8644 441862 8696
rect 106366 8576 106372 8628
rect 106424 8616 106430 8628
rect 133138 8616 133144 8628
rect 106424 8588 133144 8616
rect 106424 8576 106430 8588
rect 133138 8576 133144 8588
rect 133196 8576 133202 8628
rect 364242 8576 364248 8628
rect 364300 8616 364306 8628
rect 445386 8616 445392 8628
rect 364300 8588 445392 8616
rect 364300 8576 364306 8588
rect 445386 8576 445392 8588
rect 445444 8576 445450 8628
rect 360010 8508 360016 8560
rect 360068 8548 360074 8560
rect 438210 8548 438216 8560
rect 360068 8520 438216 8548
rect 360068 8508 360074 8520
rect 438210 8508 438216 8520
rect 438268 8508 438274 8560
rect 358630 8440 358636 8492
rect 358688 8480 358694 8492
rect 434622 8480 434628 8492
rect 358688 8452 434628 8480
rect 358688 8440 358694 8452
rect 434622 8440 434628 8452
rect 434680 8440 434686 8492
rect 125597 8347 125655 8353
rect 125597 8313 125609 8347
rect 125643 8344 125655 8347
rect 129274 8344 129280 8356
rect 125643 8316 129280 8344
rect 125643 8313 125655 8316
rect 125597 8307 125655 8313
rect 129274 8304 129280 8316
rect 129332 8304 129338 8356
rect 301869 8347 301927 8353
rect 301869 8313 301881 8347
rect 301915 8344 301927 8347
rect 302050 8344 302056 8356
rect 301915 8316 302056 8344
rect 301915 8313 301927 8316
rect 301869 8307 301927 8313
rect 302050 8304 302056 8316
rect 302108 8304 302114 8356
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 131758 8276 131764 8288
rect 3476 8248 131764 8276
rect 3476 8236 3482 8248
rect 131758 8236 131764 8248
rect 131816 8236 131822 8288
rect 133782 8236 133788 8288
rect 133840 8276 133846 8288
rect 203058 8276 203064 8288
rect 133840 8248 203064 8276
rect 133840 8236 133846 8248
rect 203058 8236 203064 8248
rect 203116 8236 203122 8288
rect 384942 8236 384948 8288
rect 385000 8276 385006 8288
rect 414753 8279 414811 8285
rect 414753 8276 414765 8279
rect 385000 8248 414765 8276
rect 385000 8236 385006 8248
rect 414753 8245 414765 8248
rect 414799 8245 414811 8279
rect 414753 8239 414811 8245
rect 415029 8279 415087 8285
rect 415029 8245 415041 8279
rect 415075 8276 415087 8279
rect 486970 8276 486976 8288
rect 415075 8248 486976 8276
rect 415075 8245 415087 8248
rect 415029 8239 415087 8245
rect 486970 8236 486976 8248
rect 487028 8236 487034 8288
rect 114738 8168 114744 8220
rect 114796 8208 114802 8220
rect 191926 8208 191932 8220
rect 114796 8180 191932 8208
rect 114796 8168 114802 8180
rect 191926 8168 191932 8180
rect 191984 8168 191990 8220
rect 387610 8168 387616 8220
rect 387668 8208 387674 8220
rect 490558 8208 490564 8220
rect 387668 8180 490564 8208
rect 387668 8168 387674 8180
rect 490558 8168 490564 8180
rect 490616 8168 490622 8220
rect 107562 8100 107568 8152
rect 107620 8140 107626 8152
rect 189166 8140 189172 8152
rect 107620 8112 189172 8140
rect 107620 8100 107626 8112
rect 189166 8100 189172 8112
rect 189224 8100 189230 8152
rect 388898 8100 388904 8152
rect 388956 8140 388962 8152
rect 494146 8140 494152 8152
rect 388956 8112 494152 8140
rect 388956 8100 388962 8112
rect 494146 8100 494152 8112
rect 494204 8100 494210 8152
rect 100478 8032 100484 8084
rect 100536 8072 100542 8084
rect 184934 8072 184940 8084
rect 100536 8044 184940 8072
rect 100536 8032 100542 8044
rect 184934 8032 184940 8044
rect 184992 8032 184998 8084
rect 390462 8032 390468 8084
rect 390520 8072 390526 8084
rect 497734 8072 497740 8084
rect 390520 8044 497740 8072
rect 390520 8032 390526 8044
rect 497734 8032 497740 8044
rect 497792 8032 497798 8084
rect 48130 7964 48136 8016
rect 48188 8004 48194 8016
rect 158806 8004 158812 8016
rect 48188 7976 158812 8004
rect 48188 7964 48194 7976
rect 158806 7964 158812 7976
rect 158864 7964 158870 8016
rect 393130 7964 393136 8016
rect 393188 8004 393194 8016
rect 501230 8004 501236 8016
rect 393188 7976 501236 8004
rect 393188 7964 393194 7976
rect 501230 7964 501236 7976
rect 501288 7964 501294 8016
rect 13630 7896 13636 7948
rect 13688 7936 13694 7948
rect 141050 7936 141056 7948
rect 13688 7908 141056 7936
rect 13688 7896 13694 7908
rect 141050 7896 141056 7908
rect 141108 7896 141114 7948
rect 394326 7896 394332 7948
rect 394384 7936 394390 7948
rect 504818 7936 504824 7948
rect 394384 7908 504824 7936
rect 394384 7896 394390 7908
rect 504818 7896 504824 7908
rect 504876 7896 504882 7948
rect 7650 7828 7656 7880
rect 7708 7868 7714 7880
rect 136726 7868 136732 7880
rect 7708 7840 136732 7868
rect 7708 7828 7714 7840
rect 136726 7828 136732 7840
rect 136784 7828 136790 7880
rect 140866 7828 140872 7880
rect 140924 7868 140930 7880
rect 205634 7868 205640 7880
rect 140924 7840 205640 7868
rect 140924 7828 140930 7840
rect 205634 7828 205640 7840
rect 205692 7828 205698 7880
rect 395890 7828 395896 7880
rect 395948 7868 395954 7880
rect 508406 7868 508412 7880
rect 395948 7840 508412 7868
rect 395948 7828 395954 7840
rect 508406 7828 508412 7840
rect 508464 7828 508470 7880
rect 4062 7760 4068 7812
rect 4120 7800 4126 7812
rect 135254 7800 135260 7812
rect 4120 7772 135260 7800
rect 4120 7760 4126 7772
rect 135254 7760 135260 7772
rect 135312 7760 135318 7812
rect 139670 7760 139676 7812
rect 139728 7800 139734 7812
rect 205726 7800 205732 7812
rect 139728 7772 205732 7800
rect 139728 7760 139734 7772
rect 205726 7760 205732 7772
rect 205784 7760 205790 7812
rect 413922 7760 413928 7812
rect 413980 7800 413986 7812
rect 541710 7800 541716 7812
rect 413980 7772 541716 7800
rect 413980 7760 413986 7772
rect 541710 7760 541716 7772
rect 541768 7760 541774 7812
rect 1670 7692 1676 7744
rect 1728 7732 1734 7744
rect 134058 7732 134064 7744
rect 1728 7704 134064 7732
rect 1728 7692 1734 7704
rect 134058 7692 134064 7704
rect 134116 7692 134122 7744
rect 136082 7692 136088 7744
rect 136140 7732 136146 7744
rect 202966 7732 202972 7744
rect 136140 7704 202972 7732
rect 136140 7692 136146 7704
rect 202966 7692 202972 7704
rect 203024 7692 203030 7744
rect 344738 7692 344744 7744
rect 344796 7732 344802 7744
rect 409690 7732 409696 7744
rect 344796 7704 409696 7732
rect 344796 7692 344802 7704
rect 409690 7692 409696 7704
rect 409748 7692 409754 7744
rect 414934 7692 414940 7744
rect 414992 7732 414998 7744
rect 545298 7732 545304 7744
rect 414992 7704 545304 7732
rect 414992 7692 414998 7704
rect 545298 7692 545304 7704
rect 545356 7692 545362 7744
rect 2866 7624 2872 7676
rect 2924 7664 2930 7676
rect 135346 7664 135352 7676
rect 2924 7636 135352 7664
rect 2924 7624 2930 7636
rect 135346 7624 135352 7636
rect 135404 7624 135410 7676
rect 137278 7624 137284 7676
rect 137336 7664 137342 7676
rect 204346 7664 204352 7676
rect 137336 7636 204352 7664
rect 137336 7624 137342 7636
rect 204346 7624 204352 7636
rect 204404 7624 204410 7676
rect 347682 7624 347688 7676
rect 347740 7664 347746 7676
rect 413278 7664 413284 7676
rect 347740 7636 413284 7664
rect 347740 7624 347746 7636
rect 413278 7624 413284 7636
rect 413336 7624 413342 7676
rect 416590 7624 416596 7676
rect 416648 7664 416654 7676
rect 548886 7664 548892 7676
rect 416648 7636 548892 7664
rect 416648 7624 416654 7636
rect 548886 7624 548892 7636
rect 548944 7624 548950 7676
rect 566 7556 572 7608
rect 624 7596 630 7608
rect 133874 7596 133880 7608
rect 624 7568 133880 7596
rect 624 7556 630 7568
rect 133874 7556 133880 7568
rect 133932 7556 133938 7608
rect 134886 7556 134892 7608
rect 134944 7596 134950 7608
rect 202874 7596 202880 7608
rect 134944 7568 202880 7596
rect 134944 7556 134950 7568
rect 202874 7556 202880 7568
rect 202932 7556 202938 7608
rect 348970 7556 348976 7608
rect 349028 7596 349034 7608
rect 412637 7599 412695 7605
rect 412637 7596 412649 7599
rect 349028 7568 412649 7596
rect 349028 7556 349034 7568
rect 412637 7565 412649 7568
rect 412683 7565 412695 7599
rect 412637 7559 412695 7565
rect 416774 7556 416780 7608
rect 416832 7596 416838 7608
rect 417970 7596 417976 7608
rect 416832 7568 417976 7596
rect 416832 7556 416838 7568
rect 417970 7556 417976 7568
rect 418028 7556 418034 7608
rect 430482 7556 430488 7608
rect 430540 7596 430546 7608
rect 573818 7596 573824 7608
rect 430540 7568 573824 7596
rect 430540 7556 430546 7568
rect 573818 7556 573824 7568
rect 573876 7556 573882 7608
rect 121822 7488 121828 7540
rect 121880 7528 121886 7540
rect 196066 7528 196072 7540
rect 121880 7500 196072 7528
rect 121880 7488 121886 7500
rect 196066 7488 196072 7500
rect 196124 7488 196130 7540
rect 383286 7488 383292 7540
rect 383344 7528 383350 7540
rect 383344 7500 477448 7528
rect 383344 7488 383350 7500
rect 126606 7420 126612 7472
rect 126664 7460 126670 7472
rect 198826 7460 198832 7472
rect 126664 7432 198832 7460
rect 126664 7420 126670 7432
rect 198826 7420 198832 7432
rect 198884 7420 198890 7472
rect 367002 7420 367008 7472
rect 367060 7460 367066 7472
rect 451274 7460 451280 7472
rect 367060 7432 451280 7460
rect 367060 7420 367066 7432
rect 451274 7420 451280 7432
rect 451332 7420 451338 7472
rect 123113 7395 123171 7401
rect 123113 7361 123125 7395
rect 123159 7392 123171 7395
rect 127618 7392 127624 7404
rect 123159 7364 127624 7392
rect 123159 7361 123171 7364
rect 123113 7355 123171 7361
rect 127618 7352 127624 7364
rect 127676 7352 127682 7404
rect 197446 7392 197452 7404
rect 127728 7364 197452 7392
rect 77846 7284 77852 7336
rect 77904 7324 77910 7336
rect 77904 7296 123616 7324
rect 77904 7284 77910 7296
rect 117130 7216 117136 7268
rect 117188 7256 117194 7268
rect 123113 7259 123171 7265
rect 123113 7256 123125 7259
rect 117188 7228 123125 7256
rect 117188 7216 117194 7228
rect 123113 7225 123125 7228
rect 123159 7225 123171 7259
rect 123113 7219 123171 7225
rect 84930 7148 84936 7200
rect 84988 7188 84994 7200
rect 123588 7188 123616 7296
rect 125410 7284 125416 7336
rect 125468 7324 125474 7336
rect 127728 7324 127756 7364
rect 197446 7352 197452 7364
rect 197504 7352 197510 7404
rect 365622 7352 365628 7404
rect 365680 7392 365686 7404
rect 447778 7392 447784 7404
rect 365680 7364 447784 7392
rect 365680 7352 365686 7364
rect 447778 7352 447784 7364
rect 447836 7352 447842 7404
rect 477420 7392 477448 7500
rect 477494 7488 477500 7540
rect 477552 7528 477558 7540
rect 478690 7528 478696 7540
rect 477552 7500 478696 7528
rect 477552 7488 477558 7500
rect 478690 7488 478696 7500
rect 478748 7488 478754 7540
rect 483474 7392 483480 7404
rect 477420 7364 483480 7392
rect 483474 7352 483480 7364
rect 483532 7352 483538 7404
rect 125468 7296 127756 7324
rect 125468 7284 125474 7296
rect 128998 7284 129004 7336
rect 129056 7324 129062 7336
rect 200206 7324 200212 7336
rect 129056 7296 200212 7324
rect 129056 7284 129062 7296
rect 200206 7284 200212 7296
rect 200264 7284 200270 7336
rect 362862 7284 362868 7336
rect 362920 7324 362926 7336
rect 444190 7324 444196 7336
rect 362920 7296 444196 7324
rect 362920 7284 362926 7296
rect 444190 7284 444196 7296
rect 444248 7284 444254 7336
rect 127802 7216 127808 7268
rect 127860 7256 127866 7268
rect 198734 7256 198740 7268
rect 127860 7228 198740 7256
rect 127860 7216 127866 7228
rect 198734 7216 198740 7228
rect 198792 7216 198798 7268
rect 361482 7216 361488 7268
rect 361540 7256 361546 7268
rect 440602 7256 440608 7268
rect 361540 7228 440608 7256
rect 361540 7216 361546 7228
rect 440602 7216 440608 7228
rect 440660 7216 440666 7268
rect 129090 7188 129096 7200
rect 84988 7160 123524 7188
rect 123588 7160 129096 7188
rect 84988 7148 84994 7160
rect 95694 7080 95700 7132
rect 95752 7120 95758 7132
rect 123496 7120 123524 7160
rect 129090 7148 129096 7160
rect 129148 7148 129154 7200
rect 131390 7148 131396 7200
rect 131448 7188 131454 7200
rect 201586 7188 201592 7200
rect 131448 7160 201592 7188
rect 131448 7148 131454 7160
rect 201586 7148 201592 7160
rect 201644 7148 201650 7200
rect 360102 7148 360108 7200
rect 360160 7188 360166 7200
rect 437014 7188 437020 7200
rect 360160 7160 437020 7188
rect 360160 7148 360166 7160
rect 437014 7148 437020 7160
rect 437072 7148 437078 7200
rect 129182 7120 129188 7132
rect 95752 7092 120764 7120
rect 123496 7092 129188 7120
rect 95752 7080 95758 7092
rect 120736 6984 120764 7092
rect 129182 7080 129188 7092
rect 129240 7080 129246 7132
rect 130194 7080 130200 7132
rect 130252 7120 130258 7132
rect 200114 7120 200120 7132
rect 130252 7092 200120 7120
rect 130252 7080 130258 7092
rect 200114 7080 200120 7092
rect 200172 7080 200178 7132
rect 358722 7080 358728 7132
rect 358780 7120 358786 7132
rect 435818 7120 435824 7132
rect 358780 7092 435824 7120
rect 358780 7080 358786 7092
rect 435818 7080 435824 7092
rect 435876 7080 435882 7132
rect 132586 7012 132592 7064
rect 132644 7052 132650 7064
rect 201494 7052 201500 7064
rect 132644 7024 201500 7052
rect 132644 7012 132650 7024
rect 201494 7012 201500 7024
rect 201552 7012 201558 7064
rect 412637 7055 412695 7061
rect 412637 7021 412649 7055
rect 412683 7052 412695 7055
rect 416866 7052 416872 7064
rect 412683 7024 416872 7052
rect 412683 7021 412695 7024
rect 412637 7015 412695 7021
rect 416866 7012 416872 7024
rect 416924 7012 416930 7064
rect 125597 6987 125655 6993
rect 125597 6984 125609 6987
rect 120736 6956 125609 6984
rect 125597 6953 125609 6956
rect 125643 6953 125655 6987
rect 125597 6947 125655 6953
rect 227806 6916 227812 6928
rect 227767 6888 227812 6916
rect 227806 6876 227812 6888
rect 227864 6876 227870 6928
rect 230106 6916 230112 6928
rect 230067 6888 230112 6916
rect 230106 6876 230112 6888
rect 230164 6876 230170 6928
rect 94498 6808 94504 6860
rect 94556 6848 94562 6860
rect 182266 6848 182272 6860
rect 94556 6820 182272 6848
rect 94556 6808 94562 6820
rect 182266 6808 182272 6820
rect 182324 6808 182330 6860
rect 317230 6808 317236 6860
rect 317288 6848 317294 6860
rect 356146 6848 356152 6860
rect 317288 6820 356152 6848
rect 317288 6808 317294 6820
rect 356146 6808 356152 6820
rect 356204 6808 356210 6860
rect 391750 6808 391756 6860
rect 391808 6848 391814 6860
rect 498930 6848 498936 6860
rect 391808 6820 498936 6848
rect 391808 6808 391814 6820
rect 498930 6808 498936 6820
rect 498988 6808 498994 6860
rect 93302 6740 93308 6792
rect 93360 6780 93366 6792
rect 180978 6780 180984 6792
rect 93360 6752 180984 6780
rect 93360 6740 93366 6752
rect 180978 6740 180984 6752
rect 181036 6740 181042 6792
rect 326890 6740 326896 6792
rect 326948 6780 326954 6792
rect 373994 6780 374000 6792
rect 326948 6752 374000 6780
rect 326948 6740 326954 6752
rect 373994 6740 374000 6752
rect 374052 6740 374058 6792
rect 393222 6740 393228 6792
rect 393280 6780 393286 6792
rect 502426 6780 502432 6792
rect 393280 6752 502432 6780
rect 393280 6740 393286 6752
rect 502426 6740 502432 6752
rect 502484 6740 502490 6792
rect 90910 6672 90916 6724
rect 90968 6712 90974 6724
rect 180886 6712 180892 6724
rect 90968 6684 180892 6712
rect 90968 6672 90974 6684
rect 180886 6672 180892 6684
rect 180944 6672 180950 6724
rect 328178 6672 328184 6724
rect 328236 6712 328242 6724
rect 377582 6712 377588 6724
rect 328236 6684 377588 6712
rect 328236 6672 328242 6684
rect 377582 6672 377588 6684
rect 377640 6672 377646 6724
rect 394602 6672 394608 6724
rect 394660 6712 394666 6724
rect 506014 6712 506020 6724
rect 394660 6684 506020 6712
rect 394660 6672 394666 6684
rect 506014 6672 506020 6684
rect 506072 6672 506078 6724
rect 86126 6604 86132 6656
rect 86184 6644 86190 6656
rect 178126 6644 178132 6656
rect 86184 6616 178132 6644
rect 86184 6604 86190 6616
rect 178126 6604 178132 6616
rect 178184 6604 178190 6656
rect 331030 6604 331036 6656
rect 331088 6644 331094 6656
rect 381170 6644 381176 6656
rect 331088 6616 381176 6644
rect 331088 6604 331094 6616
rect 381170 6604 381176 6616
rect 381228 6604 381234 6656
rect 397362 6604 397368 6656
rect 397420 6644 397426 6656
rect 509602 6644 509608 6656
rect 397420 6616 509608 6644
rect 397420 6604 397426 6616
rect 509602 6604 509608 6616
rect 509660 6604 509666 6656
rect 82630 6536 82636 6588
rect 82688 6576 82694 6588
rect 175366 6576 175372 6588
rect 82688 6548 175372 6576
rect 82688 6536 82694 6548
rect 175366 6536 175372 6548
rect 175424 6536 175430 6588
rect 332410 6536 332416 6588
rect 332468 6576 332474 6588
rect 384666 6576 384672 6588
rect 332468 6548 384672 6576
rect 332468 6536 332474 6548
rect 384666 6536 384672 6548
rect 384724 6536 384730 6588
rect 398650 6536 398656 6588
rect 398708 6576 398714 6588
rect 513190 6576 513196 6588
rect 398708 6548 513196 6576
rect 398708 6536 398714 6548
rect 513190 6536 513196 6548
rect 513248 6536 513254 6588
rect 8846 6468 8852 6520
rect 8904 6508 8910 6520
rect 103514 6508 103520 6520
rect 8904 6480 103520 6508
rect 8904 6468 8910 6480
rect 103514 6468 103520 6480
rect 103572 6468 103578 6520
rect 105170 6468 105176 6520
rect 105228 6508 105234 6520
rect 187694 6508 187700 6520
rect 105228 6480 187700 6508
rect 105228 6468 105234 6480
rect 187694 6468 187700 6480
rect 187752 6468 187758 6520
rect 336642 6468 336648 6520
rect 336700 6508 336706 6520
rect 391842 6508 391848 6520
rect 336700 6480 391848 6508
rect 336700 6468 336706 6480
rect 391842 6468 391848 6480
rect 391900 6468 391906 6520
rect 399938 6468 399944 6520
rect 399996 6508 400002 6520
rect 516778 6508 516784 6520
rect 399996 6480 516784 6508
rect 399996 6468 400002 6480
rect 516778 6468 516784 6480
rect 516836 6468 516842 6520
rect 75454 6400 75460 6452
rect 75512 6440 75518 6452
rect 172606 6440 172612 6452
rect 75512 6412 172612 6440
rect 75512 6400 75518 6412
rect 172606 6400 172612 6412
rect 172664 6400 172670 6452
rect 333698 6400 333704 6452
rect 333756 6440 333762 6452
rect 388254 6440 388260 6452
rect 333756 6412 388260 6440
rect 333756 6400 333762 6412
rect 388254 6400 388260 6412
rect 388312 6400 388318 6452
rect 402790 6400 402796 6452
rect 402848 6440 402854 6452
rect 520274 6440 520280 6452
rect 402848 6412 520280 6440
rect 402848 6400 402854 6412
rect 520274 6400 520280 6412
rect 520332 6400 520338 6452
rect 68278 6332 68284 6384
rect 68336 6372 68342 6384
rect 168374 6372 168380 6384
rect 68336 6344 168380 6372
rect 68336 6332 68342 6344
rect 168374 6332 168380 6344
rect 168432 6332 168438 6384
rect 337930 6332 337936 6384
rect 337988 6372 337994 6384
rect 395430 6372 395436 6384
rect 337988 6344 395436 6372
rect 337988 6332 337994 6344
rect 395430 6332 395436 6344
rect 395488 6332 395494 6384
rect 404170 6332 404176 6384
rect 404228 6372 404234 6384
rect 523862 6372 523868 6384
rect 404228 6344 523868 6372
rect 404228 6332 404234 6344
rect 523862 6332 523868 6344
rect 523920 6332 523926 6384
rect 61194 6264 61200 6316
rect 61252 6304 61258 6316
rect 164418 6304 164424 6316
rect 61252 6276 164424 6304
rect 61252 6264 61258 6276
rect 164418 6264 164424 6276
rect 164476 6264 164482 6316
rect 342162 6264 342168 6316
rect 342220 6304 342226 6316
rect 402514 6304 402520 6316
rect 342220 6276 402520 6304
rect 342220 6264 342226 6276
rect 402514 6264 402520 6276
rect 402572 6264 402578 6316
rect 408402 6264 408408 6316
rect 408460 6304 408466 6316
rect 531038 6304 531044 6316
rect 408460 6276 531044 6304
rect 408460 6264 408466 6276
rect 531038 6264 531044 6276
rect 531096 6264 531102 6316
rect 54018 6196 54024 6248
rect 54076 6236 54082 6248
rect 161474 6236 161480 6248
rect 54076 6208 161480 6236
rect 54076 6196 54082 6208
rect 161474 6196 161480 6208
rect 161532 6196 161538 6248
rect 339310 6196 339316 6248
rect 339368 6236 339374 6248
rect 399018 6236 399024 6248
rect 339368 6208 399024 6236
rect 339368 6196 339374 6208
rect 399018 6196 399024 6208
rect 399076 6196 399082 6248
rect 405550 6196 405556 6248
rect 405608 6236 405614 6248
rect 527450 6236 527456 6248
rect 405608 6208 527456 6236
rect 405608 6196 405614 6208
rect 527450 6196 527456 6208
rect 527508 6196 527514 6248
rect 44542 6128 44548 6180
rect 44600 6168 44606 6180
rect 155954 6168 155960 6180
rect 44600 6140 155960 6168
rect 44600 6128 44606 6140
rect 155954 6128 155960 6140
rect 156012 6128 156018 6180
rect 157518 6128 157524 6180
rect 157576 6168 157582 6180
rect 214190 6168 214196 6180
rect 157576 6140 214196 6168
rect 157576 6128 157582 6140
rect 214190 6128 214196 6140
rect 214248 6128 214254 6180
rect 343450 6128 343456 6180
rect 343508 6168 343514 6180
rect 406102 6168 406108 6180
rect 343508 6140 406108 6168
rect 343508 6128 343514 6140
rect 406102 6128 406108 6140
rect 406160 6128 406166 6180
rect 409598 6128 409604 6180
rect 409656 6168 409662 6180
rect 534534 6168 534540 6180
rect 409656 6140 534540 6168
rect 409656 6128 409662 6140
rect 534534 6128 534540 6140
rect 534592 6128 534598 6180
rect 101582 6060 101588 6112
rect 101640 6100 101646 6112
rect 186498 6100 186504 6112
rect 101640 6072 186504 6100
rect 101640 6060 101646 6072
rect 186498 6060 186504 6072
rect 186556 6060 186562 6112
rect 318702 6060 318708 6112
rect 318760 6100 318766 6112
rect 358538 6100 358544 6112
rect 318760 6072 358544 6100
rect 318760 6060 318766 6072
rect 358538 6060 358544 6072
rect 358596 6060 358602 6112
rect 388990 6060 388996 6112
rect 389048 6100 389054 6112
rect 495342 6100 495348 6112
rect 389048 6072 495348 6100
rect 389048 6060 389054 6072
rect 495342 6060 495348 6072
rect 495400 6060 495406 6112
rect 98086 5992 98092 6044
rect 98144 6032 98150 6044
rect 183830 6032 183836 6044
rect 98144 6004 183836 6032
rect 98144 5992 98150 6004
rect 183830 5992 183836 6004
rect 183888 5992 183894 6044
rect 317138 5992 317144 6044
rect 317196 6032 317202 6044
rect 354950 6032 354956 6044
rect 317196 6004 354956 6032
rect 317196 5992 317202 6004
rect 354950 5992 354956 6004
rect 355008 5992 355014 6044
rect 387702 5992 387708 6044
rect 387760 6032 387766 6044
rect 491754 6032 491760 6044
rect 387760 6004 491760 6032
rect 387760 5992 387766 6004
rect 491754 5992 491760 6004
rect 491812 5992 491818 6044
rect 108758 5924 108764 5976
rect 108816 5964 108822 5976
rect 189074 5964 189080 5976
rect 108816 5936 189080 5964
rect 108816 5924 108822 5936
rect 189074 5924 189080 5936
rect 189132 5924 189138 5976
rect 315942 5924 315948 5976
rect 316000 5964 316006 5976
rect 352558 5964 352564 5976
rect 316000 5936 352564 5964
rect 316000 5924 316006 5936
rect 352558 5924 352564 5936
rect 352616 5924 352622 5976
rect 383470 5924 383476 5976
rect 383528 5964 383534 5976
rect 484578 5964 484584 5976
rect 383528 5936 484584 5964
rect 383528 5924 383534 5936
rect 484578 5924 484584 5936
rect 484636 5924 484642 5976
rect 112346 5856 112352 5908
rect 112404 5896 112410 5908
rect 191834 5896 191840 5908
rect 112404 5868 191840 5896
rect 112404 5856 112410 5868
rect 191834 5856 191840 5868
rect 191892 5856 191898 5908
rect 315850 5856 315856 5908
rect 315908 5896 315914 5908
rect 351362 5896 351368 5908
rect 315908 5868 351368 5896
rect 315908 5856 315914 5868
rect 351362 5856 351368 5868
rect 351420 5856 351426 5908
rect 386322 5856 386328 5908
rect 386380 5896 386386 5908
rect 488166 5896 488172 5908
rect 386380 5868 488172 5896
rect 386380 5856 386386 5868
rect 488166 5856 488172 5868
rect 488224 5856 488230 5908
rect 113542 5788 113548 5840
rect 113600 5828 113606 5840
rect 192202 5828 192208 5840
rect 113600 5800 192208 5828
rect 113600 5788 113606 5800
rect 192202 5788 192208 5800
rect 192260 5788 192266 5840
rect 379330 5788 379336 5840
rect 379388 5828 379394 5840
rect 476298 5828 476304 5840
rect 379388 5800 476304 5828
rect 379388 5788 379394 5800
rect 476298 5788 476304 5800
rect 476356 5788 476362 5840
rect 115934 5720 115940 5772
rect 115992 5760 115998 5772
rect 193214 5760 193220 5772
rect 115992 5732 193220 5760
rect 115992 5720 115998 5732
rect 193214 5720 193220 5732
rect 193272 5720 193278 5772
rect 382182 5720 382188 5772
rect 382240 5760 382246 5772
rect 479886 5760 479892 5772
rect 382240 5732 479892 5760
rect 382240 5720 382246 5732
rect 479886 5720 479892 5732
rect 479944 5720 479950 5772
rect 119430 5652 119436 5704
rect 119488 5692 119494 5704
rect 194686 5692 194692 5704
rect 119488 5664 194692 5692
rect 119488 5652 119494 5664
rect 194686 5652 194692 5664
rect 194744 5652 194750 5704
rect 378042 5652 378048 5704
rect 378100 5692 378106 5704
rect 472710 5692 472716 5704
rect 378100 5664 472716 5692
rect 378100 5652 378106 5664
rect 472710 5652 472716 5664
rect 472768 5652 472774 5704
rect 123018 5584 123024 5636
rect 123076 5624 123082 5636
rect 197354 5624 197360 5636
rect 123076 5596 197360 5624
rect 123076 5584 123082 5596
rect 197354 5584 197360 5596
rect 197412 5584 197418 5636
rect 373902 5584 373908 5636
rect 373960 5624 373966 5636
rect 465626 5624 465632 5636
rect 373960 5596 465632 5624
rect 373960 5584 373966 5596
rect 465626 5584 465632 5596
rect 465684 5584 465690 5636
rect 150434 5516 150440 5568
rect 150492 5556 150498 5568
rect 211246 5556 211252 5568
rect 150492 5528 211252 5556
rect 150492 5516 150498 5528
rect 211246 5516 211252 5528
rect 211304 5516 211310 5568
rect 376662 5516 376668 5568
rect 376720 5556 376726 5568
rect 469122 5556 469128 5568
rect 376720 5528 469128 5556
rect 376720 5516 376726 5528
rect 469122 5516 469128 5528
rect 469180 5516 469186 5568
rect 73062 5448 73068 5500
rect 73120 5488 73126 5500
rect 171226 5488 171232 5500
rect 73120 5460 171232 5488
rect 73120 5448 73126 5460
rect 171226 5448 171232 5460
rect 171284 5448 171290 5500
rect 171686 5448 171692 5500
rect 171744 5488 171750 5500
rect 211154 5488 211160 5500
rect 171744 5460 211160 5488
rect 171744 5448 171750 5460
rect 211154 5448 211160 5460
rect 211212 5448 211218 5500
rect 335170 5448 335176 5500
rect 335228 5488 335234 5500
rect 390646 5488 390652 5500
rect 335228 5460 390652 5488
rect 335228 5448 335234 5460
rect 390646 5448 390652 5460
rect 390704 5448 390710 5500
rect 415302 5448 415308 5500
rect 415360 5488 415366 5500
rect 544102 5488 544108 5500
rect 415360 5460 544108 5488
rect 415360 5448 415366 5460
rect 544102 5448 544108 5460
rect 544160 5448 544166 5500
rect 69474 5380 69480 5432
rect 69532 5420 69538 5432
rect 169938 5420 169944 5432
rect 69532 5392 169944 5420
rect 69532 5380 69538 5392
rect 169938 5380 169944 5392
rect 169996 5380 170002 5432
rect 187234 5380 187240 5432
rect 187292 5420 187298 5432
rect 229094 5420 229100 5432
rect 187292 5392 229100 5420
rect 187292 5380 187298 5392
rect 229094 5380 229100 5392
rect 229152 5380 229158 5432
rect 339402 5380 339408 5432
rect 339460 5420 339466 5432
rect 397822 5420 397828 5432
rect 339460 5392 397828 5420
rect 339460 5380 339466 5392
rect 397822 5380 397828 5392
rect 397880 5380 397886 5432
rect 416682 5380 416688 5432
rect 416740 5420 416746 5432
rect 547690 5420 547696 5432
rect 416740 5392 547696 5420
rect 416740 5380 416746 5392
rect 547690 5380 547696 5392
rect 547748 5380 547754 5432
rect 65978 5312 65984 5364
rect 66036 5352 66042 5364
rect 166994 5352 167000 5364
rect 66036 5324 167000 5352
rect 66036 5312 66042 5324
rect 166994 5312 167000 5324
rect 167052 5312 167058 5364
rect 170582 5312 170588 5364
rect 170640 5352 170646 5364
rect 220998 5352 221004 5364
rect 170640 5324 221004 5352
rect 170640 5312 170646 5324
rect 220998 5312 221004 5324
rect 221056 5312 221062 5364
rect 340690 5312 340696 5364
rect 340748 5352 340754 5364
rect 401318 5352 401324 5364
rect 340748 5324 401324 5352
rect 340748 5312 340754 5324
rect 401318 5312 401324 5324
rect 401376 5312 401382 5364
rect 418062 5312 418068 5364
rect 418120 5352 418126 5364
rect 551186 5352 551192 5364
rect 418120 5324 551192 5352
rect 418120 5312 418126 5324
rect 551186 5312 551192 5324
rect 551244 5312 551250 5364
rect 62390 5244 62396 5296
rect 62448 5284 62454 5296
rect 165706 5284 165712 5296
rect 62448 5256 165712 5284
rect 62448 5244 62454 5256
rect 165706 5244 165712 5256
rect 165764 5244 165770 5296
rect 167086 5244 167092 5296
rect 167144 5284 167150 5296
rect 219526 5284 219532 5296
rect 167144 5256 219532 5284
rect 167144 5244 167150 5256
rect 219526 5244 219532 5256
rect 219584 5244 219590 5296
rect 343542 5244 343548 5296
rect 343600 5284 343606 5296
rect 404906 5284 404912 5296
rect 343600 5256 404912 5284
rect 343600 5244 343606 5256
rect 404906 5244 404912 5256
rect 404964 5244 404970 5296
rect 420822 5244 420828 5296
rect 420880 5284 420886 5296
rect 554774 5284 554780 5296
rect 420880 5256 554780 5284
rect 420880 5244 420886 5256
rect 554774 5244 554780 5256
rect 554832 5244 554838 5296
rect 37366 5176 37372 5228
rect 37424 5216 37430 5228
rect 153286 5216 153292 5228
rect 37424 5188 153292 5216
rect 37424 5176 37430 5188
rect 153286 5176 153292 5188
rect 153344 5176 153350 5228
rect 163498 5176 163504 5228
rect 163556 5216 163562 5228
rect 218146 5216 218152 5228
rect 163556 5188 218152 5216
rect 163556 5176 163562 5188
rect 218146 5176 218152 5188
rect 218204 5176 218210 5228
rect 344830 5176 344836 5228
rect 344888 5216 344894 5228
rect 408678 5216 408684 5228
rect 344888 5188 408684 5216
rect 344888 5176 344894 5188
rect 408678 5176 408684 5188
rect 408736 5176 408742 5228
rect 422202 5176 422208 5228
rect 422260 5216 422266 5228
rect 558362 5216 558368 5228
rect 422260 5188 558368 5216
rect 422260 5176 422266 5188
rect 558362 5176 558368 5188
rect 558420 5176 558426 5228
rect 33870 5108 33876 5160
rect 33928 5148 33934 5160
rect 150710 5148 150716 5160
rect 33928 5120 150716 5148
rect 33928 5108 33934 5120
rect 150710 5108 150716 5120
rect 150768 5108 150774 5160
rect 158714 5108 158720 5160
rect 158772 5148 158778 5160
rect 215294 5148 215300 5160
rect 158772 5120 215300 5148
rect 158772 5108 158778 5120
rect 215294 5108 215300 5120
rect 215352 5108 215358 5160
rect 346302 5108 346308 5160
rect 346360 5148 346366 5160
rect 412082 5148 412088 5160
rect 346360 5120 412088 5148
rect 346360 5108 346366 5120
rect 412082 5108 412088 5120
rect 412140 5108 412146 5160
rect 426342 5108 426348 5160
rect 426400 5148 426406 5160
rect 565538 5148 565544 5160
rect 426400 5120 565544 5148
rect 426400 5108 426406 5120
rect 565538 5108 565544 5120
rect 565596 5108 565602 5160
rect 29086 5040 29092 5092
rect 29144 5080 29150 5092
rect 148042 5080 148048 5092
rect 29144 5052 148048 5080
rect 29144 5040 29150 5052
rect 148042 5040 148048 5052
rect 148100 5040 148106 5092
rect 155126 5040 155132 5092
rect 155184 5080 155190 5092
rect 213914 5080 213920 5092
rect 155184 5052 213920 5080
rect 155184 5040 155190 5052
rect 213914 5040 213920 5052
rect 213972 5040 213978 5092
rect 349062 5040 349068 5092
rect 349120 5080 349126 5092
rect 415670 5080 415676 5092
rect 349120 5052 415676 5080
rect 349120 5040 349126 5052
rect 415670 5040 415676 5052
rect 415728 5040 415734 5092
rect 423582 5040 423588 5092
rect 423640 5080 423646 5092
rect 561950 5080 561956 5092
rect 423640 5052 561956 5080
rect 423640 5040 423646 5052
rect 561950 5040 561956 5052
rect 562008 5040 562014 5092
rect 26694 4972 26700 5024
rect 26752 5012 26758 5024
rect 147766 5012 147772 5024
rect 26752 4984 147772 5012
rect 26752 4972 26758 4984
rect 147766 4972 147772 4984
rect 147824 4972 147830 5024
rect 152734 4972 152740 5024
rect 152792 5012 152798 5024
rect 212626 5012 212632 5024
rect 152792 4984 212632 5012
rect 152792 4972 152798 4984
rect 212626 4972 212632 4984
rect 212684 4972 212690 5024
rect 219342 4972 219348 5024
rect 219400 5012 219406 5024
rect 246022 5012 246028 5024
rect 219400 4984 246028 5012
rect 219400 4972 219406 4984
rect 246022 4972 246028 4984
rect 246080 4972 246086 5024
rect 350442 4972 350448 5024
rect 350500 5012 350506 5024
rect 419166 5012 419172 5024
rect 350500 4984 419172 5012
rect 350500 4972 350506 4984
rect 419166 4972 419172 4984
rect 419224 4972 419230 5024
rect 427722 4972 427728 5024
rect 427780 5012 427786 5024
rect 569034 5012 569040 5024
rect 427780 4984 569040 5012
rect 427780 4972 427786 4984
rect 569034 4972 569040 4984
rect 569092 4972 569098 5024
rect 21910 4904 21916 4956
rect 21968 4944 21974 4956
rect 145098 4944 145104 4956
rect 21968 4916 145104 4944
rect 21968 4904 21974 4916
rect 145098 4904 145104 4916
rect 145156 4904 145162 4956
rect 149238 4904 149244 4956
rect 149296 4944 149302 4956
rect 209866 4944 209872 4956
rect 149296 4916 209872 4944
rect 149296 4904 149302 4916
rect 209866 4904 209872 4916
rect 209924 4904 209930 4956
rect 215846 4904 215852 4956
rect 215904 4944 215910 4956
rect 244550 4944 244556 4956
rect 215904 4916 244556 4944
rect 215904 4904 215910 4916
rect 244550 4904 244556 4916
rect 244608 4904 244614 4956
rect 310422 4904 310428 4956
rect 310480 4944 310486 4956
rect 341886 4944 341892 4956
rect 310480 4916 341892 4944
rect 310480 4904 310486 4916
rect 341886 4904 341892 4916
rect 341944 4904 341950 4956
rect 351730 4904 351736 4956
rect 351788 4944 351794 4956
rect 422754 4944 422760 4956
rect 351788 4916 422760 4944
rect 351788 4904 351794 4916
rect 422754 4904 422760 4916
rect 422812 4904 422818 4956
rect 429102 4904 429108 4956
rect 429160 4944 429166 4956
rect 572622 4944 572628 4956
rect 429160 4916 572628 4944
rect 429160 4904 429166 4916
rect 572622 4904 572628 4916
rect 572680 4904 572686 4956
rect 12434 4836 12440 4888
rect 12492 4876 12498 4888
rect 139394 4876 139400 4888
rect 12492 4848 139400 4876
rect 12492 4836 12498 4848
rect 139394 4836 139400 4848
rect 139452 4836 139458 4888
rect 142062 4836 142068 4888
rect 142120 4876 142126 4888
rect 207014 4876 207020 4888
rect 142120 4848 207020 4876
rect 142120 4836 142126 4848
rect 207014 4836 207020 4848
rect 207072 4836 207078 4888
rect 212258 4836 212264 4888
rect 212316 4876 212322 4888
rect 242986 4876 242992 4888
rect 212316 4848 242992 4876
rect 212316 4836 212322 4848
rect 242986 4836 242992 4848
rect 243044 4836 243050 4888
rect 314562 4836 314568 4888
rect 314620 4876 314626 4888
rect 349062 4876 349068 4888
rect 314620 4848 349068 4876
rect 314620 4836 314626 4848
rect 349062 4836 349068 4848
rect 349120 4836 349126 4888
rect 354582 4836 354588 4888
rect 354640 4876 354646 4888
rect 426342 4876 426348 4888
rect 354640 4848 426348 4876
rect 354640 4836 354646 4848
rect 426342 4836 426348 4848
rect 426400 4836 426406 4888
rect 431862 4836 431868 4888
rect 431920 4876 431926 4888
rect 576210 4876 576216 4888
rect 431920 4848 576216 4876
rect 431920 4836 431926 4848
rect 576210 4836 576216 4848
rect 576268 4836 576274 4888
rect 17218 4768 17224 4820
rect 17276 4808 17282 4820
rect 142246 4808 142252 4820
rect 17276 4780 142252 4808
rect 17276 4768 17282 4780
rect 142246 4768 142252 4780
rect 142304 4768 142310 4820
rect 145650 4768 145656 4820
rect 145708 4808 145714 4820
rect 208394 4808 208400 4820
rect 145708 4780 208400 4808
rect 145708 4768 145714 4780
rect 208394 4768 208400 4780
rect 208452 4768 208458 4820
rect 208670 4768 208676 4820
rect 208728 4808 208734 4820
rect 240134 4808 240140 4820
rect 208728 4780 240140 4808
rect 208728 4768 208734 4780
rect 240134 4768 240140 4780
rect 240192 4768 240198 4820
rect 313090 4768 313096 4820
rect 313148 4808 313154 4820
rect 347866 4808 347872 4820
rect 313148 4780 347872 4808
rect 313148 4768 313154 4780
rect 347866 4768 347872 4780
rect 347924 4768 347930 4820
rect 355962 4768 355968 4820
rect 356020 4808 356026 4820
rect 429930 4808 429936 4820
rect 356020 4780 429936 4808
rect 356020 4768 356026 4780
rect 429930 4768 429936 4780
rect 429988 4768 429994 4820
rect 433242 4768 433248 4820
rect 433300 4808 433306 4820
rect 579798 4808 579804 4820
rect 433300 4780 579804 4808
rect 433300 4768 433306 4780
rect 579798 4768 579804 4780
rect 579856 4768 579862 4820
rect 76650 4700 76656 4752
rect 76708 4740 76714 4752
rect 172514 4740 172520 4752
rect 76708 4712 172520 4740
rect 76708 4700 76714 4712
rect 172514 4700 172520 4712
rect 172572 4700 172578 4752
rect 203794 4700 203800 4752
rect 203852 4740 203858 4752
rect 237466 4740 237472 4752
rect 203852 4712 237472 4740
rect 203852 4700 203858 4712
rect 237466 4700 237472 4712
rect 237524 4700 237530 4752
rect 338022 4700 338028 4752
rect 338080 4740 338086 4752
rect 394234 4740 394240 4752
rect 338080 4712 394240 4740
rect 338080 4700 338086 4712
rect 394234 4700 394240 4712
rect 394292 4700 394298 4752
rect 412542 4700 412548 4752
rect 412600 4740 412606 4752
rect 540514 4740 540520 4752
rect 412600 4712 540520 4740
rect 412600 4700 412606 4712
rect 540514 4700 540520 4712
rect 540572 4700 540578 4752
rect 80238 4632 80244 4684
rect 80296 4672 80302 4684
rect 175550 4672 175556 4684
rect 80296 4644 175556 4672
rect 80296 4632 80302 4644
rect 175550 4632 175556 4644
rect 175608 4632 175614 4684
rect 205082 4632 205088 4684
rect 205140 4672 205146 4684
rect 238938 4672 238944 4684
rect 205140 4644 238944 4672
rect 205140 4632 205146 4644
rect 238938 4632 238944 4644
rect 238996 4632 239002 4684
rect 333790 4632 333796 4684
rect 333848 4672 333854 4684
rect 387058 4672 387064 4684
rect 333848 4644 387064 4672
rect 333848 4632 333854 4644
rect 387058 4632 387064 4644
rect 387116 4632 387122 4684
rect 411162 4632 411168 4684
rect 411220 4672 411226 4684
rect 536926 4672 536932 4684
rect 411220 4644 536932 4672
rect 411220 4632 411226 4644
rect 536926 4632 536932 4644
rect 536984 4632 536990 4684
rect 83826 4564 83832 4616
rect 83884 4604 83890 4616
rect 176746 4604 176752 4616
rect 83884 4576 176752 4604
rect 83884 4564 83890 4576
rect 176746 4564 176752 4576
rect 176804 4564 176810 4616
rect 204162 4564 204168 4616
rect 204220 4604 204226 4616
rect 234614 4604 234620 4616
rect 204220 4576 234620 4604
rect 204220 4564 204226 4576
rect 234614 4564 234620 4576
rect 234672 4564 234678 4616
rect 332502 4564 332508 4616
rect 332560 4604 332566 4616
rect 383562 4604 383568 4616
rect 332560 4576 383568 4604
rect 332560 4564 332566 4576
rect 383562 4564 383568 4576
rect 383620 4564 383626 4616
rect 409782 4564 409788 4616
rect 409840 4604 409846 4616
rect 533430 4604 533436 4616
rect 409840 4576 533436 4604
rect 409840 4564 409846 4576
rect 533430 4564 533436 4576
rect 533488 4564 533494 4616
rect 87322 4496 87328 4548
rect 87380 4536 87386 4548
rect 178034 4536 178040 4548
rect 87380 4508 178040 4536
rect 87380 4496 87386 4508
rect 178034 4496 178040 4508
rect 178092 4496 178098 4548
rect 329742 4496 329748 4548
rect 329800 4536 329806 4548
rect 379974 4536 379980 4548
rect 329800 4508 379980 4536
rect 329800 4496 329806 4508
rect 379974 4496 379980 4508
rect 380032 4496 380038 4548
rect 406930 4496 406936 4548
rect 406988 4536 406994 4548
rect 529842 4536 529848 4548
rect 406988 4508 529848 4536
rect 406988 4496 406994 4508
rect 529842 4496 529848 4508
rect 529900 4496 529906 4548
rect 49326 4428 49332 4480
rect 49384 4468 49390 4480
rect 130378 4468 130384 4480
rect 49384 4440 130384 4468
rect 49384 4428 49390 4440
rect 130378 4428 130384 4440
rect 130436 4428 130442 4480
rect 138474 4428 138480 4480
rect 138532 4468 138538 4480
rect 204254 4468 204260 4480
rect 138532 4440 204260 4468
rect 138532 4428 138538 4440
rect 204254 4428 204260 4440
rect 204312 4428 204318 4480
rect 328270 4428 328276 4480
rect 328328 4468 328334 4480
rect 376386 4468 376392 4480
rect 328328 4440 376392 4468
rect 328328 4428 328334 4440
rect 376386 4428 376392 4440
rect 376444 4428 376450 4480
rect 405642 4428 405648 4480
rect 405700 4468 405706 4480
rect 526254 4468 526260 4480
rect 405700 4440 526260 4468
rect 405700 4428 405706 4440
rect 526254 4428 526260 4440
rect 526312 4428 526318 4480
rect 52822 4360 52828 4412
rect 52880 4400 52886 4412
rect 122098 4400 122104 4412
rect 52880 4372 122104 4400
rect 52880 4360 52886 4372
rect 122098 4360 122104 4372
rect 122156 4360 122162 4412
rect 124214 4360 124220 4412
rect 124272 4400 124278 4412
rect 125962 4400 125968 4412
rect 124272 4372 125968 4400
rect 124272 4360 124278 4372
rect 125962 4360 125968 4372
rect 126020 4360 126026 4412
rect 214006 4400 214012 4412
rect 162872 4372 214012 4400
rect 63586 4292 63592 4344
rect 63644 4332 63650 4344
rect 128814 4332 128820 4344
rect 63644 4304 128820 4332
rect 63644 4292 63650 4304
rect 128814 4292 128820 4304
rect 128872 4292 128878 4344
rect 70670 4224 70676 4276
rect 70728 4264 70734 4276
rect 120718 4264 120724 4276
rect 70728 4236 120724 4264
rect 70728 4224 70734 4236
rect 120718 4224 120724 4236
rect 120776 4224 120782 4276
rect 123478 4224 123484 4276
rect 123536 4224 123542 4276
rect 109954 4156 109960 4208
rect 110012 4196 110018 4208
rect 123496 4196 123524 4224
rect 110012 4168 123524 4196
rect 148980 4168 149192 4196
rect 110012 4156 110018 4168
rect 46934 4088 46940 4140
rect 46992 4128 46998 4140
rect 55217 4131 55275 4137
rect 55217 4128 55229 4131
rect 46992 4100 55229 4128
rect 46992 4088 46998 4100
rect 55217 4097 55229 4100
rect 55263 4097 55275 4131
rect 55217 4091 55275 4097
rect 64785 4131 64843 4137
rect 64785 4097 64797 4131
rect 64831 4128 64843 4131
rect 74537 4131 74595 4137
rect 74537 4128 74549 4131
rect 64831 4100 74549 4128
rect 64831 4097 64843 4100
rect 64785 4091 64843 4097
rect 74537 4097 74549 4100
rect 74583 4097 74595 4131
rect 74537 4091 74595 4097
rect 84105 4131 84163 4137
rect 84105 4097 84117 4131
rect 84151 4128 84163 4131
rect 93857 4131 93915 4137
rect 93857 4128 93869 4131
rect 84151 4100 93869 4128
rect 84151 4097 84163 4100
rect 84105 4091 84163 4097
rect 93857 4097 93869 4100
rect 93903 4097 93915 4131
rect 93857 4091 93915 4097
rect 103425 4131 103483 4137
rect 103425 4097 103437 4131
rect 103471 4128 103483 4131
rect 113177 4131 113235 4137
rect 113177 4128 113189 4131
rect 103471 4100 113189 4128
rect 103471 4097 103483 4100
rect 103425 4091 103483 4097
rect 113177 4097 113189 4100
rect 113223 4097 113235 4131
rect 113177 4091 113235 4097
rect 123481 4131 123539 4137
rect 123481 4097 123493 4131
rect 123527 4128 123539 4131
rect 133141 4131 133199 4137
rect 133141 4128 133153 4131
rect 123527 4100 133153 4128
rect 123527 4097 123539 4100
rect 123481 4091 123539 4097
rect 133141 4097 133153 4100
rect 133187 4097 133199 4131
rect 133141 4091 133199 4097
rect 142801 4131 142859 4137
rect 142801 4097 142813 4131
rect 142847 4128 142859 4131
rect 148873 4131 148931 4137
rect 148873 4128 148885 4131
rect 142847 4100 148885 4128
rect 142847 4097 142859 4100
rect 142801 4091 142859 4097
rect 148873 4097 148885 4100
rect 148919 4097 148931 4131
rect 148873 4091 148931 4097
rect 39758 4020 39764 4072
rect 39816 4060 39822 4072
rect 148980 4060 149008 4168
rect 149164 4128 149192 4168
rect 153194 4128 153200 4140
rect 149164 4100 153200 4128
rect 153194 4088 153200 4100
rect 153252 4088 153258 4140
rect 156322 4088 156328 4140
rect 156380 4128 156386 4140
rect 162872 4128 162900 4372
rect 214006 4360 214012 4372
rect 214064 4360 214070 4412
rect 326982 4360 326988 4412
rect 327040 4400 327046 4412
rect 372798 4400 372804 4412
rect 327040 4372 372804 4400
rect 327040 4360 327046 4372
rect 372798 4360 372804 4372
rect 372856 4360 372862 4412
rect 401502 4360 401508 4412
rect 401560 4400 401566 4412
rect 519078 4400 519084 4412
rect 401560 4372 519084 4400
rect 401560 4360 401566 4372
rect 519078 4360 519084 4372
rect 519136 4360 519142 4412
rect 165614 4292 165620 4344
rect 165672 4332 165678 4344
rect 215570 4332 215576 4344
rect 165672 4304 215576 4332
rect 165672 4292 165678 4304
rect 215570 4292 215576 4304
rect 215628 4292 215634 4344
rect 324130 4292 324136 4344
rect 324188 4332 324194 4344
rect 369210 4332 369216 4344
rect 324188 4304 369216 4332
rect 324188 4292 324194 4304
rect 369210 4292 369216 4304
rect 369268 4292 369274 4344
rect 404262 4292 404268 4344
rect 404320 4332 404326 4344
rect 522666 4332 522672 4344
rect 404320 4304 522672 4332
rect 404320 4292 404326 4304
rect 522666 4292 522672 4304
rect 522724 4292 522730 4344
rect 168282 4224 168288 4276
rect 168340 4264 168346 4276
rect 208486 4264 208492 4276
rect 168340 4236 208492 4264
rect 168340 4224 168346 4236
rect 208486 4224 208492 4236
rect 208544 4224 208550 4276
rect 322566 4224 322572 4276
rect 322624 4264 322630 4276
rect 365714 4264 365720 4276
rect 322624 4236 365720 4264
rect 322624 4224 322630 4236
rect 365714 4224 365720 4236
rect 365772 4224 365778 4276
rect 400030 4224 400036 4276
rect 400088 4264 400094 4276
rect 515582 4264 515588 4276
rect 400088 4236 515588 4264
rect 400088 4224 400094 4236
rect 515582 4224 515588 4236
rect 515640 4224 515646 4276
rect 321370 4156 321376 4208
rect 321428 4196 321434 4208
rect 362126 4196 362132 4208
rect 321428 4168 362132 4196
rect 321428 4156 321434 4168
rect 362126 4156 362132 4168
rect 362184 4156 362190 4208
rect 398742 4156 398748 4208
rect 398800 4196 398806 4208
rect 511994 4196 512000 4208
rect 398800 4168 512000 4196
rect 398800 4156 398806 4168
rect 511994 4156 512000 4168
rect 512052 4156 512058 4208
rect 156380 4100 162900 4128
rect 156380 4088 156386 4100
rect 171778 4088 171784 4140
rect 171836 4128 171842 4140
rect 174538 4128 174544 4140
rect 171836 4100 174544 4128
rect 171836 4088 171842 4100
rect 174538 4088 174544 4100
rect 174596 4088 174602 4140
rect 177758 4088 177764 4140
rect 177816 4128 177822 4140
rect 185670 4128 185676 4140
rect 177816 4100 185676 4128
rect 177816 4088 177822 4100
rect 185670 4088 185676 4100
rect 185728 4088 185734 4140
rect 189626 4088 189632 4140
rect 189684 4128 189690 4140
rect 190362 4128 190368 4140
rect 189684 4100 190368 4128
rect 189684 4088 189690 4100
rect 190362 4088 190368 4100
rect 190420 4088 190426 4140
rect 190822 4088 190828 4140
rect 190880 4128 190886 4140
rect 190880 4100 225092 4128
rect 190880 4088 190886 4100
rect 39816 4032 149008 4060
rect 149057 4063 149115 4069
rect 39816 4020 39822 4032
rect 149057 4029 149069 4063
rect 149103 4060 149115 4063
rect 157334 4060 157340 4072
rect 149103 4032 157340 4060
rect 149103 4029 149115 4032
rect 149057 4023 149115 4029
rect 157334 4020 157340 4032
rect 157392 4020 157398 4072
rect 170398 4060 170404 4072
rect 168116 4032 170404 4060
rect 34974 3952 34980 4004
rect 35032 3992 35038 4004
rect 151906 3992 151912 4004
rect 35032 3964 151912 3992
rect 35032 3952 35038 3964
rect 151906 3952 151912 3964
rect 151964 3952 151970 4004
rect 161106 3952 161112 4004
rect 161164 3992 161170 4004
rect 168116 3992 168144 4032
rect 170398 4020 170404 4032
rect 170456 4020 170462 4072
rect 174170 4020 174176 4072
rect 174228 4060 174234 4072
rect 185578 4060 185584 4072
rect 174228 4032 185584 4060
rect 174228 4020 174234 4032
rect 185578 4020 185584 4032
rect 185636 4020 185642 4072
rect 188430 4020 188436 4072
rect 188488 4060 188494 4072
rect 218057 4063 218115 4069
rect 218057 4060 218069 4063
rect 188488 4032 218069 4060
rect 188488 4020 188494 4032
rect 218057 4029 218069 4032
rect 218103 4029 218115 4063
rect 218057 4023 218115 4029
rect 218146 4020 218152 4072
rect 218204 4060 218210 4072
rect 219250 4060 219256 4072
rect 218204 4032 219256 4060
rect 218204 4020 218210 4032
rect 219250 4020 219256 4032
rect 219308 4020 219314 4072
rect 222930 4020 222936 4072
rect 222988 4060 222994 4072
rect 223482 4060 223488 4072
rect 222988 4032 223488 4060
rect 222988 4020 222994 4032
rect 223482 4020 223488 4032
rect 223540 4020 223546 4072
rect 225064 4060 225092 4100
rect 226518 4088 226524 4140
rect 226576 4128 226582 4140
rect 227622 4128 227628 4140
rect 226576 4100 227628 4128
rect 226576 4088 226582 4100
rect 227622 4088 227628 4100
rect 227680 4088 227686 4140
rect 227714 4088 227720 4140
rect 227772 4128 227778 4140
rect 229002 4128 229008 4140
rect 227772 4100 229008 4128
rect 227772 4088 227778 4100
rect 229002 4088 229008 4100
rect 229060 4088 229066 4140
rect 231302 4088 231308 4140
rect 231360 4128 231366 4140
rect 231762 4128 231768 4140
rect 231360 4100 231768 4128
rect 231360 4088 231366 4100
rect 231762 4088 231768 4100
rect 231820 4088 231826 4140
rect 232498 4088 232504 4140
rect 232556 4128 232562 4140
rect 233142 4128 233148 4140
rect 232556 4100 233148 4128
rect 232556 4088 232562 4100
rect 233142 4088 233148 4100
rect 233200 4088 233206 4140
rect 233694 4088 233700 4140
rect 233752 4128 233758 4140
rect 234522 4128 234528 4140
rect 233752 4100 234528 4128
rect 233752 4088 233758 4100
rect 234522 4088 234528 4100
rect 234580 4088 234586 4140
rect 235994 4088 236000 4140
rect 236052 4128 236058 4140
rect 237190 4128 237196 4140
rect 236052 4100 237196 4128
rect 236052 4088 236058 4100
rect 237190 4088 237196 4100
rect 237248 4088 237254 4140
rect 239582 4088 239588 4140
rect 239640 4128 239646 4140
rect 240042 4128 240048 4140
rect 239640 4100 240048 4128
rect 239640 4088 239646 4100
rect 240042 4088 240048 4100
rect 240100 4088 240106 4140
rect 240778 4088 240784 4140
rect 240836 4128 240842 4140
rect 241422 4128 241428 4140
rect 240836 4100 241428 4128
rect 240836 4088 240842 4100
rect 241422 4088 241428 4100
rect 241480 4088 241486 4140
rect 243170 4088 243176 4140
rect 243228 4128 243234 4140
rect 244182 4128 244188 4140
rect 243228 4100 244188 4128
rect 243228 4088 243234 4100
rect 244182 4088 244188 4100
rect 244240 4088 244246 4140
rect 251450 4088 251456 4140
rect 251508 4128 251514 4140
rect 252462 4128 252468 4140
rect 251508 4100 252468 4128
rect 251508 4088 251514 4100
rect 252462 4088 252468 4100
rect 252520 4088 252526 4140
rect 265802 4088 265808 4140
rect 265860 4128 265866 4140
rect 266262 4128 266268 4140
rect 265860 4100 266268 4128
rect 265860 4088 265866 4100
rect 266262 4088 266268 4100
rect 266320 4088 266326 4140
rect 268102 4088 268108 4140
rect 268160 4128 268166 4140
rect 269758 4128 269764 4140
rect 268160 4100 269764 4128
rect 268160 4088 268166 4100
rect 269758 4088 269764 4100
rect 269816 4088 269822 4140
rect 271690 4088 271696 4140
rect 271748 4128 271754 4140
rect 272518 4128 272524 4140
rect 271748 4100 272524 4128
rect 271748 4088 271754 4100
rect 272518 4088 272524 4100
rect 272576 4088 272582 4140
rect 274082 4088 274088 4140
rect 274140 4128 274146 4140
rect 274542 4128 274548 4140
rect 274140 4100 274548 4128
rect 274140 4088 274146 4100
rect 274542 4088 274548 4100
rect 274600 4088 274606 4140
rect 280062 4088 280068 4140
rect 280120 4128 280126 4140
rect 282454 4128 282460 4140
rect 280120 4100 282460 4128
rect 280120 4088 280126 4100
rect 282454 4088 282460 4100
rect 282512 4088 282518 4140
rect 284938 4088 284944 4140
rect 284996 4128 285002 4140
rect 288342 4128 288348 4140
rect 284996 4100 288348 4128
rect 284996 4088 285002 4100
rect 288342 4088 288348 4100
rect 288400 4088 288406 4140
rect 292390 4088 292396 4140
rect 292448 4128 292454 4140
rect 307386 4128 307392 4140
rect 292448 4100 307392 4128
rect 292448 4088 292454 4100
rect 307386 4088 307392 4100
rect 307444 4088 307450 4140
rect 315298 4088 315304 4140
rect 315356 4128 315362 4140
rect 315850 4128 315856 4140
rect 315356 4100 315856 4128
rect 315356 4088 315362 4100
rect 315850 4088 315856 4100
rect 315908 4088 315914 4140
rect 321462 4088 321468 4140
rect 321520 4128 321526 4140
rect 321520 4100 355456 4128
rect 321520 4088 321526 4100
rect 231946 4060 231952 4072
rect 225064 4032 231952 4060
rect 231946 4020 231952 4032
rect 232004 4020 232010 4072
rect 241974 4020 241980 4072
rect 242032 4060 242038 4072
rect 243538 4060 243544 4072
rect 242032 4032 243544 4060
rect 242032 4020 242038 4032
rect 243538 4020 243544 4032
rect 243596 4020 243602 4072
rect 283558 4020 283564 4072
rect 283616 4060 283622 4072
rect 287146 4060 287152 4072
rect 283616 4032 287152 4060
rect 283616 4020 283622 4032
rect 287146 4020 287152 4032
rect 287204 4020 287210 4072
rect 297910 4020 297916 4072
rect 297968 4020 297974 4072
rect 298002 4020 298008 4072
rect 298060 4060 298066 4072
rect 316954 4060 316960 4072
rect 298060 4032 316960 4060
rect 298060 4020 298066 4032
rect 316954 4020 316960 4032
rect 317012 4020 317018 4072
rect 324222 4020 324228 4072
rect 324280 4060 324286 4072
rect 355321 4063 355379 4069
rect 355321 4060 355333 4063
rect 324280 4032 355333 4060
rect 324280 4020 324286 4032
rect 355321 4029 355333 4032
rect 355367 4029 355379 4063
rect 355321 4023 355379 4029
rect 161164 3964 168144 3992
rect 161164 3952 161170 3964
rect 168190 3952 168196 4004
rect 168248 3992 168254 4004
rect 176010 3992 176016 4004
rect 168248 3964 176016 3992
rect 168248 3952 168254 3964
rect 176010 3952 176016 3964
rect 176068 3952 176074 4004
rect 183738 3952 183744 4004
rect 183796 3992 183802 4004
rect 227806 3992 227812 4004
rect 183796 3964 227812 3992
rect 183796 3952 183802 3964
rect 227806 3952 227812 3964
rect 227864 3952 227870 4004
rect 269298 3952 269304 4004
rect 269356 3992 269362 4004
rect 272150 3992 272156 4004
rect 269356 3964 272156 3992
rect 269356 3952 269362 3964
rect 272150 3952 272156 3964
rect 272208 3952 272214 4004
rect 293126 3992 293132 4004
rect 287348 3964 293132 3992
rect 32674 3884 32680 3936
rect 32732 3924 32738 3936
rect 150618 3924 150624 3936
rect 32732 3896 150624 3924
rect 32732 3884 32738 3896
rect 150618 3884 150624 3896
rect 150676 3884 150682 3936
rect 164694 3884 164700 3936
rect 164752 3924 164758 3936
rect 175918 3924 175924 3936
rect 164752 3896 175924 3924
rect 164752 3884 164758 3896
rect 175918 3884 175924 3896
rect 175976 3884 175982 3936
rect 180150 3884 180156 3936
rect 180208 3924 180214 3936
rect 226426 3924 226432 3936
rect 180208 3896 226432 3924
rect 180208 3884 180214 3896
rect 226426 3884 226432 3896
rect 226484 3884 226490 3936
rect 229741 3927 229799 3933
rect 229741 3893 229753 3927
rect 229787 3924 229799 3927
rect 236638 3924 236644 3936
rect 229787 3896 236644 3924
rect 229787 3893 229799 3896
rect 229741 3887 229799 3893
rect 236638 3884 236644 3896
rect 236696 3884 236702 3936
rect 285582 3884 285588 3936
rect 285640 3924 285646 3936
rect 287348 3924 287376 3964
rect 293126 3952 293132 3964
rect 293184 3952 293190 4004
rect 297928 3992 297956 4020
rect 318058 3992 318064 4004
rect 297928 3964 318064 3992
rect 318058 3952 318064 3964
rect 318116 3952 318122 4004
rect 322842 3952 322848 4004
rect 322900 3992 322906 4004
rect 355229 3995 355287 4001
rect 355229 3992 355241 3995
rect 322900 3964 355241 3992
rect 322900 3952 322906 3964
rect 355229 3961 355241 3964
rect 355275 3961 355287 3995
rect 355428 3992 355456 4100
rect 358078 4088 358084 4140
rect 358136 4128 358142 4140
rect 360930 4128 360936 4140
rect 358136 4100 360936 4128
rect 358136 4088 358142 4100
rect 360930 4088 360936 4100
rect 360988 4088 360994 4140
rect 363598 4088 363604 4140
rect 363656 4128 363662 4140
rect 364518 4128 364524 4140
rect 363656 4100 364524 4128
rect 363656 4088 363662 4100
rect 364518 4088 364524 4100
rect 364576 4088 364582 4140
rect 391750 4088 391756 4140
rect 391808 4128 391814 4140
rect 500126 4128 500132 4140
rect 391808 4100 500132 4128
rect 391808 4088 391814 4100
rect 500126 4088 500132 4100
rect 500184 4088 500190 4140
rect 500218 4088 500224 4140
rect 500276 4128 500282 4140
rect 504545 4131 504603 4137
rect 504545 4128 504557 4131
rect 500276 4100 504557 4128
rect 500276 4088 500282 4100
rect 504545 4097 504557 4100
rect 504591 4097 504603 4131
rect 504545 4091 504603 4097
rect 507118 4088 507124 4140
rect 507176 4128 507182 4140
rect 571426 4128 571432 4140
rect 507176 4100 571432 4128
rect 507176 4088 507182 4100
rect 571426 4088 571432 4100
rect 571484 4088 571490 4140
rect 355505 4063 355563 4069
rect 355505 4029 355517 4063
rect 355551 4060 355563 4063
rect 368014 4060 368020 4072
rect 355551 4032 368020 4060
rect 355551 4029 355563 4032
rect 355505 4023 355563 4029
rect 368014 4020 368020 4032
rect 368072 4020 368078 4072
rect 395982 4020 395988 4072
rect 396040 4060 396046 4072
rect 507210 4060 507216 4072
rect 396040 4032 507216 4060
rect 396040 4020 396046 4032
rect 507210 4020 507216 4032
rect 507268 4020 507274 4072
rect 511258 4020 511264 4072
rect 511316 4060 511322 4072
rect 578602 4060 578608 4072
rect 511316 4032 578608 4060
rect 511316 4020 511322 4032
rect 578602 4020 578608 4032
rect 578660 4020 578666 4072
rect 363322 3992 363328 4004
rect 355428 3964 363328 3992
rect 355229 3955 355287 3961
rect 363322 3952 363328 3964
rect 363380 3952 363386 4004
rect 400122 3952 400128 4004
rect 400180 3992 400186 4004
rect 514386 3992 514392 4004
rect 400180 3964 514392 3992
rect 400180 3952 400186 3964
rect 514386 3952 514392 3964
rect 514444 3952 514450 4004
rect 285640 3896 287376 3924
rect 285640 3884 285646 3896
rect 288250 3884 288256 3936
rect 288308 3924 288314 3936
rect 297910 3924 297916 3936
rect 288308 3896 297916 3924
rect 288308 3884 288314 3896
rect 297910 3884 297916 3896
rect 297968 3884 297974 3936
rect 302142 3884 302148 3936
rect 302200 3924 302206 3936
rect 324038 3924 324044 3936
rect 302200 3896 324044 3924
rect 302200 3884 302206 3896
rect 324038 3884 324044 3896
rect 324096 3884 324102 3936
rect 326338 3884 326344 3936
rect 326396 3924 326402 3936
rect 370406 3924 370412 3936
rect 326396 3896 370412 3924
rect 326396 3884 326402 3896
rect 370406 3884 370412 3896
rect 370464 3884 370470 3936
rect 374638 3884 374644 3936
rect 374696 3924 374702 3936
rect 374696 3896 375420 3924
rect 374696 3884 374702 3896
rect 25498 3816 25504 3868
rect 25556 3856 25562 3868
rect 146386 3856 146392 3868
rect 25556 3828 146392 3856
rect 25556 3816 25562 3828
rect 146386 3816 146392 3828
rect 146444 3816 146450 3868
rect 153930 3816 153936 3868
rect 153988 3856 153994 3868
rect 171502 3856 171508 3868
rect 153988 3828 171508 3856
rect 153988 3816 153994 3828
rect 171502 3816 171508 3828
rect 171560 3816 171566 3868
rect 176562 3816 176568 3868
rect 176620 3856 176626 3868
rect 217873 3859 217931 3865
rect 217873 3856 217885 3859
rect 176620 3828 217885 3856
rect 176620 3816 176626 3828
rect 217873 3825 217885 3828
rect 217919 3825 217931 3859
rect 222378 3856 222384 3868
rect 217873 3819 217931 3825
rect 217980 3828 222384 3856
rect 24302 3748 24308 3800
rect 24360 3788 24366 3800
rect 146294 3788 146300 3800
rect 24360 3760 146300 3788
rect 24360 3748 24366 3760
rect 146294 3748 146300 3760
rect 146352 3748 146358 3800
rect 151538 3748 151544 3800
rect 151596 3788 151602 3800
rect 171686 3788 171692 3800
rect 151596 3760 171692 3788
rect 151596 3748 151602 3760
rect 171686 3748 171692 3760
rect 171744 3748 171750 3800
rect 172974 3748 172980 3800
rect 173032 3788 173038 3800
rect 217980 3788 218008 3828
rect 222378 3816 222384 3828
rect 222436 3816 222442 3868
rect 225233 3859 225291 3865
rect 225233 3825 225245 3859
rect 225279 3856 225291 3859
rect 233418 3856 233424 3868
rect 225279 3828 233424 3856
rect 225279 3825 225291 3828
rect 225233 3819 225291 3825
rect 233418 3816 233424 3828
rect 233476 3816 233482 3868
rect 286962 3816 286968 3868
rect 287020 3856 287026 3868
rect 295518 3856 295524 3868
rect 287020 3828 295524 3856
rect 287020 3816 287026 3828
rect 295518 3816 295524 3828
rect 295576 3816 295582 3868
rect 299382 3816 299388 3868
rect 299440 3856 299446 3868
rect 320450 3856 320456 3868
rect 299440 3828 320456 3856
rect 299440 3816 299446 3828
rect 320450 3816 320456 3828
rect 320508 3816 320514 3868
rect 328362 3816 328368 3868
rect 328420 3856 328426 3868
rect 375190 3856 375196 3868
rect 328420 3828 375196 3856
rect 328420 3816 328426 3828
rect 375190 3816 375196 3828
rect 375248 3816 375254 3868
rect 375392 3856 375420 3896
rect 402882 3884 402888 3936
rect 402940 3924 402946 3936
rect 521470 3924 521476 3936
rect 402940 3896 521476 3924
rect 402940 3884 402946 3896
rect 521470 3884 521476 3896
rect 521528 3884 521534 3936
rect 393038 3856 393044 3868
rect 375392 3828 393044 3856
rect 393038 3816 393044 3828
rect 393096 3816 393102 3868
rect 398837 3859 398895 3865
rect 398837 3825 398849 3859
rect 398883 3856 398895 3859
rect 398883 3828 403848 3856
rect 398883 3825 398895 3828
rect 398837 3819 398895 3825
rect 173032 3760 218008 3788
rect 218057 3791 218115 3797
rect 173032 3748 173038 3760
rect 218057 3757 218069 3791
rect 218103 3788 218115 3791
rect 230566 3788 230572 3800
rect 218103 3760 230572 3788
rect 218103 3757 218115 3760
rect 218057 3751 218115 3757
rect 230566 3748 230572 3760
rect 230624 3748 230630 3800
rect 234798 3748 234804 3800
rect 234856 3788 234862 3800
rect 250438 3788 250444 3800
rect 234856 3760 250444 3788
rect 234856 3748 234862 3760
rect 250438 3748 250444 3760
rect 250496 3748 250502 3800
rect 288066 3748 288072 3800
rect 288124 3788 288130 3800
rect 299106 3788 299112 3800
rect 288124 3760 299112 3788
rect 288124 3748 288130 3760
rect 299106 3748 299112 3760
rect 299164 3748 299170 3800
rect 302050 3748 302056 3800
rect 302108 3788 302114 3800
rect 325234 3788 325240 3800
rect 302108 3760 325240 3788
rect 302108 3748 302114 3760
rect 325234 3748 325240 3760
rect 325292 3748 325298 3800
rect 326154 3748 326160 3800
rect 326212 3788 326218 3800
rect 326433 3791 326491 3797
rect 326433 3788 326445 3791
rect 326212 3760 326445 3788
rect 326212 3748 326218 3760
rect 326433 3757 326445 3760
rect 326479 3757 326491 3791
rect 326433 3751 326491 3757
rect 334618 3748 334624 3800
rect 334676 3788 334682 3800
rect 335906 3788 335912 3800
rect 334676 3760 335912 3788
rect 334676 3748 334682 3760
rect 335906 3748 335912 3760
rect 335964 3748 335970 3800
rect 385862 3788 385868 3800
rect 340156 3760 385868 3788
rect 19518 3680 19524 3732
rect 19576 3720 19582 3732
rect 143534 3720 143540 3732
rect 19576 3692 143540 3720
rect 19576 3680 19582 3692
rect 143534 3680 143540 3692
rect 143592 3680 143598 3732
rect 146846 3680 146852 3732
rect 146904 3720 146910 3732
rect 168282 3720 168288 3732
rect 146904 3692 168288 3720
rect 146904 3680 146910 3692
rect 168282 3680 168288 3692
rect 168340 3680 168346 3732
rect 169386 3680 169392 3732
rect 169444 3720 169450 3732
rect 220814 3720 220820 3732
rect 169444 3692 220820 3720
rect 169444 3680 169450 3692
rect 220814 3680 220820 3692
rect 220872 3680 220878 3732
rect 221734 3680 221740 3732
rect 221792 3720 221798 3732
rect 240686 3720 240692 3732
rect 221792 3692 240692 3720
rect 221792 3680 221798 3692
rect 240686 3680 240692 3692
rect 240744 3680 240750 3732
rect 286870 3680 286876 3732
rect 286928 3720 286934 3732
rect 296714 3720 296720 3732
rect 286928 3692 296720 3720
rect 286928 3680 286934 3692
rect 296714 3680 296720 3692
rect 296772 3680 296778 3732
rect 303522 3680 303528 3732
rect 303580 3720 303586 3732
rect 327626 3720 327632 3732
rect 303580 3692 327632 3720
rect 303580 3680 303586 3692
rect 327626 3680 327632 3692
rect 327684 3680 327690 3732
rect 333882 3680 333888 3732
rect 333940 3720 333946 3732
rect 340156 3720 340184 3760
rect 385862 3748 385868 3760
rect 385920 3748 385926 3800
rect 389818 3748 389824 3800
rect 389876 3788 389882 3800
rect 403710 3788 403716 3800
rect 389876 3760 403716 3788
rect 389876 3748 389882 3760
rect 403710 3748 403716 3760
rect 403768 3748 403774 3800
rect 403820 3788 403848 3828
rect 407022 3816 407028 3868
rect 407080 3856 407086 3868
rect 528646 3856 528652 3868
rect 407080 3828 528652 3856
rect 407080 3816 407086 3828
rect 528646 3816 528652 3828
rect 528704 3816 528710 3868
rect 407393 3791 407451 3797
rect 407393 3788 407405 3791
rect 403820 3760 407405 3788
rect 407393 3757 407405 3760
rect 407439 3757 407451 3791
rect 407393 3751 407451 3757
rect 409506 3748 409512 3800
rect 409564 3788 409570 3800
rect 535730 3788 535736 3800
rect 409564 3760 535736 3788
rect 409564 3748 409570 3760
rect 535730 3748 535736 3760
rect 535788 3748 535794 3800
rect 333940 3692 340184 3720
rect 340233 3723 340291 3729
rect 333940 3680 333946 3692
rect 340233 3689 340245 3723
rect 340279 3720 340291 3723
rect 382366 3720 382372 3732
rect 340279 3692 382372 3720
rect 340279 3689 340291 3692
rect 340233 3683 340291 3689
rect 382366 3680 382372 3692
rect 382424 3680 382430 3732
rect 384298 3680 384304 3732
rect 384356 3720 384362 3732
rect 396626 3720 396632 3732
rect 384356 3692 396632 3720
rect 384356 3680 384362 3692
rect 396626 3680 396632 3692
rect 396684 3680 396690 3732
rect 396718 3680 396724 3732
rect 396776 3720 396782 3732
rect 410886 3720 410892 3732
rect 396776 3692 410892 3720
rect 396776 3680 396782 3692
rect 410886 3680 410892 3692
rect 410944 3680 410950 3732
rect 418154 3680 418160 3732
rect 418212 3720 418218 3732
rect 542906 3720 542912 3732
rect 418212 3692 542912 3720
rect 418212 3680 418218 3692
rect 542906 3680 542912 3692
rect 542964 3680 542970 3732
rect 14826 3612 14832 3664
rect 14884 3652 14890 3664
rect 140774 3652 140780 3664
rect 14884 3624 140780 3652
rect 14884 3612 14890 3624
rect 140774 3612 140780 3624
rect 140832 3612 140838 3664
rect 165890 3612 165896 3664
rect 165948 3652 165954 3664
rect 219618 3652 219624 3664
rect 165948 3624 219624 3652
rect 165948 3612 165954 3624
rect 219618 3612 219624 3624
rect 219676 3612 219682 3664
rect 224126 3612 224132 3664
rect 224184 3652 224190 3664
rect 228821 3655 228879 3661
rect 228821 3652 228833 3655
rect 224184 3624 228833 3652
rect 224184 3612 224190 3624
rect 228821 3621 228833 3624
rect 228867 3621 228879 3655
rect 228821 3615 228879 3621
rect 228910 3612 228916 3664
rect 228968 3652 228974 3664
rect 247678 3652 247684 3664
rect 228968 3624 247684 3652
rect 228968 3612 228974 3624
rect 247678 3612 247684 3624
rect 247736 3612 247742 3664
rect 284202 3612 284208 3664
rect 284260 3652 284266 3664
rect 289538 3652 289544 3664
rect 284260 3624 289544 3652
rect 284260 3612 284266 3624
rect 289538 3612 289544 3624
rect 289596 3612 289602 3664
rect 290918 3612 290924 3664
rect 290976 3652 290982 3664
rect 303798 3652 303804 3664
rect 290976 3624 303804 3652
rect 290976 3612 290982 3624
rect 303798 3612 303804 3624
rect 303856 3612 303862 3664
rect 306282 3612 306288 3664
rect 306340 3652 306346 3664
rect 332410 3652 332416 3664
rect 306340 3624 332416 3652
rect 306340 3612 306346 3624
rect 332410 3612 332416 3624
rect 332468 3612 332474 3664
rect 335262 3612 335268 3664
rect 335320 3652 335326 3664
rect 389450 3652 389456 3664
rect 335320 3624 389456 3652
rect 335320 3612 335326 3624
rect 389450 3612 389456 3624
rect 389508 3612 389514 3664
rect 393958 3612 393964 3664
rect 394016 3652 394022 3664
rect 398837 3655 398895 3661
rect 398837 3652 398849 3655
rect 394016 3624 398849 3652
rect 394016 3612 394022 3624
rect 398837 3621 398849 3624
rect 398883 3621 398895 3655
rect 398837 3615 398895 3621
rect 413186 3612 413192 3664
rect 413244 3652 413250 3664
rect 417973 3655 418031 3661
rect 417973 3652 417985 3655
rect 413244 3624 417985 3652
rect 413244 3612 413250 3624
rect 417973 3621 417985 3624
rect 418019 3621 418031 3655
rect 417973 3615 418031 3621
rect 420178 3612 420184 3664
rect 420236 3652 420242 3664
rect 553578 3652 553584 3664
rect 420236 3624 553584 3652
rect 420236 3612 420242 3624
rect 553578 3612 553584 3624
rect 553636 3612 553642 3664
rect 16022 3544 16028 3596
rect 16080 3584 16086 3596
rect 142338 3584 142344 3596
rect 16080 3556 142344 3584
rect 16080 3544 16086 3556
rect 142338 3544 142344 3556
rect 142396 3544 142402 3596
rect 162302 3544 162308 3596
rect 162360 3584 162366 3596
rect 216858 3584 216864 3596
rect 162360 3556 216864 3584
rect 162360 3544 162366 3556
rect 216858 3544 216864 3556
rect 216916 3544 216922 3596
rect 217873 3587 217931 3593
rect 217873 3553 217885 3587
rect 217919 3584 217931 3587
rect 223574 3584 223580 3596
rect 217919 3556 223580 3584
rect 217919 3553 217931 3556
rect 217873 3547 217931 3553
rect 223574 3544 223580 3556
rect 223632 3544 223638 3596
rect 234617 3587 234675 3593
rect 234617 3553 234629 3587
rect 234663 3584 234675 3587
rect 248598 3584 248604 3596
rect 234663 3556 248604 3584
rect 234663 3553 234675 3556
rect 234617 3547 234675 3553
rect 248598 3544 248604 3556
rect 248656 3544 248662 3596
rect 291102 3544 291108 3596
rect 291160 3584 291166 3596
rect 302602 3584 302608 3596
rect 291160 3556 302608 3584
rect 291160 3544 291166 3556
rect 302602 3544 302608 3556
rect 302660 3544 302666 3596
rect 303430 3544 303436 3596
rect 303488 3584 303494 3596
rect 328822 3584 328828 3596
rect 303488 3556 328828 3584
rect 303488 3544 303494 3556
rect 328822 3544 328828 3556
rect 328880 3544 328886 3596
rect 331122 3544 331128 3596
rect 331180 3584 331186 3596
rect 340233 3587 340291 3593
rect 340233 3584 340245 3587
rect 331180 3556 340245 3584
rect 331180 3544 331186 3556
rect 340233 3553 340245 3556
rect 340279 3553 340291 3587
rect 340233 3547 340291 3553
rect 341610 3544 341616 3596
rect 341668 3584 341674 3596
rect 343082 3584 343088 3596
rect 341668 3556 343088 3584
rect 341668 3544 341674 3556
rect 343082 3544 343088 3556
rect 343140 3544 343146 3596
rect 355229 3587 355287 3593
rect 355229 3553 355241 3587
rect 355275 3584 355287 3587
rect 366910 3584 366916 3596
rect 355275 3556 366916 3584
rect 355275 3553 355287 3556
rect 355229 3547 355287 3553
rect 366910 3544 366916 3556
rect 366968 3544 366974 3596
rect 398098 3544 398104 3596
rect 398156 3584 398162 3596
rect 408310 3584 408316 3596
rect 398156 3556 408316 3584
rect 398156 3544 398162 3556
rect 408310 3544 408316 3556
rect 408368 3544 408374 3596
rect 408494 3544 408500 3596
rect 408552 3584 408558 3596
rect 427630 3584 427636 3596
rect 408552 3556 427636 3584
rect 408552 3544 408558 3556
rect 427630 3544 427636 3556
rect 427688 3544 427694 3596
rect 427725 3587 427783 3593
rect 427725 3553 427737 3587
rect 427771 3584 427783 3587
rect 560754 3584 560760 3596
rect 427771 3556 560760 3584
rect 427771 3553 427783 3556
rect 427725 3547 427783 3553
rect 560754 3544 560760 3556
rect 560812 3544 560818 3596
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 138014 3516 138020 3528
rect 10100 3488 138020 3516
rect 10100 3476 10106 3488
rect 138014 3476 138020 3488
rect 138072 3476 138078 3528
rect 159910 3476 159916 3528
rect 159968 3516 159974 3528
rect 165614 3516 165620 3528
rect 159968 3488 165620 3516
rect 159968 3476 159974 3488
rect 165614 3476 165620 3488
rect 165672 3476 165678 3528
rect 175366 3476 175372 3528
rect 175424 3516 175430 3528
rect 177298 3516 177304 3528
rect 175424 3488 177304 3516
rect 175424 3476 175430 3488
rect 177298 3476 177304 3488
rect 177356 3476 177362 3528
rect 196802 3476 196808 3528
rect 196860 3516 196866 3528
rect 197262 3516 197268 3528
rect 196860 3488 197268 3516
rect 196860 3476 196866 3488
rect 197262 3476 197268 3488
rect 197320 3476 197326 3528
rect 200390 3476 200396 3528
rect 200448 3516 200454 3528
rect 201402 3516 201408 3528
rect 200448 3488 201408 3516
rect 200448 3476 200454 3488
rect 201402 3476 201408 3488
rect 201460 3476 201466 3528
rect 207474 3476 207480 3528
rect 207532 3516 207538 3528
rect 208302 3516 208308 3528
rect 207532 3488 208308 3516
rect 207532 3476 207538 3488
rect 208302 3476 208308 3488
rect 208360 3476 208366 3528
rect 209866 3476 209872 3528
rect 209924 3516 209930 3528
rect 211062 3516 211068 3528
rect 209924 3488 211068 3516
rect 209924 3476 209930 3488
rect 211062 3476 211068 3488
rect 211120 3476 211126 3528
rect 217229 3519 217287 3525
rect 217229 3485 217241 3519
rect 217275 3516 217287 3519
rect 229741 3519 229799 3525
rect 229741 3516 229753 3519
rect 217275 3488 229753 3516
rect 217275 3485 217287 3488
rect 217229 3479 217287 3485
rect 229741 3485 229753 3488
rect 229787 3485 229799 3519
rect 229741 3479 229799 3485
rect 257430 3476 257436 3528
rect 257488 3516 257494 3528
rect 257982 3516 257988 3528
rect 257488 3488 257988 3516
rect 257488 3476 257494 3488
rect 257982 3476 257988 3488
rect 258040 3476 258046 3528
rect 259822 3476 259828 3528
rect 259880 3516 259886 3528
rect 261478 3516 261484 3528
rect 259880 3488 261484 3516
rect 259880 3476 259886 3488
rect 261478 3476 261484 3488
rect 261536 3476 261542 3528
rect 262214 3476 262220 3528
rect 262272 3516 262278 3528
rect 263502 3516 263508 3528
rect 262272 3488 263508 3516
rect 262272 3476 262278 3488
rect 263502 3476 263508 3488
rect 263560 3476 263566 3528
rect 291010 3476 291016 3528
rect 291068 3516 291074 3528
rect 304994 3516 305000 3528
rect 291068 3488 305000 3516
rect 291068 3476 291074 3488
rect 304994 3476 305000 3488
rect 305052 3476 305058 3528
rect 305638 3476 305644 3528
rect 305696 3516 305702 3528
rect 306282 3516 306288 3528
rect 305696 3488 306288 3516
rect 305696 3476 305702 3488
rect 306282 3476 306288 3488
rect 306340 3476 306346 3528
rect 309042 3476 309048 3528
rect 309100 3516 309106 3528
rect 339494 3516 339500 3528
rect 309100 3488 339500 3516
rect 309100 3476 309106 3488
rect 339494 3476 339500 3488
rect 339552 3476 339558 3528
rect 344922 3476 344928 3528
rect 344980 3516 344986 3528
rect 407298 3516 407304 3528
rect 344980 3488 407304 3516
rect 344980 3476 344986 3488
rect 407298 3476 407304 3488
rect 407356 3476 407362 3528
rect 407393 3519 407451 3525
rect 407393 3485 407405 3519
rect 407439 3516 407451 3519
rect 417878 3516 417884 3528
rect 407439 3488 417884 3516
rect 407439 3485 407451 3488
rect 407393 3479 407451 3485
rect 417878 3476 417884 3488
rect 417936 3476 417942 3528
rect 417973 3519 418031 3525
rect 417973 3485 417985 3519
rect 418019 3516 418031 3519
rect 418157 3519 418215 3525
rect 418157 3516 418169 3519
rect 418019 3488 418169 3516
rect 418019 3485 418031 3488
rect 417973 3479 418031 3485
rect 418157 3485 418169 3488
rect 418203 3485 418215 3519
rect 421558 3516 421564 3528
rect 418157 3479 418215 3485
rect 418264 3488 421564 3516
rect 6454 3408 6460 3460
rect 6512 3448 6518 3460
rect 136910 3448 136916 3460
rect 6512 3420 136916 3448
rect 6512 3408 6518 3420
rect 136910 3408 136916 3420
rect 136968 3408 136974 3460
rect 144454 3408 144460 3460
rect 144512 3448 144518 3460
rect 208578 3448 208584 3460
rect 144512 3420 208584 3448
rect 144512 3408 144518 3420
rect 208578 3408 208584 3420
rect 208636 3408 208642 3460
rect 210053 3451 210111 3457
rect 210053 3417 210065 3451
rect 210099 3448 210111 3451
rect 214558 3448 214564 3460
rect 210099 3420 214564 3448
rect 210099 3417 210111 3420
rect 210053 3411 210111 3417
rect 214558 3408 214564 3420
rect 214616 3408 214622 3460
rect 217042 3408 217048 3460
rect 217100 3448 217106 3460
rect 243630 3448 243636 3460
rect 217100 3420 243636 3448
rect 217100 3408 217106 3420
rect 243630 3408 243636 3420
rect 243688 3408 243694 3460
rect 270494 3408 270500 3460
rect 270552 3448 270558 3460
rect 273346 3448 273352 3460
rect 270552 3420 273352 3448
rect 270552 3408 270558 3420
rect 273346 3408 273352 3420
rect 273404 3408 273410 3460
rect 285490 3408 285496 3460
rect 285548 3448 285554 3460
rect 294322 3448 294328 3460
rect 285548 3420 294328 3448
rect 285548 3408 285554 3420
rect 294322 3408 294328 3420
rect 294380 3408 294386 3460
rect 295242 3408 295248 3460
rect 295300 3448 295306 3460
rect 310974 3448 310980 3460
rect 295300 3420 310980 3448
rect 295300 3408 295306 3420
rect 310974 3408 310980 3420
rect 311032 3408 311038 3460
rect 313182 3408 313188 3460
rect 313240 3448 313246 3460
rect 346670 3448 346676 3460
rect 313240 3420 346676 3448
rect 313240 3408 313246 3420
rect 346670 3408 346676 3420
rect 346728 3408 346734 3460
rect 351822 3408 351828 3460
rect 351880 3448 351886 3460
rect 418264 3448 418292 3488
rect 421558 3476 421564 3488
rect 421616 3476 421622 3528
rect 427814 3476 427820 3528
rect 427872 3516 427878 3528
rect 439406 3516 439412 3528
rect 427872 3488 439412 3516
rect 427872 3476 427878 3488
rect 439406 3476 439412 3488
rect 439464 3476 439470 3528
rect 442261 3519 442319 3525
rect 442261 3485 442273 3519
rect 442307 3516 442319 3519
rect 567838 3516 567844 3528
rect 442307 3488 567844 3516
rect 442307 3485 442319 3488
rect 442261 3479 442319 3485
rect 567838 3476 567844 3488
rect 567896 3476 567902 3528
rect 351880 3420 418292 3448
rect 351880 3408 351886 3420
rect 418338 3408 418344 3460
rect 418396 3448 418402 3460
rect 432322 3448 432328 3460
rect 418396 3420 432328 3448
rect 418396 3408 418402 3420
rect 432322 3408 432328 3420
rect 432380 3408 432386 3460
rect 432509 3451 432567 3457
rect 432509 3417 432521 3451
rect 432555 3448 432567 3451
rect 437385 3451 437443 3457
rect 437385 3448 437397 3451
rect 432555 3420 437397 3448
rect 432555 3417 432567 3420
rect 432509 3411 432567 3417
rect 437385 3417 437397 3420
rect 437431 3417 437443 3451
rect 437385 3411 437443 3417
rect 442166 3408 442172 3460
rect 442224 3448 442230 3460
rect 582190 3448 582196 3460
rect 442224 3420 582196 3448
rect 442224 3408 442230 3420
rect 582190 3408 582196 3420
rect 582248 3408 582254 3460
rect 27890 3340 27896 3392
rect 27948 3380 27954 3392
rect 28902 3380 28908 3392
rect 27948 3352 28908 3380
rect 27948 3340 27954 3352
rect 28902 3340 28908 3352
rect 28960 3340 28966 3392
rect 50522 3340 50528 3392
rect 50580 3380 50586 3392
rect 158898 3380 158904 3392
rect 50580 3352 158904 3380
rect 50580 3340 50586 3352
rect 158898 3340 158904 3352
rect 158956 3340 158962 3392
rect 194410 3340 194416 3392
rect 194468 3380 194474 3392
rect 225233 3383 225291 3389
rect 225233 3380 225245 3383
rect 194468 3352 225245 3380
rect 194468 3340 194474 3352
rect 225233 3349 225245 3352
rect 225279 3349 225291 3383
rect 225233 3343 225291 3349
rect 225322 3340 225328 3392
rect 225380 3380 225386 3392
rect 226242 3380 226248 3392
rect 225380 3352 226248 3380
rect 225380 3340 225386 3352
rect 226242 3340 226248 3352
rect 226300 3340 226306 3392
rect 228821 3383 228879 3389
rect 228821 3349 228833 3383
rect 228867 3380 228879 3383
rect 234617 3383 234675 3389
rect 234617 3380 234629 3383
rect 228867 3352 234629 3380
rect 228867 3349 228879 3352
rect 228821 3343 228879 3349
rect 234617 3349 234629 3352
rect 234663 3349 234675 3383
rect 234617 3343 234675 3349
rect 250346 3340 250352 3392
rect 250404 3380 250410 3392
rect 251082 3380 251088 3392
rect 250404 3352 251088 3380
rect 250404 3340 250410 3352
rect 251082 3340 251088 3352
rect 251140 3340 251146 3392
rect 293862 3340 293868 3392
rect 293920 3380 293926 3392
rect 308582 3380 308588 3392
rect 293920 3352 308588 3380
rect 293920 3340 293926 3352
rect 308582 3340 308588 3352
rect 308640 3340 308646 3392
rect 320082 3340 320088 3392
rect 320140 3380 320146 3392
rect 359734 3380 359740 3392
rect 320140 3352 359740 3380
rect 320140 3340 320146 3352
rect 359734 3340 359740 3352
rect 359792 3340 359798 3392
rect 389082 3340 389088 3392
rect 389140 3380 389146 3392
rect 492950 3380 492956 3392
rect 389140 3352 492956 3380
rect 389140 3340 389146 3352
rect 492950 3340 492956 3352
rect 493008 3340 493014 3392
rect 496078 3340 496084 3392
rect 496136 3380 496142 3392
rect 504361 3383 504419 3389
rect 504361 3380 504373 3383
rect 496136 3352 504373 3380
rect 496136 3340 496142 3352
rect 504361 3349 504373 3352
rect 504407 3349 504419 3383
rect 564342 3380 564348 3392
rect 504361 3343 504419 3349
rect 504468 3352 564348 3380
rect 42150 3272 42156 3324
rect 42208 3312 42214 3324
rect 42702 3312 42708 3324
rect 42208 3284 42708 3312
rect 42208 3272 42214 3284
rect 42702 3272 42708 3284
rect 42760 3272 42766 3324
rect 45738 3272 45744 3324
rect 45796 3312 45802 3324
rect 143718 3312 143724 3324
rect 45796 3284 143724 3312
rect 45796 3272 45802 3284
rect 143718 3272 143724 3284
rect 143776 3272 143782 3324
rect 182542 3272 182548 3324
rect 182600 3312 182606 3324
rect 183462 3312 183468 3324
rect 182600 3284 183468 3312
rect 182600 3272 182606 3284
rect 183462 3272 183468 3284
rect 183520 3272 183526 3324
rect 193214 3272 193220 3324
rect 193272 3312 193278 3324
rect 194502 3312 194508 3324
rect 193272 3284 194508 3312
rect 193272 3272 193278 3284
rect 194502 3272 194508 3284
rect 194560 3272 194566 3324
rect 194597 3315 194655 3321
rect 194597 3281 194609 3315
rect 194643 3312 194655 3315
rect 232130 3312 232136 3324
rect 194643 3284 232136 3312
rect 194643 3281 194655 3284
rect 194597 3275 194655 3281
rect 232130 3272 232136 3284
rect 232188 3272 232194 3324
rect 244366 3272 244372 3324
rect 244424 3312 244430 3324
rect 245470 3312 245476 3324
rect 244424 3284 245476 3312
rect 244424 3272 244430 3284
rect 245470 3272 245476 3284
rect 245528 3272 245534 3324
rect 249150 3272 249156 3324
rect 249208 3312 249214 3324
rect 249702 3312 249708 3324
rect 249208 3284 249708 3312
rect 249208 3272 249214 3284
rect 249702 3272 249708 3284
rect 249760 3272 249766 3324
rect 253842 3272 253848 3324
rect 253900 3312 253906 3324
rect 257338 3312 257344 3324
rect 253900 3284 257344 3312
rect 253900 3272 253906 3284
rect 257338 3272 257344 3284
rect 257396 3272 257402 3324
rect 266998 3272 267004 3324
rect 267056 3312 267062 3324
rect 267642 3312 267648 3324
rect 267056 3284 267648 3312
rect 267056 3272 267062 3284
rect 267642 3272 267648 3284
rect 267700 3272 267706 3324
rect 292482 3272 292488 3324
rect 292540 3312 292546 3324
rect 306190 3312 306196 3324
rect 292540 3284 306196 3312
rect 292540 3272 292546 3284
rect 306190 3272 306196 3284
rect 306248 3272 306254 3324
rect 306282 3272 306288 3324
rect 306340 3312 306346 3324
rect 314562 3312 314568 3324
rect 306340 3284 314568 3312
rect 306340 3272 306346 3284
rect 314562 3272 314568 3284
rect 314620 3272 314626 3324
rect 317322 3272 317328 3324
rect 317380 3312 317386 3324
rect 353754 3312 353760 3324
rect 317380 3284 353760 3312
rect 317380 3272 317386 3284
rect 353754 3272 353760 3284
rect 353812 3272 353818 3324
rect 358170 3272 358176 3324
rect 358228 3312 358234 3324
rect 378778 3312 378784 3324
rect 358228 3284 378784 3312
rect 358228 3272 358234 3284
rect 378778 3272 378784 3284
rect 378836 3272 378842 3324
rect 383470 3272 383476 3324
rect 383528 3312 383534 3324
rect 482278 3312 482284 3324
rect 383528 3284 482284 3312
rect 383528 3272 383534 3284
rect 482278 3272 482284 3284
rect 482336 3272 482342 3324
rect 482373 3315 482431 3321
rect 482373 3281 482385 3315
rect 482419 3312 482431 3315
rect 485685 3315 485743 3321
rect 485685 3312 485697 3315
rect 482419 3284 485697 3312
rect 482419 3281 482431 3284
rect 482373 3275 482431 3281
rect 485685 3281 485697 3284
rect 485731 3281 485743 3315
rect 485685 3275 485743 3281
rect 486418 3272 486424 3324
rect 486476 3312 486482 3324
rect 489549 3315 489607 3321
rect 489549 3312 489561 3315
rect 486476 3284 489561 3312
rect 486476 3272 486482 3284
rect 489549 3281 489561 3284
rect 489595 3281 489607 3315
rect 489549 3275 489607 3281
rect 489641 3315 489699 3321
rect 489641 3281 489653 3315
rect 489687 3312 489699 3315
rect 489687 3284 493272 3312
rect 489687 3281 489699 3284
rect 489641 3275 489699 3281
rect 59998 3204 60004 3256
rect 60056 3244 60062 3256
rect 60642 3244 60648 3256
rect 60056 3216 60648 3244
rect 60056 3204 60062 3216
rect 60642 3204 60648 3216
rect 60700 3204 60706 3256
rect 73798 3204 73804 3256
rect 73856 3244 73862 3256
rect 74258 3244 74264 3256
rect 73856 3216 74264 3244
rect 73856 3204 73862 3216
rect 74258 3204 74264 3216
rect 74316 3204 74322 3256
rect 81434 3204 81440 3256
rect 81492 3244 81498 3256
rect 82722 3244 82728 3256
rect 81492 3216 82728 3244
rect 81492 3204 81498 3216
rect 82722 3204 82728 3216
rect 82780 3204 82786 3256
rect 89714 3204 89720 3256
rect 89772 3244 89778 3256
rect 179874 3244 179880 3256
rect 89772 3216 179880 3244
rect 89772 3204 89778 3216
rect 179874 3204 179880 3216
rect 179932 3204 179938 3256
rect 181346 3204 181352 3256
rect 181404 3244 181410 3256
rect 210053 3247 210111 3253
rect 210053 3244 210065 3247
rect 181404 3216 210065 3244
rect 181404 3204 181410 3216
rect 210053 3213 210065 3216
rect 210099 3213 210111 3247
rect 210053 3207 210111 3213
rect 211062 3204 211068 3256
rect 211120 3244 211126 3256
rect 217229 3247 217287 3253
rect 217229 3244 217241 3247
rect 211120 3216 217241 3244
rect 211120 3204 211126 3216
rect 217229 3213 217241 3216
rect 217275 3213 217287 3247
rect 217229 3207 217287 3213
rect 220538 3204 220544 3256
rect 220596 3244 220602 3256
rect 238018 3244 238024 3256
rect 220596 3216 238024 3244
rect 220596 3204 220602 3216
rect 238018 3204 238024 3216
rect 238076 3204 238082 3256
rect 246758 3204 246764 3256
rect 246816 3244 246822 3256
rect 250530 3244 250536 3256
rect 246816 3216 250536 3244
rect 246816 3204 246822 3216
rect 250530 3204 250536 3216
rect 250588 3204 250594 3256
rect 261018 3204 261024 3256
rect 261076 3244 261082 3256
rect 262122 3244 262128 3256
rect 261076 3216 262128 3244
rect 261076 3204 261082 3216
rect 262122 3204 262128 3216
rect 262180 3204 262186 3256
rect 281442 3204 281448 3256
rect 281500 3244 281506 3256
rect 285950 3244 285956 3256
rect 281500 3216 285956 3244
rect 281500 3204 281506 3216
rect 285950 3204 285956 3216
rect 286008 3204 286014 3256
rect 294598 3204 294604 3256
rect 294656 3244 294662 3256
rect 301406 3244 301412 3256
rect 294656 3216 301412 3244
rect 294656 3204 294662 3216
rect 301406 3204 301412 3216
rect 301464 3204 301470 3256
rect 315850 3204 315856 3256
rect 315908 3244 315914 3256
rect 321646 3244 321652 3256
rect 315908 3216 321652 3244
rect 315908 3204 315914 3216
rect 321646 3204 321652 3216
rect 321704 3204 321710 3256
rect 322198 3204 322204 3256
rect 322256 3244 322262 3256
rect 357342 3244 357348 3256
rect 322256 3216 357348 3244
rect 322256 3204 322262 3216
rect 357342 3204 357348 3216
rect 357400 3204 357406 3256
rect 379422 3204 379428 3256
rect 379480 3244 379486 3256
rect 475102 3244 475108 3256
rect 379480 3216 475108 3244
rect 379480 3204 379486 3216
rect 475102 3204 475108 3216
rect 475160 3204 475166 3256
rect 475378 3204 475384 3256
rect 475436 3244 475442 3256
rect 480901 3247 480959 3253
rect 480901 3244 480913 3247
rect 475436 3216 480913 3244
rect 475436 3204 475442 3216
rect 480901 3213 480913 3216
rect 480947 3213 480959 3247
rect 480901 3207 480959 3213
rect 480993 3247 481051 3253
rect 480993 3213 481005 3247
rect 481039 3244 481051 3247
rect 485133 3247 485191 3253
rect 485133 3244 485145 3247
rect 481039 3216 485145 3244
rect 481039 3213 481051 3216
rect 480993 3207 481051 3213
rect 485133 3213 485145 3216
rect 485179 3213 485191 3247
rect 493244 3244 493272 3284
rect 493318 3272 493324 3324
rect 493376 3312 493382 3324
rect 496633 3315 496691 3321
rect 496633 3312 496645 3315
rect 493376 3284 496645 3312
rect 493376 3272 493382 3284
rect 496633 3281 496645 3284
rect 496679 3281 496691 3315
rect 496633 3275 496691 3281
rect 502978 3272 502984 3324
rect 503036 3312 503042 3324
rect 504468 3312 504496 3352
rect 564342 3340 564348 3352
rect 564400 3340 564406 3392
rect 503036 3284 504496 3312
rect 504545 3315 504603 3321
rect 503036 3272 503042 3284
rect 504545 3281 504557 3315
rect 504591 3312 504603 3315
rect 557166 3312 557172 3324
rect 504591 3284 557172 3312
rect 504591 3281 504603 3284
rect 504545 3275 504603 3281
rect 557166 3272 557172 3284
rect 557224 3272 557230 3324
rect 503622 3244 503628 3256
rect 493244 3216 503628 3244
rect 485133 3207 485191 3213
rect 503622 3204 503628 3216
rect 503680 3204 503686 3256
rect 504361 3247 504419 3253
rect 504361 3213 504373 3247
rect 504407 3244 504419 3247
rect 550082 3244 550088 3256
rect 504407 3216 550088 3244
rect 504407 3213 504419 3216
rect 504361 3207 504419 3213
rect 550082 3204 550088 3216
rect 550140 3204 550146 3256
rect 55217 3179 55275 3185
rect 55217 3145 55229 3179
rect 55263 3176 55275 3179
rect 64785 3179 64843 3185
rect 64785 3176 64797 3179
rect 55263 3148 64797 3176
rect 55263 3145 55275 3148
rect 55217 3139 55275 3145
rect 64785 3145 64797 3148
rect 64831 3145 64843 3179
rect 64785 3139 64843 3145
rect 74537 3179 74595 3185
rect 74537 3145 74549 3179
rect 74583 3176 74595 3179
rect 84105 3179 84163 3185
rect 84105 3176 84117 3179
rect 74583 3148 84117 3176
rect 74583 3145 74595 3148
rect 74537 3139 74595 3145
rect 84105 3145 84117 3148
rect 84151 3145 84163 3179
rect 97258 3176 97264 3188
rect 84105 3139 84163 3145
rect 95528 3148 97264 3176
rect 92106 3068 92112 3120
rect 92164 3108 92170 3120
rect 95528 3108 95556 3148
rect 97258 3136 97264 3148
rect 97316 3136 97322 3188
rect 97994 3136 98000 3188
rect 98052 3176 98058 3188
rect 99282 3176 99288 3188
rect 98052 3148 99288 3176
rect 98052 3136 98058 3148
rect 99282 3136 99288 3148
rect 99340 3136 99346 3188
rect 183554 3176 183560 3188
rect 99392 3148 183560 3176
rect 92164 3080 95556 3108
rect 92164 3068 92170 3080
rect 96890 3068 96896 3120
rect 96948 3108 96954 3120
rect 99392 3108 99420 3148
rect 183554 3136 183560 3148
rect 183612 3136 183618 3188
rect 184842 3136 184848 3188
rect 184900 3176 184906 3188
rect 184900 3148 190132 3176
rect 184900 3136 184906 3148
rect 96948 3080 99420 3108
rect 96948 3068 96954 3080
rect 103974 3068 103980 3120
rect 104032 3108 104038 3120
rect 186590 3108 186596 3120
rect 104032 3080 186596 3108
rect 104032 3068 104038 3080
rect 186590 3068 186596 3080
rect 186648 3068 186654 3120
rect 190104 3108 190132 3148
rect 192018 3136 192024 3188
rect 192076 3176 192082 3188
rect 194597 3179 194655 3185
rect 194597 3176 194609 3179
rect 192076 3148 194609 3176
rect 192076 3136 192082 3148
rect 194597 3145 194609 3148
rect 194643 3145 194655 3179
rect 194597 3139 194655 3145
rect 203886 3136 203892 3188
rect 203944 3176 203950 3188
rect 233878 3176 233884 3188
rect 203944 3148 233884 3176
rect 203944 3136 203950 3148
rect 233878 3136 233884 3148
rect 233936 3136 233942 3188
rect 281350 3136 281356 3188
rect 281408 3176 281414 3188
rect 284754 3176 284760 3188
rect 281408 3148 284760 3176
rect 281408 3136 281414 3148
rect 284754 3136 284760 3148
rect 284812 3136 284818 3188
rect 297358 3136 297364 3188
rect 297416 3176 297422 3188
rect 300302 3176 300308 3188
rect 297416 3148 300308 3176
rect 297416 3136 297422 3148
rect 300302 3136 300308 3148
rect 300360 3136 300366 3188
rect 302878 3136 302884 3188
rect 302936 3176 302942 3188
rect 309778 3176 309784 3188
rect 302936 3148 309784 3176
rect 302936 3136 302942 3148
rect 309778 3136 309784 3148
rect 309836 3136 309842 3188
rect 320818 3136 320824 3188
rect 320876 3176 320882 3188
rect 350258 3176 350264 3188
rect 320876 3148 350264 3176
rect 320876 3136 320882 3148
rect 350258 3136 350264 3148
rect 350316 3136 350322 3188
rect 375282 3136 375288 3188
rect 375340 3176 375346 3188
rect 467926 3176 467932 3188
rect 375340 3148 467932 3176
rect 375340 3136 375346 3148
rect 467926 3136 467932 3148
rect 467984 3136 467990 3188
rect 473998 3136 474004 3188
rect 474056 3176 474062 3188
rect 496538 3176 496544 3188
rect 474056 3148 496544 3176
rect 474056 3136 474062 3148
rect 496538 3136 496544 3148
rect 496596 3136 496602 3188
rect 496633 3179 496691 3185
rect 496633 3145 496645 3179
rect 496679 3176 496691 3179
rect 546494 3176 546500 3188
rect 496679 3148 546500 3176
rect 496679 3145 496691 3148
rect 496633 3139 496691 3145
rect 546494 3136 546500 3148
rect 546552 3136 546558 3188
rect 193858 3108 193864 3120
rect 190104 3080 193864 3108
rect 193858 3068 193864 3080
rect 193916 3068 193922 3120
rect 202690 3068 202696 3120
rect 202748 3108 202754 3120
rect 231118 3108 231124 3120
rect 202748 3080 231124 3108
rect 202748 3068 202754 3080
rect 231118 3068 231124 3080
rect 231176 3068 231182 3120
rect 258626 3068 258632 3120
rect 258684 3108 258690 3120
rect 259362 3108 259368 3120
rect 258684 3080 259368 3108
rect 258684 3068 258690 3080
rect 259362 3068 259368 3080
rect 259420 3068 259426 3120
rect 264606 3068 264612 3120
rect 264664 3108 264670 3120
rect 268378 3108 268384 3120
rect 264664 3080 268384 3108
rect 264664 3068 264670 3080
rect 268378 3068 268384 3080
rect 268436 3068 268442 3120
rect 372522 3068 372528 3120
rect 372580 3108 372586 3120
rect 460842 3108 460848 3120
rect 372580 3080 460848 3108
rect 372580 3068 372586 3080
rect 460842 3068 460848 3080
rect 460900 3068 460906 3120
rect 469858 3068 469864 3120
rect 469916 3108 469922 3120
rect 489362 3108 489368 3120
rect 469916 3080 489368 3108
rect 469916 3068 469922 3080
rect 489362 3068 489368 3080
rect 489420 3068 489426 3120
rect 539318 3108 539324 3120
rect 489472 3080 539324 3108
rect 111150 3000 111156 3052
rect 111208 3040 111214 3052
rect 190730 3040 190736 3052
rect 111208 3012 190736 3040
rect 111208 3000 111214 3012
rect 190730 3000 190736 3012
rect 190788 3000 190794 3052
rect 199194 3000 199200 3052
rect 199252 3040 199258 3052
rect 225598 3040 225604 3052
rect 199252 3012 225604 3040
rect 199252 3000 199258 3012
rect 225598 3000 225604 3012
rect 225656 3000 225662 3052
rect 252646 3000 252652 3052
rect 252704 3040 252710 3052
rect 254578 3040 254584 3052
rect 252704 3012 254584 3040
rect 252704 3000 252710 3012
rect 254578 3000 254584 3012
rect 254636 3000 254642 3052
rect 377398 3000 377404 3052
rect 377456 3040 377462 3052
rect 453666 3040 453672 3052
rect 377456 3012 453672 3040
rect 377456 3000 377462 3012
rect 453666 3000 453672 3012
rect 453724 3000 453730 3052
rect 463697 3043 463755 3049
rect 463697 3009 463709 3043
rect 463743 3040 463755 3043
rect 473265 3043 473323 3049
rect 473265 3040 473277 3043
rect 463743 3012 473277 3040
rect 463743 3009 463755 3012
rect 463697 3003 463755 3009
rect 473265 3009 473277 3012
rect 473311 3009 473323 3043
rect 473265 3003 473323 3009
rect 480901 3043 480959 3049
rect 480901 3009 480913 3043
rect 480947 3040 480959 3043
rect 489089 3043 489147 3049
rect 489089 3040 489101 3043
rect 480947 3012 489101 3040
rect 480947 3009 480959 3012
rect 480901 3003 480959 3009
rect 489089 3009 489101 3012
rect 489135 3009 489147 3043
rect 489089 3003 489147 3009
rect 489178 3000 489184 3052
rect 489236 3040 489242 3052
rect 489472 3040 489500 3080
rect 539318 3068 539324 3080
rect 539376 3068 539382 3120
rect 489236 3012 489500 3040
rect 489549 3043 489607 3049
rect 489236 3000 489242 3012
rect 489549 3009 489561 3043
rect 489595 3040 489607 3043
rect 532234 3040 532240 3052
rect 489595 3012 532240 3040
rect 489595 3009 489607 3012
rect 489549 3003 489607 3009
rect 532234 3000 532240 3012
rect 532292 3000 532298 3052
rect 93857 2975 93915 2981
rect 93857 2941 93869 2975
rect 93903 2972 93915 2975
rect 103425 2975 103483 2981
rect 103425 2972 103437 2975
rect 93903 2944 103437 2972
rect 93903 2941 93915 2944
rect 93857 2935 93915 2941
rect 103425 2941 103437 2944
rect 103471 2941 103483 2975
rect 103425 2935 103483 2941
rect 118234 2932 118240 2984
rect 118292 2972 118298 2984
rect 194778 2972 194784 2984
rect 118292 2944 194784 2972
rect 118292 2932 118298 2944
rect 194778 2932 194784 2944
rect 194836 2932 194842 2984
rect 197998 2932 198004 2984
rect 198056 2972 198062 2984
rect 204162 2972 204168 2984
rect 198056 2944 204168 2972
rect 198056 2932 198062 2944
rect 204162 2932 204168 2944
rect 204220 2932 204226 2984
rect 206278 2932 206284 2984
rect 206336 2972 206342 2984
rect 232406 2972 232412 2984
rect 206336 2944 232412 2972
rect 206336 2932 206342 2944
rect 232406 2932 232412 2944
rect 232464 2932 232470 2984
rect 308398 2932 308404 2984
rect 308456 2972 308462 2984
rect 313366 2972 313372 2984
rect 308456 2944 313372 2972
rect 308456 2932 308462 2944
rect 313366 2932 313372 2944
rect 313424 2932 313430 2984
rect 369118 2932 369124 2984
rect 369176 2972 369182 2984
rect 371602 2972 371608 2984
rect 369176 2944 371608 2972
rect 369176 2932 369182 2944
rect 371602 2932 371608 2944
rect 371660 2932 371666 2984
rect 376018 2932 376024 2984
rect 376076 2972 376082 2984
rect 414474 2972 414480 2984
rect 376076 2944 414480 2972
rect 376076 2932 376082 2944
rect 414474 2932 414480 2944
rect 414532 2932 414538 2984
rect 416038 2932 416044 2984
rect 416096 2972 416102 2984
rect 418154 2972 418160 2984
rect 416096 2944 418160 2972
rect 416096 2932 416102 2944
rect 418154 2932 418160 2944
rect 418212 2932 418218 2984
rect 418249 2975 418307 2981
rect 418249 2941 418261 2975
rect 418295 2972 418307 2975
rect 422297 2975 422355 2981
rect 422297 2972 422309 2975
rect 418295 2944 422309 2972
rect 418295 2941 418307 2944
rect 418249 2935 418307 2941
rect 422297 2941 422309 2944
rect 422343 2941 422355 2975
rect 422297 2935 422355 2941
rect 424318 2932 424324 2984
rect 424376 2972 424382 2984
rect 427725 2975 427783 2981
rect 427725 2972 427737 2975
rect 424376 2944 427737 2972
rect 424376 2932 424382 2944
rect 427725 2941 427737 2944
rect 427771 2941 427783 2975
rect 427725 2935 427783 2941
rect 437385 2975 437443 2981
rect 437385 2941 437397 2975
rect 437431 2972 437443 2975
rect 437431 2944 456840 2972
rect 437431 2941 437443 2944
rect 437385 2935 437443 2941
rect 113177 2907 113235 2913
rect 113177 2873 113189 2907
rect 113223 2904 113235 2907
rect 123481 2907 123539 2913
rect 123481 2904 123493 2907
rect 113223 2876 123493 2904
rect 113223 2873 113235 2876
rect 113177 2867 113235 2873
rect 123481 2873 123493 2876
rect 123527 2873 123539 2907
rect 123481 2867 123539 2873
rect 133141 2907 133199 2913
rect 133141 2873 133153 2907
rect 133187 2904 133199 2907
rect 142801 2907 142859 2913
rect 142801 2904 142813 2907
rect 133187 2876 142813 2904
rect 133187 2873 133199 2876
rect 133141 2867 133199 2873
rect 142801 2873 142813 2876
rect 142847 2873 142859 2907
rect 142801 2867 142859 2873
rect 201494 2864 201500 2916
rect 201552 2904 201558 2916
rect 203794 2904 203800 2916
rect 201552 2876 203800 2904
rect 201552 2864 201558 2876
rect 203794 2864 203800 2876
rect 203852 2864 203858 2916
rect 214650 2864 214656 2916
rect 214708 2904 214714 2916
rect 239398 2904 239404 2916
rect 214708 2876 239404 2904
rect 214708 2864 214714 2876
rect 239398 2864 239404 2876
rect 239456 2864 239462 2916
rect 369394 2864 369400 2916
rect 369452 2904 369458 2916
rect 428734 2904 428740 2916
rect 369452 2876 428740 2904
rect 369452 2864 369458 2876
rect 428734 2864 428740 2876
rect 428792 2864 428798 2916
rect 429838 2864 429844 2916
rect 429896 2904 429902 2916
rect 442261 2907 442319 2913
rect 442261 2904 442273 2907
rect 429896 2876 442273 2904
rect 429896 2864 429902 2876
rect 442261 2873 442273 2876
rect 442307 2873 442319 2907
rect 456812 2904 456840 2944
rect 478138 2932 478144 2984
rect 478196 2972 478202 2984
rect 480993 2975 481051 2981
rect 480993 2972 481005 2975
rect 478196 2944 481005 2972
rect 478196 2932 478202 2944
rect 480993 2941 481005 2944
rect 481039 2941 481051 2975
rect 480993 2935 481051 2941
rect 481085 2975 481143 2981
rect 481085 2941 481097 2975
rect 481131 2972 481143 2975
rect 482097 2975 482155 2981
rect 482097 2972 482109 2975
rect 481131 2944 482109 2972
rect 481131 2941 481143 2944
rect 481085 2935 481143 2941
rect 482097 2941 482109 2944
rect 482143 2941 482155 2975
rect 482097 2935 482155 2941
rect 482186 2932 482192 2984
rect 482244 2972 482250 2984
rect 485041 2975 485099 2981
rect 485041 2972 485053 2975
rect 482244 2944 485053 2972
rect 482244 2932 482250 2944
rect 485041 2941 485053 2944
rect 485087 2941 485099 2975
rect 485041 2935 485099 2941
rect 485133 2975 485191 2981
rect 485133 2941 485145 2975
rect 485179 2972 485191 2975
rect 510798 2972 510804 2984
rect 485179 2944 510804 2972
rect 485179 2941 485191 2944
rect 485133 2935 485191 2941
rect 510798 2932 510804 2944
rect 510856 2932 510862 2984
rect 463697 2907 463755 2913
rect 463697 2904 463709 2907
rect 456812 2876 463709 2904
rect 442261 2867 442319 2873
rect 463697 2873 463709 2876
rect 463743 2873 463755 2907
rect 463697 2867 463755 2873
rect 485685 2907 485743 2913
rect 485685 2873 485697 2907
rect 485731 2904 485743 2907
rect 485774 2904 485780 2916
rect 485731 2876 485780 2904
rect 485731 2873 485743 2876
rect 485685 2867 485743 2873
rect 485774 2864 485780 2876
rect 485832 2864 485838 2916
rect 525058 2904 525064 2916
rect 485884 2876 525064 2904
rect 148042 2796 148048 2848
rect 148100 2836 148106 2848
rect 209958 2836 209964 2848
rect 148100 2808 209964 2836
rect 148100 2796 148106 2808
rect 209958 2796 209964 2808
rect 210016 2796 210022 2848
rect 340782 2796 340788 2848
rect 340840 2836 340846 2848
rect 400214 2836 400220 2848
rect 340840 2808 400220 2836
rect 340840 2796 340846 2808
rect 400214 2796 400220 2808
rect 400272 2796 400278 2848
rect 402238 2796 402244 2848
rect 402296 2836 402302 2848
rect 446582 2836 446588 2848
rect 402296 2808 446588 2836
rect 402296 2796 402302 2808
rect 446582 2796 446588 2808
rect 446640 2796 446646 2848
rect 473265 2839 473323 2845
rect 473265 2805 473277 2839
rect 473311 2836 473323 2839
rect 480809 2839 480867 2845
rect 480809 2836 480821 2839
rect 473311 2808 480821 2836
rect 473311 2805 473323 2808
rect 473265 2799 473323 2805
rect 480809 2805 480821 2808
rect 480855 2805 480867 2839
rect 480809 2799 480867 2805
rect 480898 2796 480904 2848
rect 480956 2836 480962 2848
rect 483017 2839 483075 2845
rect 483017 2836 483029 2839
rect 480956 2808 483029 2836
rect 480956 2796 480962 2808
rect 483017 2805 483029 2808
rect 483063 2805 483075 2839
rect 483017 2799 483075 2805
rect 485041 2839 485099 2845
rect 485041 2805 485053 2839
rect 485087 2836 485099 2839
rect 485884 2836 485912 2876
rect 525058 2864 525064 2876
rect 525116 2864 525122 2916
rect 517882 2836 517888 2848
rect 485087 2808 485912 2836
rect 485976 2808 517888 2836
rect 485087 2805 485099 2808
rect 485041 2799 485099 2805
rect 422297 2771 422355 2777
rect 422297 2737 422309 2771
rect 422343 2768 422355 2771
rect 432509 2771 432567 2777
rect 432509 2768 432521 2771
rect 422343 2740 432521 2768
rect 422343 2737 422355 2740
rect 422297 2731 422355 2737
rect 432509 2737 432521 2740
rect 432555 2737 432567 2771
rect 432509 2731 432567 2737
rect 483017 2703 483075 2709
rect 483017 2669 483029 2703
rect 483063 2700 483075 2703
rect 485976 2700 486004 2808
rect 517882 2796 517888 2808
rect 517940 2796 517946 2848
rect 483063 2672 486004 2700
rect 483063 2669 483075 2672
rect 483017 2663 483075 2669
rect 23106 552 23112 604
rect 23164 592 23170 604
rect 23382 592 23388 604
rect 23164 564 23388 592
rect 23164 552 23170 564
rect 23382 552 23388 564
rect 23440 552 23446 604
rect 178954 552 178960 604
rect 179012 592 179018 604
rect 179322 592 179328 604
rect 179012 564 179328 592
rect 179012 552 179018 564
rect 179322 552 179328 564
rect 179380 552 179386 604
rect 272886 552 272892 604
rect 272944 592 272950 604
rect 273162 592 273168 604
rect 272944 564 273168 592
rect 272944 552 272950 564
rect 273162 552 273168 564
rect 273220 552 273226 604
rect 290090 552 290096 604
rect 290148 592 290154 604
rect 290734 592 290740 604
rect 290148 564 290740 592
rect 290148 552 290154 564
rect 290734 552 290740 564
rect 290792 552 290798 604
rect 291378 552 291384 604
rect 291436 592 291442 604
rect 291930 592 291936 604
rect 291436 564 291936 592
rect 291436 552 291442 564
rect 291930 552 291936 564
rect 291988 552 291994 604
rect 318978 552 318984 604
rect 319036 592 319042 604
rect 319254 592 319260 604
rect 319036 564 319260 592
rect 319036 552 319042 564
rect 319254 552 319260 564
rect 319312 552 319318 604
rect 326430 592 326436 604
rect 326391 564 326436 592
rect 326430 552 326436 564
rect 326488 552 326494 604
rect 332870 552 332876 604
rect 332928 592 332934 604
rect 333606 592 333612 604
rect 332928 564 333612 592
rect 332928 552 332934 564
rect 333606 552 333612 564
rect 333664 552 333670 604
rect 336918 552 336924 604
rect 336976 592 336982 604
rect 337102 592 337108 604
rect 336976 564 337108 592
rect 336976 552 336982 564
rect 337102 552 337108 564
rect 337160 552 337166 604
rect 343910 552 343916 604
rect 343968 592 343974 604
rect 344278 592 344284 604
rect 343968 564 344284 592
rect 343968 552 343974 564
rect 344278 552 344284 564
rect 344336 552 344342 604
rect 425146 552 425152 604
rect 425204 592 425210 604
rect 425330 592 425336 604
rect 425204 564 425336 592
rect 425204 552 425210 564
rect 425330 552 425336 564
rect 425388 552 425394 604
rect 456794 552 456800 604
rect 456852 592 456858 604
rect 457254 592 457260 604
rect 456852 564 457260 592
rect 456852 552 456858 564
rect 457254 552 457260 564
rect 457312 552 457318 604
rect 470594 552 470600 604
rect 470652 592 470658 604
rect 471514 592 471520 604
rect 470652 564 471520 592
rect 470652 552 470658 564
rect 471514 552 471520 564
rect 471572 552 471578 604
rect 473354 552 473360 604
rect 473412 592 473418 604
rect 473906 592 473912 604
rect 473412 564 473912 592
rect 473412 552 473418 564
rect 473906 552 473912 564
rect 473964 552 473970 604
<< via1 >>
rect 133972 700952 134024 701004
rect 267648 700952 267700 701004
rect 133788 700884 133840 700936
rect 283840 700884 283892 700936
rect 300124 700884 300176 700936
rect 434076 700884 434128 700936
rect 132500 700816 132552 700868
rect 332508 700816 332560 700868
rect 133696 700748 133748 700800
rect 218980 700748 219032 700800
rect 235172 700748 235224 700800
rect 434168 700748 434220 700800
rect 131120 700680 131172 700732
rect 348792 700680 348844 700732
rect 364984 700680 365036 700732
rect 433984 700680 434036 700732
rect 170312 700612 170364 700664
rect 434352 700612 434404 700664
rect 131212 700544 131264 700596
rect 397460 700544 397512 700596
rect 132316 700476 132368 700528
rect 413652 700476 413704 700528
rect 105452 700408 105504 700460
rect 434444 700408 434496 700460
rect 438124 700408 438176 700460
rect 494796 700408 494848 700460
rect 8116 700340 8168 700392
rect 13084 700340 13136 700392
rect 89168 700340 89220 700392
rect 126244 700340 126296 700392
rect 132592 700340 132644 700392
rect 462320 700340 462372 700392
rect 40500 700272 40552 700324
rect 434260 700272 434312 700324
rect 447784 700272 447836 700324
rect 559656 700272 559708 700324
rect 133420 700204 133472 700256
rect 202788 700204 202840 700256
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 72424 699660 72476 699712
rect 72976 699660 73028 699712
rect 133328 699660 133380 699712
rect 137836 699660 137888 699712
rect 429844 699660 429896 699712
rect 433892 699660 433944 699712
rect 153568 698232 153620 698284
rect 154212 698232 154264 698284
rect 147588 697076 147640 697128
rect 154488 697076 154540 697128
rect 166908 697076 166960 697128
rect 173808 697076 173860 697128
rect 186228 697076 186280 697128
rect 193128 697076 193180 697128
rect 205548 697076 205600 697128
rect 212448 697076 212500 697128
rect 224868 697076 224920 697128
rect 231768 697076 231820 697128
rect 244188 697076 244240 697128
rect 251088 697076 251140 697128
rect 263508 697076 263560 697128
rect 270408 697076 270460 697128
rect 282828 697076 282880 697128
rect 289728 697076 289780 697128
rect 302148 697076 302200 697128
rect 309048 697076 309100 697128
rect 321468 697076 321520 697128
rect 328368 697076 328420 697128
rect 154580 686264 154632 686316
rect 159456 686264 159508 686316
rect 135260 686128 135312 686180
rect 142896 686128 142948 686180
rect 153292 685924 153344 685976
rect 153660 685924 153712 685976
rect 153292 684428 153344 684480
rect 3516 681708 3568 681760
rect 434720 681708 434772 681760
rect 446404 673480 446456 673532
rect 580172 673480 580224 673532
rect 3424 667904 3476 667956
rect 19984 667904 20036 667956
rect 153660 666544 153712 666596
rect 153476 656863 153528 656872
rect 153476 656829 153485 656863
rect 153485 656829 153519 656863
rect 153519 656829 153528 656863
rect 153476 656820 153528 656829
rect 154580 650360 154632 650412
rect 159456 650360 159508 650412
rect 135260 650224 135312 650276
rect 142896 650224 142948 650276
rect 153568 647232 153620 647284
rect 153292 637644 153344 637696
rect 153568 637644 153620 637696
rect 153384 630708 153436 630760
rect 153568 630504 153620 630556
rect 445024 626560 445076 626612
rect 580172 626560 580224 626612
rect 153568 626492 153620 626544
rect 153752 626492 153804 626544
rect 3424 623772 3476 623824
rect 434812 623772 434864 623824
rect 153568 611192 153620 611244
rect 153752 611192 153804 611244
rect 3424 609968 3476 610020
rect 21364 609968 21416 610020
rect 153384 598952 153436 599004
rect 153568 598952 153620 599004
rect 4068 594804 4120 594856
rect 4896 594804 4948 594856
rect 153292 591948 153344 592000
rect 153568 591948 153620 592000
rect 175924 583652 175976 583704
rect 302792 583652 302844 583704
rect 270408 583584 270460 583636
rect 307024 583584 307076 583636
rect 286324 583516 286376 583568
rect 319720 583516 319772 583568
rect 129280 583448 129332 583500
rect 347504 583448 347556 583500
rect 126336 583380 126388 583432
rect 324136 583380 324188 583432
rect 85396 583312 85448 583364
rect 334624 583312 334676 583364
rect 85580 583244 85632 583296
rect 345296 583244 345348 583296
rect 291844 583176 291896 583228
rect 328368 583176 328420 583228
rect 298928 583108 298980 583160
rect 341064 583108 341116 583160
rect 294604 583040 294656 583092
rect 338856 583040 338908 583092
rect 281356 582972 281408 583024
rect 326160 582972 326212 583024
rect 299020 582904 299072 582956
rect 353760 582904 353812 582956
rect 298652 582836 298704 582888
rect 355968 582836 356020 582888
rect 291108 582768 291160 582820
rect 351736 582768 351788 582820
rect 298744 582700 298796 582752
rect 360200 582700 360252 582752
rect 300492 582632 300544 582684
rect 362408 582632 362460 582684
rect 366640 582632 366692 582684
rect 378876 582632 378928 582684
rect 298836 582564 298888 582616
rect 332600 582564 332652 582616
rect 357992 582564 358044 582616
rect 378416 582564 378468 582616
rect 298468 582496 298520 582548
rect 321928 582496 321980 582548
rect 370872 582496 370924 582548
rect 378692 582496 378744 582548
rect 287704 582428 287756 582480
rect 313464 582428 313516 582480
rect 298560 582360 298612 582412
rect 309232 582360 309284 582412
rect 372896 582360 372948 582412
rect 378600 582360 378652 582412
rect 299388 579640 299440 579692
rect 304816 579640 304868 579692
rect 442264 579640 442316 579692
rect 580172 579640 580224 579692
rect 153384 579615 153436 579624
rect 153384 579581 153393 579615
rect 153393 579581 153427 579615
rect 153427 579581 153436 579615
rect 153384 579572 153436 579581
rect 299480 579300 299532 579352
rect 300676 579300 300728 579352
rect 310980 579343 311032 579352
rect 310980 579309 310989 579343
rect 310989 579309 311023 579343
rect 311023 579309 311032 579343
rect 310980 579300 311032 579309
rect 315212 579343 315264 579352
rect 315212 579309 315221 579343
rect 315221 579309 315255 579343
rect 315255 579309 315264 579343
rect 315212 579300 315264 579309
rect 317420 579343 317472 579352
rect 317420 579309 317429 579343
rect 317429 579309 317463 579343
rect 317463 579309 317472 579343
rect 317420 579300 317472 579309
rect 330208 579300 330260 579352
rect 336648 579343 336700 579352
rect 336648 579309 336657 579343
rect 336657 579309 336691 579343
rect 336691 579309 336700 579343
rect 336648 579300 336700 579309
rect 342996 579343 343048 579352
rect 342996 579309 343005 579343
rect 343005 579309 343039 579343
rect 343039 579309 343048 579343
rect 342996 579300 343048 579309
rect 364248 579343 364300 579352
rect 364248 579309 364257 579343
rect 364257 579309 364291 579343
rect 364291 579309 364300 579343
rect 364248 579300 364300 579309
rect 375380 579300 375432 579352
rect 378508 579300 378560 579352
rect 129004 578756 129056 578808
rect 130384 578688 130436 578740
rect 122748 578552 122800 578604
rect 115388 578416 115440 578468
rect 119344 578348 119396 578400
rect 115204 578280 115256 578332
rect 129188 578212 129240 578264
rect 110328 575492 110380 575544
rect 296720 575492 296772 575544
rect 153476 569916 153528 569968
rect 272524 569916 272576 569968
rect 298008 569916 298060 569968
rect 153476 563116 153528 563168
rect 129556 563048 129608 563100
rect 296904 563048 296956 563100
rect 153292 563023 153344 563032
rect 153292 562989 153301 563023
rect 153301 562989 153335 563023
rect 153335 562989 153344 563023
rect 153292 562980 153344 562989
rect 195888 561960 195940 562012
rect 197084 561892 197136 561944
rect 208676 561892 208728 561944
rect 217876 561892 217928 561944
rect 196992 561824 197044 561876
rect 205548 561824 205600 561876
rect 197268 561756 197320 561808
rect 214748 561756 214800 561808
rect 153292 560235 153344 560244
rect 153292 560201 153301 560235
rect 153301 560201 153335 560235
rect 153335 560201 153344 560235
rect 153292 560192 153344 560201
rect 197176 560192 197228 560244
rect 202052 560192 202104 560244
rect 420184 556248 420236 556300
rect 511264 556248 511316 556300
rect 273168 556180 273220 556232
rect 297088 556180 297140 556232
rect 378784 556180 378836 556232
rect 484400 556180 484452 556232
rect 109408 554752 109460 554804
rect 110328 554752 110380 554804
rect 115940 554752 115992 554804
rect 92112 553936 92164 553988
rect 115296 553936 115348 553988
rect 89168 553868 89220 553920
rect 162124 553868 162176 553920
rect 115112 553800 115164 553852
rect 128360 553800 128412 553852
rect 129280 553800 129332 553852
rect 95056 553732 95108 553784
rect 120724 553732 120776 553784
rect 100760 553664 100812 553716
rect 129096 553664 129148 553716
rect 106464 553596 106516 553648
rect 140044 553596 140096 553648
rect 103704 553528 103756 553580
rect 151084 553528 151136 553580
rect 97816 553460 97868 553512
rect 157984 553460 158036 553512
rect 112352 553392 112404 553444
rect 116032 553392 116084 553444
rect 3148 552032 3200 552084
rect 28264 552032 28316 552084
rect 153476 550604 153528 550656
rect 85488 549856 85540 549908
rect 86408 549856 86460 549908
rect 115388 549856 115440 549908
rect 153292 543600 153344 543652
rect 153476 543600 153528 543652
rect 286876 538228 286928 538280
rect 297732 538228 297784 538280
rect 117320 536800 117372 536852
rect 146944 536800 146996 536852
rect 118240 534012 118292 534064
rect 118516 534012 118568 534064
rect 153292 534012 153344 534064
rect 153476 534012 153528 534064
rect 295984 532856 296036 532908
rect 297456 532856 297508 532908
rect 117320 532720 117372 532772
rect 160744 532720 160796 532772
rect 514024 532720 514076 532772
rect 580172 532720 580224 532772
rect 117964 529864 118016 529916
rect 119344 529864 119396 529916
rect 117320 525036 117372 525088
rect 129188 525036 129240 525088
rect 70308 524424 70360 524476
rect 82820 524424 82872 524476
rect 118516 524492 118568 524544
rect 118424 524356 118476 524408
rect 128912 521636 128964 521688
rect 129188 521636 129240 521688
rect 153568 521636 153620 521688
rect 153752 521636 153804 521688
rect 280068 521636 280120 521688
rect 297088 521636 297140 521688
rect 295340 521568 295392 521620
rect 295984 521568 296036 521620
rect 85304 521228 85356 521280
rect 295340 521228 295392 521280
rect 199384 521092 199436 521144
rect 222384 521092 222436 521144
rect 199476 521024 199528 521076
rect 222568 521024 222620 521076
rect 198280 520956 198332 521008
rect 222660 520956 222712 521008
rect 117320 520888 117372 520940
rect 128452 520888 128504 520940
rect 129004 520888 129056 520940
rect 198188 520888 198240 520940
rect 222476 520888 222528 520940
rect 86592 518712 86644 518764
rect 122748 518916 122800 518968
rect 279424 518916 279476 518968
rect 297732 518916 297784 518968
rect 89352 518848 89404 518900
rect 129832 518848 129884 518900
rect 130384 518848 130436 518900
rect 109592 518780 109644 518832
rect 113824 518780 113876 518832
rect 115204 518780 115256 518832
rect 127716 518780 127768 518832
rect 98000 518372 98052 518424
rect 144184 518372 144236 518424
rect 106648 518304 106700 518356
rect 153844 518304 153896 518356
rect 100944 518236 100996 518288
rect 159364 518236 159416 518288
rect 198096 518236 198148 518288
rect 218980 518236 219032 518288
rect 92296 518168 92348 518220
rect 126980 518168 127032 518220
rect 297456 518168 297508 518220
rect 205640 517488 205692 517540
rect 206652 517488 206704 517540
rect 284944 516128 284996 516180
rect 297732 516128 297784 516180
rect 118240 511980 118292 512032
rect 118516 511980 118568 512032
rect 293868 509260 293920 509312
rect 297640 509260 297692 509312
rect 192484 506472 192536 506524
rect 297640 506472 297692 506524
rect 153384 505155 153436 505164
rect 153384 505121 153393 505155
rect 153393 505121 153427 505155
rect 153427 505121 153436 505155
rect 153384 505112 153436 505121
rect 380716 503115 380768 503124
rect 380716 503081 380725 503115
rect 380725 503081 380759 503115
rect 380759 503081 380768 503115
rect 380716 503072 380768 503081
rect 118332 502324 118384 502376
rect 118516 502324 118568 502376
rect 128544 502324 128596 502376
rect 128820 502324 128872 502376
rect 153384 502367 153436 502376
rect 153384 502333 153393 502367
rect 153393 502333 153427 502367
rect 153427 502333 153436 502367
rect 153384 502324 153436 502333
rect 96528 500896 96580 500948
rect 380440 500896 380492 500948
rect 103520 500828 103572 500880
rect 104808 500828 104860 500880
rect 380440 500760 380492 500812
rect 380716 500760 380768 500812
rect 70216 500216 70268 500268
rect 95240 500216 95292 500268
rect 96528 500216 96580 500268
rect 300492 499128 300544 499180
rect 311900 499128 311952 499180
rect 298928 499060 298980 499112
rect 310612 499060 310664 499112
rect 324228 499060 324280 499112
rect 378416 499060 378468 499112
rect 299020 498992 299072 499044
rect 314844 498992 314896 499044
rect 321468 498992 321520 499044
rect 378508 498992 378560 499044
rect 298652 498924 298704 498976
rect 316040 498924 316092 498976
rect 317328 498924 317380 498976
rect 378876 498924 378928 498976
rect 298836 498856 298888 498908
rect 309140 498856 309192 498908
rect 310428 498856 310480 498908
rect 378692 498856 378744 498908
rect 298468 498788 298520 498840
rect 306472 498788 306524 498840
rect 309048 498788 309100 498840
rect 378600 498788 378652 498840
rect 298560 498244 298612 498296
rect 302424 498244 302476 498296
rect 132132 498176 132184 498228
rect 580172 498176 580224 498228
rect 129096 498108 129148 498160
rect 364248 498108 364300 498160
rect 116032 498040 116084 498092
rect 347320 498040 347372 498092
rect 120724 497972 120776 498024
rect 121368 497972 121420 498024
rect 338856 497972 338908 498024
rect 111708 497904 111760 497956
rect 115296 497904 115348 497956
rect 313280 497904 313332 497956
rect 320088 497904 320140 497956
rect 357992 497904 358044 497956
rect 144184 497836 144236 497888
rect 334440 497836 334492 497888
rect 338764 497836 338816 497888
rect 362224 497836 362276 497888
rect 284116 497768 284168 497820
rect 368480 497768 368532 497820
rect 291016 497700 291068 497752
rect 377128 497700 377180 497752
rect 284208 497632 284260 497684
rect 374920 497632 374972 497684
rect 108948 497564 109000 497616
rect 116032 497564 116084 497616
rect 118056 497564 118108 497616
rect 302608 497564 302660 497616
rect 304540 497564 304592 497616
rect 366456 497564 366508 497616
rect 83924 497496 83976 497548
rect 127072 497496 127124 497548
rect 360016 497496 360068 497548
rect 111800 497428 111852 497480
rect 125876 497428 125928 497480
rect 372712 497428 372764 497480
rect 285588 497360 285640 497412
rect 345112 497360 345164 497412
rect 292304 497292 292356 497344
rect 351552 497292 351604 497344
rect 277308 497224 277360 497276
rect 317512 497224 317564 497276
rect 337384 497224 337436 497276
rect 355784 497224 355836 497276
rect 276664 497156 276716 497208
rect 311072 497156 311124 497208
rect 315948 497156 316000 497208
rect 349344 497156 349396 497208
rect 321744 497088 321796 497140
rect 301504 497020 301556 497072
rect 325976 497020 326028 497072
rect 286416 496952 286468 497004
rect 306840 496952 306892 497004
rect 308956 496952 309008 497004
rect 321744 496952 321796 497004
rect 305644 496884 305696 496936
rect 323952 496884 324004 496936
rect 302148 496816 302200 496868
rect 302608 496816 302660 496868
rect 308404 496816 308456 496868
rect 315304 496816 315356 496868
rect 330484 496816 330536 496868
rect 336648 496816 336700 496868
rect 340144 496816 340196 496868
rect 343088 496816 343140 496868
rect 3332 495456 3384 495508
rect 31024 495456 31076 495508
rect 153384 495388 153436 495440
rect 153568 495388 153620 495440
rect 288348 492711 288400 492720
rect 288348 492677 288357 492711
rect 288357 492677 288391 492711
rect 288391 492677 288400 492711
rect 288348 492668 288400 492677
rect 118332 492600 118384 492652
rect 118516 492600 118568 492652
rect 128544 492600 128596 492652
rect 128728 492600 128780 492652
rect 153292 492600 153344 492652
rect 153568 492600 153620 492652
rect 288348 485868 288400 485920
rect 288256 485664 288308 485716
rect 299940 485800 299992 485852
rect 300584 485800 300636 485852
rect 304172 485800 304224 485852
rect 438216 485800 438268 485852
rect 580172 485800 580224 485852
rect 304264 485664 304316 485716
rect 288256 482987 288308 482996
rect 288256 482953 288265 482987
rect 288265 482953 288299 482987
rect 288299 482953 288308 482987
rect 288256 482944 288308 482953
rect 304264 482944 304316 482996
rect 304448 482944 304500 482996
rect 4068 480632 4120 480684
rect 4988 480632 5040 480684
rect 153292 476076 153344 476128
rect 153476 476076 153528 476128
rect 299756 476076 299808 476128
rect 299940 476076 299992 476128
rect 288256 476051 288308 476060
rect 288256 476017 288265 476051
rect 288265 476017 288299 476051
rect 288299 476017 288308 476051
rect 288256 476008 288308 476017
rect 299848 473331 299900 473340
rect 299848 473297 299857 473331
rect 299857 473297 299891 473331
rect 299891 473297 299900 473331
rect 299848 473288 299900 473297
rect 304264 473288 304316 473340
rect 304356 473288 304408 473340
rect 118424 466488 118476 466540
rect 288348 466488 288400 466540
rect 153384 466420 153436 466472
rect 118332 466352 118384 466404
rect 153476 466352 153528 466404
rect 299848 466395 299900 466404
rect 299848 466361 299857 466395
rect 299857 466361 299891 466395
rect 299891 466361 299900 466395
rect 299848 466352 299900 466361
rect 288256 463811 288308 463820
rect 288256 463777 288265 463811
rect 288265 463777 288299 463811
rect 288299 463777 288308 463811
rect 288256 463768 288308 463777
rect 118056 463632 118108 463684
rect 118332 463632 118384 463684
rect 153476 463675 153528 463684
rect 153476 463641 153485 463675
rect 153485 463641 153519 463675
rect 153519 463641 153528 463675
rect 153476 463632 153528 463641
rect 288256 463675 288308 463684
rect 288256 463641 288265 463675
rect 288265 463641 288299 463675
rect 288299 463641 288308 463675
rect 288256 463632 288308 463641
rect 133144 462340 133196 462392
rect 579804 462340 579856 462392
rect 304264 456832 304316 456884
rect 299756 456764 299808 456816
rect 299940 456764 299992 456816
rect 153476 456739 153528 456748
rect 153476 456705 153485 456739
rect 153485 456705 153519 456739
rect 153519 456705 153528 456739
rect 153476 456696 153528 456705
rect 288256 456739 288308 456748
rect 288256 456705 288265 456739
rect 288265 456705 288299 456739
rect 288299 456705 288308 456739
rect 288256 456696 288308 456705
rect 304264 456696 304316 456748
rect 299848 454019 299900 454028
rect 299848 453985 299857 454019
rect 299857 453985 299891 454019
rect 299891 453985 299900 454019
rect 299848 453976 299900 453985
rect 304264 453976 304316 454028
rect 304356 453976 304408 454028
rect 304356 452548 304408 452600
rect 3056 451324 3108 451376
rect 267280 451324 267332 451376
rect 133236 451256 133288 451308
rect 580172 451256 580224 451308
rect 288348 447219 288400 447228
rect 288348 447185 288357 447219
rect 288357 447185 288391 447219
rect 288391 447185 288400 447219
rect 288348 447176 288400 447185
rect 118240 447108 118292 447160
rect 153384 447108 153436 447160
rect 153568 447108 153620 447160
rect 118332 447040 118384 447092
rect 299848 447083 299900 447092
rect 299848 447049 299857 447083
rect 299857 447049 299891 447083
rect 299891 447049 299900 447083
rect 299848 447040 299900 447049
rect 288348 444431 288400 444440
rect 288348 444397 288357 444431
rect 288357 444397 288391 444431
rect 288391 444397 288400 444431
rect 288348 444388 288400 444397
rect 118056 444320 118108 444372
rect 118332 444320 118384 444372
rect 153384 444363 153436 444372
rect 153384 444329 153393 444363
rect 153393 444329 153427 444363
rect 153427 444329 153436 444363
rect 153384 444320 153436 444329
rect 288256 444363 288308 444372
rect 288256 444329 288265 444363
rect 288265 444329 288299 444363
rect 288299 444329 288308 444363
rect 288256 444320 288308 444329
rect 436744 438880 436796 438932
rect 580172 438880 580224 438932
rect 299756 437452 299808 437504
rect 299940 437452 299992 437504
rect 153384 437427 153436 437436
rect 153384 437393 153393 437427
rect 153393 437393 153427 437427
rect 153427 437393 153436 437427
rect 153384 437384 153436 437393
rect 288256 437427 288308 437436
rect 288256 437393 288265 437427
rect 288265 437393 288299 437427
rect 288299 437393 288308 437427
rect 288256 437384 288308 437393
rect 304172 434775 304224 434784
rect 304172 434741 304181 434775
rect 304181 434741 304215 434775
rect 304215 434741 304224 434775
rect 304172 434732 304224 434741
rect 299848 434707 299900 434716
rect 299848 434673 299857 434707
rect 299857 434673 299891 434707
rect 299891 434673 299900 434707
rect 299848 434664 299900 434673
rect 288348 427907 288400 427916
rect 288348 427873 288357 427907
rect 288357 427873 288391 427907
rect 288391 427873 288400 427907
rect 288348 427864 288400 427873
rect 118240 427796 118292 427848
rect 118332 427728 118384 427780
rect 299848 427771 299900 427780
rect 299848 427737 299857 427771
rect 299857 427737 299891 427771
rect 299891 427737 299900 427771
rect 299848 427728 299900 427737
rect 288348 425119 288400 425128
rect 288348 425085 288357 425119
rect 288357 425085 288391 425119
rect 288391 425085 288400 425119
rect 288348 425076 288400 425085
rect 288072 425008 288124 425060
rect 288256 425008 288308 425060
rect 4068 423648 4120 423700
rect 5080 423648 5132 423700
rect 153292 418208 153344 418260
rect 299756 418140 299808 418192
rect 299940 418140 299992 418192
rect 304264 418208 304316 418260
rect 153200 418072 153252 418124
rect 304172 418072 304224 418124
rect 132960 415420 133012 415472
rect 579804 415420 579856 415472
rect 118424 415395 118476 415404
rect 118424 415361 118433 415395
rect 118433 415361 118467 415395
rect 118467 415361 118476 415395
rect 118424 415352 118476 415361
rect 128636 415352 128688 415404
rect 299848 415395 299900 415404
rect 299848 415361 299857 415395
rect 299857 415361 299891 415395
rect 299891 415361 299900 415395
rect 299848 415352 299900 415361
rect 248972 410796 249024 410848
rect 266544 410796 266596 410848
rect 246028 410728 246080 410780
rect 267740 410728 267792 410780
rect 234620 410660 234672 410712
rect 266636 410660 266688 410712
rect 228916 410592 228968 410644
rect 267004 410592 267056 410644
rect 223396 410524 223448 410576
rect 266912 410524 266964 410576
rect 211988 410456 212040 410508
rect 267096 410456 267148 410508
rect 206284 410388 206336 410440
rect 266360 410388 266412 410440
rect 243268 410320 243320 410372
rect 266820 410320 266872 410372
rect 240324 410252 240376 410304
rect 266728 410252 266780 410304
rect 237564 410184 237616 410236
rect 267648 410184 267700 410236
rect 196900 410116 196952 410168
rect 200580 410116 200632 410168
rect 257436 410116 257488 410168
rect 268752 410116 268804 410168
rect 199752 410048 199804 410100
rect 217692 410048 217744 410100
rect 254676 410048 254728 410100
rect 268844 410048 268896 410100
rect 199936 409980 199988 410032
rect 220452 409980 220504 410032
rect 251732 409980 251784 410032
rect 266452 409980 266504 410032
rect 200028 409912 200080 409964
rect 214748 409912 214800 409964
rect 260380 409912 260432 409964
rect 267556 409912 267608 409964
rect 199844 409844 199896 409896
rect 209044 409844 209096 409896
rect 265900 409844 265952 409896
rect 268936 409844 268988 409896
rect 199568 409640 199620 409692
rect 202880 409640 202932 409692
rect 199660 409572 199712 409624
rect 205640 409572 205692 409624
rect 196808 409504 196860 409556
rect 209780 409504 209832 409556
rect 195704 409436 195756 409488
rect 212540 409436 212592 409488
rect 195796 409368 195848 409420
rect 215300 409368 215352 409420
rect 196716 409300 196768 409352
rect 222752 409300 222804 409352
rect 196624 409232 196676 409284
rect 222844 409232 222896 409284
rect 195612 409164 195664 409216
rect 222200 409164 222252 409216
rect 195520 409096 195572 409148
rect 222292 409096 222344 409148
rect 153200 408484 153252 408536
rect 153384 408416 153436 408468
rect 287980 408348 288032 408400
rect 288348 408348 288400 408400
rect 380624 407872 380676 407924
rect 70124 407804 70176 407856
rect 104808 407804 104860 407856
rect 416964 407804 417016 407856
rect 71596 407736 71648 407788
rect 85580 407736 85632 407788
rect 402980 407736 403032 407788
rect 198004 407192 198056 407244
rect 411260 407192 411312 407244
rect 130384 407124 130436 407176
rect 416872 407124 416924 407176
rect 295340 406716 295392 406768
rect 197728 406512 197780 406564
rect 295340 405832 295392 405884
rect 295984 405832 296036 405884
rect 118516 405696 118568 405748
rect 128544 405739 128596 405748
rect 128544 405705 128553 405739
rect 128553 405705 128587 405739
rect 128587 405705 128596 405739
rect 128544 405696 128596 405705
rect 132868 405739 132920 405748
rect 132868 405705 132877 405739
rect 132877 405705 132911 405739
rect 132911 405705 132920 405739
rect 132868 405696 132920 405705
rect 299940 405696 299992 405748
rect 128544 404311 128596 404320
rect 128544 404277 128553 404311
rect 128553 404277 128587 404311
rect 128587 404277 128596 404311
rect 128544 404268 128596 404277
rect 153384 398939 153436 398948
rect 153384 398905 153393 398939
rect 153393 398905 153427 398939
rect 153427 398905 153436 398939
rect 153384 398896 153436 398905
rect 304264 398896 304316 398948
rect 71688 398828 71740 398880
rect 85488 398828 85540 398880
rect 120908 398828 120960 398880
rect 121368 398828 121420 398880
rect 125692 398828 125744 398880
rect 117320 398760 117372 398812
rect 118608 398760 118660 398812
rect 129740 398760 129792 398812
rect 132684 398760 132736 398812
rect 132868 398760 132920 398812
rect 304264 398760 304316 398812
rect 85488 398692 85540 398744
rect 90272 398692 90324 398744
rect 129740 398284 129792 398336
rect 130384 398284 130436 398336
rect 100668 398216 100720 398268
rect 113824 398216 113876 398268
rect 129464 398216 129516 398268
rect 85948 398148 86000 398200
rect 117320 398148 117372 398200
rect 75828 398080 75880 398132
rect 115940 398080 115992 398132
rect 127164 398080 127216 398132
rect 133052 398080 133104 398132
rect 175924 398080 175976 398132
rect 80796 397808 80848 397860
rect 126152 397808 126204 397860
rect 126336 397808 126388 397860
rect 115848 397740 115900 397792
rect 126428 397740 126480 397792
rect 110972 397672 111024 397724
rect 111708 397672 111760 397724
rect 127256 397672 127308 397724
rect 106004 397604 106056 397656
rect 127624 397604 127676 397656
rect 95884 397536 95936 397588
rect 133052 397536 133104 397588
rect 125600 397468 125652 397520
rect 144184 397468 144236 397520
rect 129464 397400 129516 397452
rect 198004 397400 198056 397452
rect 69940 396720 69992 396772
rect 117964 396720 118016 396772
rect 126520 396720 126572 396772
rect 153384 396083 153436 396092
rect 153384 396049 153393 396083
rect 153393 396049 153427 396083
rect 153427 396049 153436 396083
rect 153384 396040 153436 396049
rect 299848 396040 299900 396092
rect 299940 396040 299992 396092
rect 153384 395904 153436 395956
rect 84016 395836 84068 395888
rect 84108 395700 84160 395752
rect 70032 395632 70084 395684
rect 108948 395632 109000 395684
rect 125784 395632 125836 395684
rect 168656 395564 168708 395616
rect 179512 395496 179564 395548
rect 128636 394680 128688 394732
rect 402980 393252 403032 393304
rect 403900 393252 403952 393304
rect 288164 391892 288216 391944
rect 288348 391892 288400 391944
rect 69664 390532 69716 390584
rect 71596 390532 71648 390584
rect 416596 389376 416648 389428
rect 464252 389376 464304 389428
rect 414664 389308 414716 389360
rect 475844 389308 475896 389360
rect 132868 389240 132920 389292
rect 418068 389240 418120 389292
rect 487436 389240 487488 389292
rect 304264 389172 304316 389224
rect 416688 389172 416740 389224
rect 499028 389172 499080 389224
rect 132868 389104 132920 389156
rect 153292 389147 153344 389156
rect 153292 389113 153301 389147
rect 153301 389113 153335 389147
rect 153335 389113 153344 389147
rect 153292 389104 153344 389113
rect 304172 389104 304224 389156
rect 128728 388424 128780 388476
rect 375288 387064 375340 387116
rect 478880 387064 478932 387116
rect 304264 386359 304316 386368
rect 304264 386325 304273 386359
rect 304273 386325 304307 386359
rect 304307 386325 304316 386359
rect 304264 386316 304316 386325
rect 344928 385772 344980 385824
rect 408868 385772 408920 385824
rect 295984 385704 296036 385756
rect 388260 385704 388312 385756
rect 267280 385636 267332 385688
rect 436100 385636 436152 385688
rect 369124 385568 369176 385620
rect 392860 385568 392912 385620
rect 349068 385500 349120 385552
rect 385868 385500 385920 385552
rect 355876 385432 355928 385484
rect 399668 385432 399720 385484
rect 357348 385364 357400 385416
rect 406660 385364 406712 385416
rect 353208 385296 353260 385348
rect 402060 385296 402112 385348
rect 347688 385228 347740 385280
rect 397460 385228 397512 385280
rect 343548 385160 343600 385212
rect 395068 385160 395120 385212
rect 355968 385092 356020 385144
rect 413468 385092 413520 385144
rect 367008 385024 367060 385076
rect 390468 385024 390520 385076
rect 126520 384276 126572 384328
rect 140780 384276 140832 384328
rect 126152 383664 126204 383716
rect 126336 383664 126388 383716
rect 301596 381488 301648 381540
rect 302148 381488 302200 381540
rect 380900 381488 380952 381540
rect 153292 379448 153344 379500
rect 153476 379448 153528 379500
rect 304264 379355 304316 379364
rect 304264 379321 304273 379355
rect 304273 379321 304307 379355
rect 304307 379321 304316 379355
rect 304264 379312 304316 379321
rect 132776 376796 132828 376848
rect 132868 376796 132920 376848
rect 128912 376728 128964 376780
rect 299848 376728 299900 376780
rect 299940 376728 299992 376780
rect 351828 376728 351880 376780
rect 380900 376728 380952 376780
rect 132684 375343 132736 375352
rect 132684 375309 132693 375343
rect 132693 375309 132727 375343
rect 132727 375309 132736 375343
rect 132684 375300 132736 375309
rect 126336 374076 126388 374128
rect 126152 374008 126204 374060
rect 364248 374008 364300 374060
rect 380900 374008 380952 374060
rect 416044 374008 416096 374060
rect 456800 374008 456852 374060
rect 288348 372580 288400 372632
rect 288532 372580 288584 372632
rect 288348 369903 288400 369912
rect 288348 369869 288357 369903
rect 288357 369869 288391 369903
rect 288391 369869 288400 369903
rect 288348 369860 288400 369869
rect 304264 369860 304316 369912
rect 347596 369860 347648 369912
rect 380900 369860 380952 369912
rect 304172 369792 304224 369844
rect 133052 367004 133104 367056
rect 133144 367047 133196 367056
rect 133144 367013 133153 367047
rect 133153 367013 133187 367047
rect 133187 367013 133196 367047
rect 133144 367004 133196 367013
rect 153568 367004 153620 367056
rect 132776 366936 132828 366988
rect 132960 366868 133012 366920
rect 133052 366800 133104 366852
rect 132960 366732 133012 366784
rect 2780 365712 2832 365764
rect 5172 365712 5224 365764
rect 129372 365644 129424 365696
rect 197728 365644 197780 365696
rect 126152 364352 126204 364404
rect 126336 364352 126388 364404
rect 288348 362967 288400 362976
rect 288348 362933 288357 362967
rect 288357 362933 288391 362967
rect 288391 362933 288400 362967
rect 288348 362924 288400 362933
rect 333888 362924 333940 362976
rect 380900 362924 380952 362976
rect 132776 360204 132828 360256
rect 288348 360247 288400 360256
rect 288348 360213 288357 360247
rect 288357 360213 288391 360247
rect 288391 360213 288400 360247
rect 288348 360204 288400 360213
rect 304172 360204 304224 360256
rect 304264 360136 304316 360188
rect 132776 360068 132828 360120
rect 133144 358683 133196 358692
rect 133144 358649 133153 358683
rect 133153 358649 133187 358683
rect 133187 358649 133196 358683
rect 133144 358640 133196 358649
rect 153476 357459 153528 357468
rect 153476 357425 153485 357459
rect 153485 357425 153519 357459
rect 153519 357425 153528 357459
rect 153476 357416 153528 357425
rect 144184 357348 144236 357400
rect 145564 357348 145616 357400
rect 304264 357255 304316 357264
rect 304264 357221 304273 357255
rect 304273 357221 304307 357255
rect 304307 357221 304316 357255
rect 304264 357212 304316 357221
rect 126336 354764 126388 354816
rect 126152 354696 126204 354748
rect 288348 353311 288400 353320
rect 288348 353277 288357 353311
rect 288357 353277 288391 353311
rect 288391 353277 288400 353311
rect 288348 353268 288400 353277
rect 354588 353268 354640 353320
rect 380900 353268 380952 353320
rect 129004 351160 129056 351212
rect 129832 351160 129884 351212
rect 130384 351160 130436 351212
rect 153476 350548 153528 350600
rect 153384 350480 153436 350532
rect 299848 350480 299900 350532
rect 299940 350412 299992 350464
rect 304264 347871 304316 347880
rect 304264 347837 304273 347871
rect 304273 347837 304307 347871
rect 304307 347837 304316 347871
rect 304264 347828 304316 347837
rect 132684 347760 132736 347812
rect 132868 347760 132920 347812
rect 381544 347692 381596 347744
rect 386788 347692 386840 347744
rect 360108 347624 360160 347676
rect 391388 347624 391440 347676
rect 362868 347556 362920 347608
rect 398196 347556 398248 347608
rect 358728 347488 358780 347540
rect 393596 347488 393648 347540
rect 362776 347420 362828 347472
rect 402796 347420 402848 347472
rect 350448 347352 350500 347404
rect 395988 347352 396040 347404
rect 342168 347284 342220 347336
rect 388996 347284 389048 347336
rect 361488 347216 361540 347268
rect 407396 347216 407448 347268
rect 354496 347148 354548 347200
rect 400588 347148 400640 347200
rect 361396 347080 361448 347132
rect 414388 347080 414440 347132
rect 333796 347012 333848 347064
rect 411996 347012 412048 347064
rect 126152 345040 126204 345092
rect 126336 345040 126388 345092
rect 504824 345040 504876 345092
rect 579988 345040 580040 345092
rect 288348 344564 288400 344616
rect 129004 342864 129056 342916
rect 130660 342864 130712 342916
rect 192484 342864 192536 342916
rect 199292 342864 199344 342916
rect 200212 342864 200264 342916
rect 130292 342048 130344 342100
rect 132684 342048 132736 342100
rect 132500 341980 132552 342032
rect 503812 341980 503864 342032
rect 504180 341980 504232 342032
rect 132500 341844 132552 341896
rect 131948 341640 132000 341692
rect 580632 341640 580684 341692
rect 132040 341572 132092 341624
rect 580816 341572 580868 341624
rect 131672 341504 131724 341556
rect 580724 341504 580776 341556
rect 153384 341003 153436 341012
rect 153384 340969 153393 341003
rect 153393 340969 153427 341003
rect 153427 340969 153436 341003
rect 153384 340960 153436 340969
rect 127256 340824 127308 340876
rect 408500 340824 408552 340876
rect 127164 340756 127216 340808
rect 404360 340756 404412 340808
rect 503904 340756 503956 340808
rect 504732 340824 504784 340876
rect 127716 340688 127768 340740
rect 381728 340688 381780 340740
rect 130384 340620 130436 340672
rect 381636 340620 381688 340672
rect 132868 340595 132920 340604
rect 132868 340561 132877 340595
rect 132877 340561 132911 340595
rect 132911 340561 132920 340595
rect 132868 340552 132920 340561
rect 140780 340552 140832 340604
rect 383660 340552 383712 340604
rect 145564 340484 145616 340536
rect 381820 340484 381872 340536
rect 153384 340459 153436 340468
rect 153384 340425 153393 340459
rect 153393 340425 153427 340459
rect 153427 340425 153436 340459
rect 153384 340416 153436 340425
rect 111708 340212 111760 340264
rect 127256 340212 127308 340264
rect 110328 340144 110380 340196
rect 127164 340144 127216 340196
rect 130752 340144 130804 340196
rect 140780 340144 140832 340196
rect 130384 339668 130436 339720
rect 130844 339668 130896 339720
rect 262128 339124 262180 339176
rect 268936 339124 268988 339176
rect 198096 338988 198148 339040
rect 209964 338988 210016 339040
rect 199476 338920 199528 338972
rect 214104 338920 214156 338972
rect 257712 338920 257764 338972
rect 267556 338920 267608 338972
rect 199384 338852 199436 338904
rect 215300 338852 215352 338904
rect 253664 338852 253716 338904
rect 268844 338852 268896 338904
rect 198280 338784 198332 338836
rect 220820 338784 220872 338836
rect 244188 338784 244240 338836
rect 268752 338784 268804 338836
rect 198188 338716 198240 338768
rect 222200 338716 222252 338768
rect 237288 338716 237340 338768
rect 267648 338716 267700 338768
rect 128912 338104 128964 338156
rect 129004 338104 129056 338156
rect 288348 338104 288400 338156
rect 107568 338036 107620 338088
rect 301596 338036 301648 338088
rect 97908 337968 97960 338020
rect 126980 337968 127032 338020
rect 132960 337968 133012 338020
rect 133052 337968 133104 338020
rect 133144 338011 133196 338020
rect 133144 337977 133153 338011
rect 133153 337977 133187 338011
rect 133187 337977 133196 338011
rect 133144 337968 133196 337977
rect 220452 337968 220504 338020
rect 238116 337968 238168 338020
rect 244924 337968 244976 338020
rect 112812 337900 112864 337952
rect 113088 337900 113140 337952
rect 127072 337900 127124 337952
rect 209044 337900 209096 337952
rect 220084 337900 220136 337952
rect 226156 337900 226208 337952
rect 248696 337900 248748 337952
rect 250996 337900 251048 337952
rect 260196 337900 260248 337952
rect 122748 337832 122800 337884
rect 127716 337832 127768 337884
rect 132960 337832 133012 337884
rect 133052 337832 133104 337884
rect 203340 337832 203392 337884
rect 215944 337832 215996 337884
rect 217508 337832 217560 337884
rect 241428 337832 241480 337884
rect 246028 337832 246080 337884
rect 253756 337832 253808 337884
rect 263140 337832 263192 337884
rect 200580 337764 200632 337816
rect 234620 337764 234672 337816
rect 237748 337764 237800 337816
rect 240048 337764 240100 337816
rect 243084 337764 243136 337816
rect 247684 337764 247736 337816
rect 257436 337764 257488 337816
rect 92756 337696 92808 337748
rect 93768 337696 93820 337748
rect 102876 337696 102928 337748
rect 103428 337696 103480 337748
rect 214748 337696 214800 337748
rect 258724 337696 258776 337748
rect 206100 337628 206152 337680
rect 251732 337628 251784 337680
rect 252468 337628 252520 337680
rect 72884 337560 72936 337612
rect 134064 337560 134116 337612
rect 299940 337560 299992 337612
rect 401508 337560 401560 337612
rect 460572 337560 460624 337612
rect 117964 337492 118016 337544
rect 124128 337492 124180 337544
rect 297364 337492 297416 337544
rect 411168 337492 411220 337544
rect 472164 337492 472216 337544
rect 77852 337424 77904 337476
rect 99288 337424 99340 337476
rect 329840 337424 329892 337476
rect 408408 337424 408460 337476
rect 483756 337424 483808 337476
rect 87788 337356 87840 337408
rect 128268 337356 128320 337408
rect 380532 337356 380584 337408
rect 413928 337356 413980 337408
rect 495348 337356 495400 337408
rect 231860 337288 231912 337340
rect 248788 337288 248840 337340
rect 255320 337288 255372 337340
rect 228916 337220 228968 337272
rect 232504 337220 232556 337272
rect 237564 337220 237616 337272
rect 243084 337220 243136 337272
rect 238024 337152 238076 337204
rect 223212 336812 223264 336864
rect 229744 336812 229796 336864
rect 244096 336812 244148 336864
rect 248604 336812 248656 336864
rect 254492 336812 254544 336864
rect 258264 336812 258316 336864
rect 2964 336744 3016 336796
rect 434904 336744 434956 336796
rect 82728 336676 82780 336728
rect 125876 336676 125928 336728
rect 257712 336676 257764 336728
rect 257804 336676 257856 336728
rect 126152 335316 126204 335368
rect 126336 335316 126388 335368
rect 257804 335248 257856 335300
rect 133144 333319 133196 333328
rect 133144 333285 133153 333319
rect 133153 333285 133187 333319
rect 133187 333285 133196 333319
rect 133144 333276 133196 333285
rect 288348 332027 288400 332036
rect 288348 331993 288357 332027
rect 288357 331993 288391 332027
rect 288391 331993 288400 332027
rect 288348 331984 288400 331993
rect 214012 331304 214064 331356
rect 503812 331236 503864 331288
rect 503628 331168 503680 331220
rect 503996 331168 504048 331220
rect 503720 328559 503772 328568
rect 503720 328525 503729 328559
rect 503729 328525 503763 328559
rect 503763 328525 503772 328559
rect 503720 328516 503772 328525
rect 209780 328448 209832 328500
rect 209964 328448 210016 328500
rect 213920 328491 213972 328500
rect 213920 328457 213929 328491
rect 213929 328457 213963 328491
rect 213963 328457 213972 328491
rect 213920 328448 213972 328457
rect 288164 328448 288216 328500
rect 129004 328423 129056 328432
rect 129004 328389 129013 328423
rect 129013 328389 129047 328423
rect 129047 328389 129056 328423
rect 129004 328380 129056 328389
rect 504272 328380 504324 328432
rect 504364 328380 504416 328432
rect 288164 328355 288216 328364
rect 288164 328321 288173 328355
rect 288173 328321 288207 328355
rect 288207 328321 288216 328355
rect 288164 328312 288216 328321
rect 504272 327063 504324 327072
rect 504272 327029 504281 327063
rect 504281 327029 504315 327063
rect 504315 327029 504324 327063
rect 504272 327020 504324 327029
rect 126152 325660 126204 325712
rect 126336 325660 126388 325712
rect 503904 321759 503956 321768
rect 503904 321725 503913 321759
rect 503913 321725 503947 321759
rect 503947 321725 503956 321759
rect 503904 321716 503956 321725
rect 503720 321691 503772 321700
rect 503720 321657 503729 321691
rect 503729 321657 503763 321691
rect 503763 321657 503772 321691
rect 503720 321648 503772 321657
rect 503996 321691 504048 321700
rect 503996 321657 504005 321691
rect 504005 321657 504039 321691
rect 504039 321657 504048 321691
rect 503996 321648 504048 321657
rect 132776 321580 132828 321632
rect 579620 321580 579672 321632
rect 503904 321555 503956 321564
rect 503904 321521 503913 321555
rect 503913 321521 503947 321555
rect 503947 321521 503956 321555
rect 503904 321512 503956 321521
rect 128820 318860 128872 318912
rect 153384 318792 153436 318844
rect 153476 318792 153528 318844
rect 288348 318792 288400 318844
rect 503996 318835 504048 318844
rect 503996 318801 504005 318835
rect 504005 318801 504039 318835
rect 504039 318801 504048 318835
rect 503996 318792 504048 318801
rect 209780 318767 209832 318776
rect 209780 318733 209789 318767
rect 209789 318733 209823 318767
rect 209823 318733 209832 318767
rect 209780 318724 209832 318733
rect 304264 318767 304316 318776
rect 304264 318733 304273 318767
rect 304273 318733 304307 318767
rect 304307 318733 304316 318767
rect 304264 318724 304316 318733
rect 257712 317475 257764 317484
rect 257712 317441 257721 317475
rect 257721 317441 257755 317475
rect 257755 317441 257764 317475
rect 257712 317432 257764 317441
rect 503720 317475 503772 317484
rect 503720 317441 503729 317475
rect 503729 317441 503763 317475
rect 503763 317441 503772 317475
rect 503720 317432 503772 317441
rect 504364 317432 504416 317484
rect 128912 317364 128964 317416
rect 126152 316004 126204 316056
rect 126336 316004 126388 316056
rect 288348 313395 288400 313404
rect 288348 313361 288357 313395
rect 288357 313361 288391 313395
rect 288391 313361 288400 313395
rect 288348 313352 288400 313361
rect 504364 312647 504416 312656
rect 504364 312613 504373 312647
rect 504373 312613 504407 312647
rect 504407 312613 504416 312647
rect 504364 312604 504416 312613
rect 153384 311924 153436 311976
rect 153476 311924 153528 311976
rect 503628 311856 503680 311908
rect 503996 311856 504048 311908
rect 503628 311720 503680 311772
rect 503996 311720 504048 311772
rect 131856 310496 131908 310548
rect 579712 310496 579764 310548
rect 304264 309247 304316 309256
rect 304264 309213 304273 309247
rect 304273 309213 304307 309247
rect 304307 309213 304316 309247
rect 304264 309204 304316 309213
rect 209780 309179 209832 309188
rect 209780 309145 209789 309179
rect 209789 309145 209823 309179
rect 209823 309145 209832 309179
rect 209780 309136 209832 309145
rect 288348 309179 288400 309188
rect 288348 309145 288357 309179
rect 288357 309145 288391 309179
rect 288391 309145 288400 309179
rect 288348 309136 288400 309145
rect 304264 309111 304316 309120
rect 304264 309077 304273 309111
rect 304273 309077 304307 309111
rect 304307 309077 304316 309111
rect 304264 309068 304316 309077
rect 132684 308252 132736 308304
rect 132868 308252 132920 308304
rect 4068 307776 4120 307828
rect 5264 307776 5316 307828
rect 128636 307819 128688 307828
rect 128636 307785 128645 307819
rect 128645 307785 128679 307819
rect 128679 307785 128688 307819
rect 128636 307776 128688 307785
rect 257804 307751 257856 307760
rect 257804 307717 257813 307751
rect 257813 307717 257847 307751
rect 257847 307717 257856 307751
rect 257804 307708 257856 307717
rect 153292 302200 153344 302252
rect 153476 302200 153528 302252
rect 288348 302243 288400 302252
rect 288348 302209 288357 302243
rect 288357 302209 288391 302243
rect 288391 302209 288400 302243
rect 288348 302200 288400 302209
rect 128636 302064 128688 302116
rect 128912 302064 128964 302116
rect 304264 301699 304316 301708
rect 304264 301665 304273 301699
rect 304273 301665 304307 301699
rect 304307 301665 304316 301699
rect 304264 301656 304316 301665
rect 288348 299523 288400 299532
rect 288348 299489 288357 299523
rect 288357 299489 288391 299523
rect 288391 299489 288400 299523
rect 288348 299480 288400 299489
rect 503628 299480 503680 299532
rect 503812 299480 503864 299532
rect 504456 299480 504508 299532
rect 209780 299455 209832 299464
rect 209780 299421 209789 299455
rect 209789 299421 209823 299455
rect 209823 299421 209832 299455
rect 209780 299412 209832 299421
rect 304264 299455 304316 299464
rect 304264 299421 304273 299455
rect 304273 299421 304307 299455
rect 304307 299421 304316 299455
rect 304264 299412 304316 299421
rect 257896 298120 257948 298172
rect 504456 298095 504508 298104
rect 504456 298061 504465 298095
rect 504465 298061 504499 298095
rect 504499 298061 504508 298095
rect 504456 298052 504508 298061
rect 126152 296692 126204 296744
rect 126336 296692 126388 296744
rect 132684 296080 132736 296132
rect 132868 296080 132920 296132
rect 288348 294083 288400 294092
rect 288348 294049 288357 294083
rect 288357 294049 288391 294083
rect 288391 294049 288400 294083
rect 288348 294040 288400 294049
rect 3332 293972 3384 294024
rect 434536 293972 434588 294024
rect 126060 292476 126112 292528
rect 126336 292476 126388 292528
rect 304264 289935 304316 289944
rect 304264 289901 304273 289935
rect 304273 289901 304307 289935
rect 304307 289901 304316 289935
rect 304264 289892 304316 289901
rect 209780 289867 209832 289876
rect 209780 289833 209789 289867
rect 209789 289833 209823 289867
rect 209823 289833 209832 289867
rect 209780 289824 209832 289833
rect 288164 289824 288216 289876
rect 128820 289799 128872 289808
rect 128820 289765 128829 289799
rect 128829 289765 128863 289799
rect 128863 289765 128872 289799
rect 128820 289756 128872 289765
rect 304264 289799 304316 289808
rect 304264 289765 304273 289799
rect 304273 289765 304307 289799
rect 304307 289765 304316 289799
rect 304264 289756 304316 289765
rect 288164 289731 288216 289740
rect 288164 289697 288173 289731
rect 288173 289697 288207 289731
rect 288207 289697 288216 289731
rect 288164 289688 288216 289697
rect 132684 288940 132736 288992
rect 132868 288940 132920 288992
rect 257804 288396 257856 288448
rect 257896 288396 257948 288448
rect 504548 288396 504600 288448
rect 257804 288303 257856 288312
rect 257804 288269 257813 288303
rect 257813 288269 257847 288303
rect 257847 288269 257856 288303
rect 257804 288260 257856 288269
rect 503720 283024 503772 283076
rect 503812 282956 503864 283008
rect 153292 282888 153344 282940
rect 153476 282888 153528 282940
rect 304264 282795 304316 282804
rect 304264 282761 304273 282795
rect 304273 282761 304307 282795
rect 304307 282761 304316 282795
rect 304264 282752 304316 282761
rect 128912 280168 128964 280220
rect 288348 280168 288400 280220
rect 126152 280100 126204 280152
rect 153384 280143 153436 280152
rect 153384 280109 153393 280143
rect 153393 280109 153427 280143
rect 153427 280109 153436 280143
rect 153384 280100 153436 280109
rect 209780 280143 209832 280152
rect 209780 280109 209789 280143
rect 209789 280109 209823 280143
rect 209823 280109 209832 280143
rect 209780 280100 209832 280109
rect 304264 280143 304316 280152
rect 304264 280109 304273 280143
rect 304273 280109 304307 280143
rect 304307 280109 304316 280143
rect 304264 280100 304316 280109
rect 257896 278740 257948 278792
rect 504456 278715 504508 278724
rect 504456 278681 504465 278715
rect 504465 278681 504499 278715
rect 504499 278681 504508 278715
rect 504456 278672 504508 278681
rect 132868 278060 132920 278112
rect 133512 278060 133564 278112
rect 288348 274771 288400 274780
rect 288348 274737 288357 274771
rect 288357 274737 288391 274771
rect 288391 274737 288400 274771
rect 288348 274728 288400 274737
rect 132684 274660 132736 274712
rect 579620 274660 579672 274712
rect 503628 273300 503680 273352
rect 503996 273300 504048 273352
rect 153568 273232 153620 273284
rect 503628 273164 503680 273216
rect 503996 273164 504048 273216
rect 304264 270623 304316 270632
rect 304264 270589 304273 270623
rect 304273 270589 304307 270623
rect 304307 270589 304316 270623
rect 304264 270580 304316 270589
rect 126060 270555 126112 270564
rect 126060 270521 126069 270555
rect 126069 270521 126103 270555
rect 126103 270521 126112 270555
rect 126060 270512 126112 270521
rect 209780 270555 209832 270564
rect 209780 270521 209789 270555
rect 209789 270521 209823 270555
rect 209823 270521 209832 270555
rect 209780 270512 209832 270521
rect 288164 270512 288216 270564
rect 153568 270487 153620 270496
rect 153568 270453 153577 270487
rect 153577 270453 153611 270487
rect 153611 270453 153620 270487
rect 153568 270444 153620 270453
rect 257804 270487 257856 270496
rect 257804 270453 257813 270487
rect 257813 270453 257847 270487
rect 257847 270453 257856 270487
rect 257804 270444 257856 270453
rect 304264 270444 304316 270496
rect 304448 270444 304500 270496
rect 288164 270419 288216 270428
rect 288164 270385 288173 270419
rect 288173 270385 288207 270419
rect 288207 270385 288216 270419
rect 288164 270376 288216 270385
rect 504640 269084 504692 269136
rect 132868 268404 132920 268456
rect 133512 268404 133564 268456
rect 2780 264936 2832 264988
rect 5448 264936 5500 264988
rect 503720 263644 503772 263696
rect 503996 263644 504048 263696
rect 128912 263619 128964 263628
rect 128912 263585 128921 263619
rect 128921 263585 128955 263619
rect 128955 263585 128964 263619
rect 128912 263576 128964 263585
rect 131580 263576 131632 263628
rect 580172 263576 580224 263628
rect 257804 263551 257856 263560
rect 257804 263517 257813 263551
rect 257813 263517 257847 263551
rect 257847 263517 257856 263551
rect 257804 263508 257856 263517
rect 503720 263508 503772 263560
rect 503996 263508 504048 263560
rect 128912 260899 128964 260908
rect 128912 260865 128921 260899
rect 128921 260865 128955 260899
rect 128955 260865 128964 260899
rect 128912 260856 128964 260865
rect 153660 260856 153712 260908
rect 288348 260856 288400 260908
rect 126152 260788 126204 260840
rect 209780 260831 209832 260840
rect 209780 260797 209789 260831
rect 209789 260797 209823 260831
rect 209823 260797 209832 260831
rect 209780 260788 209832 260797
rect 257804 260831 257856 260840
rect 257804 260797 257813 260831
rect 257813 260797 257847 260831
rect 257847 260797 257856 260831
rect 257804 260788 257856 260797
rect 304080 260831 304132 260840
rect 304080 260797 304089 260831
rect 304089 260797 304123 260831
rect 304123 260797 304132 260831
rect 304080 260788 304132 260797
rect 504272 260831 504324 260840
rect 504272 260797 504281 260831
rect 504281 260797 504315 260831
rect 504315 260797 504324 260831
rect 504272 260788 504324 260797
rect 128728 260720 128780 260772
rect 128912 260720 128964 260772
rect 132868 258748 132920 258800
rect 133512 258748 133564 258800
rect 153660 253988 153712 254040
rect 503628 253988 503680 254040
rect 503996 253988 504048 254040
rect 153568 253852 153620 253904
rect 503628 253852 503680 253904
rect 503996 253852 504048 253904
rect 257804 253827 257856 253836
rect 257804 253793 257813 253827
rect 257813 253793 257847 253827
rect 257847 253793 257856 253827
rect 257804 253784 257856 253793
rect 504272 253827 504324 253836
rect 504272 253793 504281 253827
rect 504281 253793 504315 253827
rect 504315 253793 504324 253827
rect 504272 253784 504324 253793
rect 126060 251311 126112 251320
rect 126060 251277 126069 251311
rect 126069 251277 126103 251311
rect 126103 251277 126112 251311
rect 126060 251268 126112 251277
rect 209780 251311 209832 251320
rect 209780 251277 209789 251311
rect 209789 251277 209823 251311
rect 209823 251277 209832 251311
rect 209780 251268 209832 251277
rect 3332 251200 3384 251252
rect 304264 251200 304316 251252
rect 435088 251200 435140 251252
rect 257804 251132 257856 251184
rect 288256 251175 288308 251184
rect 288256 251141 288265 251175
rect 288265 251141 288299 251175
rect 288299 251141 288308 251175
rect 288256 251132 288308 251141
rect 504272 251175 504324 251184
rect 504272 251141 504281 251175
rect 504281 251141 504315 251175
rect 504315 251141 504324 251175
rect 504272 251132 504324 251141
rect 132868 249092 132920 249144
rect 133512 249092 133564 249144
rect 503720 244400 503772 244452
rect 503812 244332 503864 244384
rect 304172 244307 304224 244316
rect 304172 244273 304181 244307
rect 304181 244273 304215 244307
rect 304215 244273 304224 244307
rect 304172 244264 304224 244273
rect 128820 244196 128872 244248
rect 129004 244196 129056 244248
rect 257712 241519 257764 241528
rect 257712 241485 257721 241519
rect 257721 241485 257755 241519
rect 257755 241485 257764 241519
rect 257712 241476 257764 241485
rect 288348 241476 288400 241528
rect 304172 241519 304224 241528
rect 304172 241485 304181 241519
rect 304181 241485 304215 241519
rect 304215 241485 304224 241519
rect 304172 241476 304224 241485
rect 504456 241476 504508 241528
rect 304172 241383 304224 241392
rect 304172 241349 304181 241383
rect 304181 241349 304215 241383
rect 304215 241349 304224 241383
rect 304172 241340 304224 241349
rect 132868 239436 132920 239488
rect 133512 239436 133564 239488
rect 129004 236759 129056 236768
rect 129004 236725 129013 236759
rect 129013 236725 129047 236759
rect 129047 236725 129056 236759
rect 129004 236716 129056 236725
rect 288348 236011 288400 236020
rect 288348 235977 288357 236011
rect 288357 235977 288391 236011
rect 288391 235977 288400 236011
rect 288348 235968 288400 235977
rect 153292 234676 153344 234728
rect 503628 234676 503680 234728
rect 503996 234676 504048 234728
rect 126152 234608 126204 234660
rect 126336 234608 126388 234660
rect 257712 234608 257764 234660
rect 153292 234540 153344 234592
rect 504456 234676 504508 234728
rect 503628 234540 503680 234592
rect 503996 234540 504048 234592
rect 504364 234540 504416 234592
rect 257804 234472 257856 234524
rect 129004 231931 129056 231940
rect 129004 231897 129013 231931
rect 129013 231897 129047 231931
rect 129047 231897 129056 231931
rect 129004 231888 129056 231897
rect 209780 231820 209832 231872
rect 209964 231820 210016 231872
rect 288164 231820 288216 231872
rect 304172 231863 304224 231872
rect 304172 231829 304181 231863
rect 304181 231829 304215 231863
rect 304215 231829 304224 231863
rect 304172 231820 304224 231829
rect 504364 231795 504416 231804
rect 504364 231761 504373 231795
rect 504373 231761 504407 231795
rect 504407 231761 504416 231795
rect 504364 231752 504416 231761
rect 132868 229712 132920 229764
rect 133512 229712 133564 229764
rect 131304 227740 131356 227792
rect 580172 227740 580224 227792
rect 503720 225088 503772 225140
rect 153200 224995 153252 225004
rect 153200 224961 153209 224995
rect 153209 224961 153243 224995
rect 153243 224961 153252 224995
rect 153200 224952 153252 224961
rect 257804 225020 257856 225072
rect 503812 225020 503864 225072
rect 126152 224884 126204 224936
rect 126336 224884 126388 224936
rect 257712 224884 257764 224936
rect 2964 222164 3016 222216
rect 14464 222164 14516 222216
rect 128636 222164 128688 222216
rect 129004 222164 129056 222216
rect 153200 222207 153252 222216
rect 153200 222173 153209 222207
rect 153209 222173 153243 222207
rect 153243 222173 153252 222207
rect 153200 222164 153252 222173
rect 288348 222164 288400 222216
rect 288532 222164 288584 222216
rect 304356 222164 304408 222216
rect 304540 222164 304592 222216
rect 504456 222164 504508 222216
rect 257712 222028 257764 222080
rect 257988 222028 258040 222080
rect 132868 220056 132920 220108
rect 133512 220056 133564 220108
rect 131488 216656 131540 216708
rect 579620 216656 579672 216708
rect 503628 215364 503680 215416
rect 503996 215364 504048 215416
rect 153200 215296 153252 215348
rect 128636 215160 128688 215212
rect 129004 215160 129056 215212
rect 504456 215364 504508 215416
rect 503628 215228 503680 215280
rect 503996 215228 504048 215280
rect 504272 215228 504324 215280
rect 153292 215160 153344 215212
rect 304172 213392 304224 213444
rect 304356 213392 304408 213444
rect 209780 212508 209832 212560
rect 209964 212508 210016 212560
rect 255320 212508 255372 212560
rect 256240 212508 256292 212560
rect 288072 212508 288124 212560
rect 288164 212508 288216 212560
rect 416412 212508 416464 212560
rect 416688 212508 416740 212560
rect 153292 212483 153344 212492
rect 153292 212449 153301 212483
rect 153301 212449 153335 212483
rect 153335 212449 153344 212483
rect 153292 212440 153344 212449
rect 132868 210400 132920 210452
rect 133512 210400 133564 210452
rect 290924 210400 290976 210452
rect 291108 210400 291160 210452
rect 244004 209720 244056 209772
rect 244188 209720 244240 209772
rect 2964 207000 3016 207052
rect 435180 207000 435232 207052
rect 503720 205776 503772 205828
rect 503812 205708 503864 205760
rect 126428 205683 126480 205692
rect 126428 205649 126437 205683
rect 126437 205649 126471 205683
rect 126471 205649 126480 205683
rect 126428 205640 126480 205649
rect 304080 205683 304132 205692
rect 304080 205649 304089 205683
rect 304089 205649 304123 205683
rect 304123 205649 304132 205683
rect 304080 205640 304132 205649
rect 503720 205640 503772 205692
rect 503996 205640 504048 205692
rect 504180 205683 504232 205692
rect 504180 205649 504189 205683
rect 504189 205649 504223 205683
rect 504223 205649 504232 205683
rect 504180 205640 504232 205649
rect 126428 205547 126480 205556
rect 126428 205513 126437 205547
rect 126437 205513 126471 205547
rect 126471 205513 126480 205547
rect 126428 205504 126480 205513
rect 196716 205300 196768 205352
rect 226892 205300 226944 205352
rect 196624 205232 196676 205284
rect 227904 205232 227956 205284
rect 195888 205164 195940 205216
rect 228640 205164 228692 205216
rect 195704 205096 195756 205148
rect 229560 205096 229612 205148
rect 195796 205028 195848 205080
rect 230480 205028 230532 205080
rect 195520 204960 195572 205012
rect 231216 204960 231268 205012
rect 195612 204892 195664 204944
rect 233240 204892 233292 204944
rect 294420 204212 294472 204264
rect 340880 204212 340932 204264
rect 345756 204212 345808 204264
rect 417056 204212 417108 204264
rect 255780 204144 255832 204196
rect 268200 204144 268252 204196
rect 297916 204144 297968 204196
rect 304264 204144 304316 204196
rect 306656 204144 306708 204196
rect 380440 204144 380492 204196
rect 253572 204076 253624 204128
rect 269028 204076 269080 204128
rect 301412 204076 301464 204128
rect 379612 204076 379664 204128
rect 250536 204008 250588 204060
rect 267924 204008 267976 204060
rect 299020 204008 299072 204060
rect 380348 204008 380400 204060
rect 199016 203940 199068 203992
rect 238760 203940 238812 203992
rect 247592 203940 247644 203992
rect 268108 203940 268160 203992
rect 294880 203940 294932 203992
rect 377404 203940 377456 203992
rect 197728 203872 197780 203924
rect 257160 203872 257212 203924
rect 292212 203872 292264 203924
rect 379796 203872 379848 203924
rect 198004 203804 198056 203856
rect 260380 203804 260432 203856
rect 292488 203804 292540 203856
rect 379888 203804 379940 203856
rect 198464 203736 198516 203788
rect 262772 203736 262824 203788
rect 286968 203736 287020 203788
rect 377312 203736 377364 203788
rect 197452 203668 197504 203720
rect 262956 203668 263008 203720
rect 287520 203668 287572 203720
rect 379704 203668 379756 203720
rect 197820 203600 197872 203652
rect 265256 203600 265308 203652
rect 271788 203600 271840 203652
rect 369860 203600 369912 203652
rect 198372 203532 198424 203584
rect 267556 203532 267608 203584
rect 280528 203532 280580 203584
rect 379980 203532 380032 203584
rect 313556 203464 313608 203516
rect 379520 203464 379572 203516
rect 296168 203396 296220 203448
rect 353300 203396 353352 203448
rect 322940 203328 322992 203380
rect 380164 203328 380216 203380
rect 302884 203260 302936 203312
rect 331220 203260 331272 203312
rect 298008 203192 298060 203244
rect 325148 203192 325200 203244
rect 126060 202852 126112 202904
rect 126612 202852 126664 202904
rect 129004 202920 129056 202972
rect 153384 202852 153436 202904
rect 257712 202852 257764 202904
rect 257988 202852 258040 202904
rect 304080 202895 304132 202904
rect 128912 202784 128964 202836
rect 162124 202784 162176 202836
rect 169116 202784 169168 202836
rect 199108 202784 199160 202836
rect 200028 202784 200080 202836
rect 239680 202784 239732 202836
rect 240140 202784 240192 202836
rect 240508 202784 240560 202836
rect 241428 202784 241480 202836
rect 242992 202784 243044 202836
rect 244096 202784 244148 202836
rect 251824 202784 251876 202836
rect 196900 202716 196952 202768
rect 241520 202716 241572 202768
rect 252376 202716 252428 202768
rect 266728 202784 266780 202836
rect 272248 202784 272300 202836
rect 273168 202784 273220 202836
rect 290556 202784 290608 202836
rect 291016 202784 291068 202836
rect 291384 202784 291436 202836
rect 292304 202784 292356 202836
rect 293132 202784 293184 202836
rect 294604 202784 294656 202836
rect 295800 202784 295852 202836
rect 296444 202784 296496 202836
rect 267832 202716 267884 202768
rect 289268 202716 289320 202768
rect 291844 202716 291896 202768
rect 199844 202648 199896 202700
rect 245200 202648 245252 202700
rect 247500 202648 247552 202700
rect 197636 202580 197688 202632
rect 244740 202580 244792 202632
rect 250904 202580 250956 202632
rect 266636 202648 266688 202700
rect 268292 202580 268344 202632
rect 288808 202580 288860 202632
rect 297916 202784 297968 202836
rect 298744 202784 298796 202836
rect 298928 202784 298980 202836
rect 301504 202784 301556 202836
rect 304080 202861 304089 202895
rect 304089 202861 304123 202895
rect 304123 202861 304132 202895
rect 304080 202852 304132 202861
rect 504180 202895 504232 202904
rect 504180 202861 504189 202895
rect 504189 202861 504223 202895
rect 504223 202861 504232 202895
rect 504180 202852 504232 202861
rect 305644 202784 305696 202836
rect 309140 202784 309192 202836
rect 309600 202784 309652 202836
rect 311900 202784 311952 202836
rect 312544 202784 312596 202836
rect 314844 202784 314896 202836
rect 315580 202784 315632 202836
rect 375748 202784 375800 202836
rect 378784 202784 378836 202836
rect 400588 202784 400640 202836
rect 401508 202784 401560 202836
rect 299112 202716 299164 202768
rect 299204 202648 299256 202700
rect 319260 202716 319312 202768
rect 320088 202716 320140 202768
rect 320548 202716 320600 202768
rect 321468 202716 321520 202768
rect 333152 202716 333204 202768
rect 333888 202716 333940 202768
rect 342076 202716 342128 202768
rect 349988 202716 350040 202768
rect 350448 202716 350500 202768
rect 351000 202716 351052 202768
rect 351828 202716 351880 202768
rect 417148 202716 417200 202768
rect 302976 202648 303028 202700
rect 299664 202580 299716 202632
rect 325700 202648 325752 202700
rect 344008 202648 344060 202700
rect 416872 202648 416924 202700
rect 338764 202580 338816 202632
rect 341432 202580 341484 202632
rect 342168 202580 342220 202632
rect 343088 202580 343140 202632
rect 343548 202580 343600 202632
rect 346676 202580 346728 202632
rect 347596 202580 347648 202632
rect 415400 202580 415452 202632
rect 159364 202512 159416 202564
rect 176936 202512 176988 202564
rect 197544 202512 197596 202564
rect 245660 202512 245712 202564
rect 160744 202444 160796 202496
rect 178040 202444 178092 202496
rect 197360 202444 197412 202496
rect 244924 202444 244976 202496
rect 246028 202444 246080 202496
rect 250076 202444 250128 202496
rect 250996 202444 251048 202496
rect 267740 202512 267792 202564
rect 271420 202512 271472 202564
rect 272524 202512 272576 202564
rect 299388 202512 299440 202564
rect 377220 202512 377272 202564
rect 400956 202512 401008 202564
rect 414664 202512 414716 202564
rect 157984 202376 158036 202428
rect 182180 202376 182232 202428
rect 199200 202376 199252 202428
rect 254032 202376 254084 202428
rect 153844 202308 153896 202360
rect 181260 202308 181312 202360
rect 140044 202240 140096 202292
rect 168380 202240 168432 202292
rect 248972 202308 249024 202360
rect 268384 202444 268436 202496
rect 273996 202444 274048 202496
rect 274548 202444 274600 202496
rect 276940 202444 276992 202496
rect 277308 202444 277360 202496
rect 278688 202444 278740 202496
rect 279424 202444 279476 202496
rect 280988 202444 281040 202496
rect 281356 202444 281408 202496
rect 297732 202444 297784 202496
rect 303896 202444 303948 202496
rect 304908 202444 304960 202496
rect 309140 202444 309192 202496
rect 310612 202444 310664 202496
rect 311256 202444 311308 202496
rect 377496 202444 377548 202496
rect 413192 202444 413244 202496
rect 416044 202444 416096 202496
rect 457444 202444 457496 202496
rect 260196 202376 260248 202428
rect 268476 202376 268528 202428
rect 275284 202376 275336 202428
rect 286416 202376 286468 202428
rect 301872 202376 301924 202428
rect 304080 202376 304132 202428
rect 307024 202376 307076 202428
rect 308404 202376 308456 202428
rect 322940 202376 322992 202428
rect 332508 202376 332560 202428
rect 261668 202308 261720 202360
rect 262128 202308 262180 202360
rect 266820 202308 266872 202360
rect 275744 202308 275796 202360
rect 286324 202308 286376 202360
rect 300124 202308 300176 202360
rect 374460 202308 374512 202360
rect 375288 202308 375340 202360
rect 378968 202308 379020 202360
rect 415768 202376 415820 202428
rect 416596 202376 416648 202428
rect 417516 202376 417568 202428
rect 418068 202376 418120 202428
rect 416780 202308 416832 202360
rect 258172 202240 258224 202292
rect 261944 202240 261996 202292
rect 277308 202240 277360 202292
rect 378140 202240 378192 202292
rect 414940 202240 414992 202292
rect 503904 202308 503956 202360
rect 103428 202172 103480 202224
rect 142528 202172 142580 202224
rect 151084 202172 151136 202224
rect 180340 202172 180392 202224
rect 198832 202172 198884 202224
rect 268568 202172 268620 202224
rect 270960 202172 271012 202224
rect 378324 202172 378376 202224
rect 411076 202172 411128 202224
rect 503812 202240 503864 202292
rect 503720 202172 503772 202224
rect 93768 202104 93820 202156
rect 134708 202104 134760 202156
rect 146944 202104 146996 202156
rect 178684 202104 178736 202156
rect 197912 202104 197964 202156
rect 269488 202104 269540 202156
rect 283564 202104 283616 202156
rect 340144 202104 340196 202156
rect 348332 202104 348384 202156
rect 353576 202104 353628 202156
rect 354588 202104 354640 202156
rect 366180 202104 366232 202156
rect 367008 202104 367060 202156
rect 376484 202104 376536 202156
rect 506480 202104 506532 202156
rect 198924 202036 198976 202088
rect 199936 202036 199988 202088
rect 229100 202036 229152 202088
rect 240968 202036 241020 202088
rect 267372 202036 267424 202088
rect 289544 202036 289596 202088
rect 199752 201968 199804 202020
rect 236644 201968 236696 202020
rect 237288 201968 237340 202020
rect 238668 201968 238720 202020
rect 241060 201968 241112 202020
rect 244648 201968 244700 202020
rect 268016 201968 268068 202020
rect 300768 201968 300820 202020
rect 315304 202036 315356 202088
rect 315948 202036 316000 202088
rect 316040 202036 316092 202088
rect 317144 202036 317196 202088
rect 318616 202036 318668 202088
rect 337384 202036 337436 202088
rect 352748 202036 352800 202088
rect 353208 202036 353260 202088
rect 198648 201900 198700 201952
rect 216036 201900 216088 201952
rect 198740 201832 198792 201884
rect 211712 201832 211764 201884
rect 215944 201832 215996 201884
rect 239220 201900 239272 201952
rect 240048 201900 240100 201952
rect 242072 201900 242124 201952
rect 247684 201900 247736 201952
rect 253112 201900 253164 201952
rect 253756 201900 253808 201952
rect 254860 201900 254912 201952
rect 266912 201900 266964 201952
rect 297824 201900 297876 201952
rect 305644 201968 305696 202020
rect 315396 201968 315448 202020
rect 320640 201968 320692 202020
rect 351736 201968 351788 202020
rect 417240 202036 417292 202088
rect 365352 201968 365404 202020
rect 369124 201968 369176 202020
rect 242164 201832 242216 201884
rect 251916 201832 251968 201884
rect 256148 201832 256200 201884
rect 196808 201764 196860 201816
rect 199292 201696 199344 201748
rect 219532 201696 219584 201748
rect 220820 201764 220872 201816
rect 221280 201764 221332 201816
rect 229100 201764 229152 201816
rect 232412 201764 232464 201816
rect 232504 201764 232556 201816
rect 236736 201764 236788 201816
rect 238116 201764 238168 201816
rect 260840 201764 260892 201816
rect 223028 201696 223080 201748
rect 243176 201696 243228 201748
rect 252468 201696 252520 201748
rect 263600 201696 263652 201748
rect 199568 201628 199620 201680
rect 218612 201628 218664 201680
rect 229744 201628 229796 201680
rect 237380 201628 237432 201680
rect 238024 201628 238076 201680
rect 259460 201628 259512 201680
rect 260104 201628 260156 201680
rect 267464 201832 267516 201884
rect 297548 201832 297600 201884
rect 311164 201900 311216 201952
rect 330484 201900 330536 201952
rect 357900 201900 357952 201952
rect 416964 201900 417016 201952
rect 266268 201764 266320 201816
rect 269120 201764 269172 201816
rect 299572 201764 299624 201816
rect 265164 201696 265216 201748
rect 267188 201696 267240 201748
rect 298376 201696 298428 201748
rect 267096 201628 267148 201680
rect 268200 201628 268252 201680
rect 273628 201628 273680 201680
rect 276664 201628 276716 201680
rect 299480 201628 299532 201680
rect 313648 201832 313700 201884
rect 322756 201832 322808 201884
rect 378232 201832 378284 201884
rect 412272 201832 412324 201884
rect 306472 201696 306524 201748
rect 307300 201696 307352 201748
rect 126428 201560 126480 201612
rect 134156 201560 134208 201612
rect 199660 201560 199712 201612
rect 216864 201560 216916 201612
rect 238208 201560 238260 201612
rect 247776 201560 247828 201612
rect 255228 201560 255280 201612
rect 258724 201560 258776 201612
rect 263876 201560 263928 201612
rect 267004 201560 267056 201612
rect 267740 201560 267792 201612
rect 279240 201560 279292 201612
rect 280068 201560 280120 201612
rect 282644 201560 282696 201612
rect 287704 201560 287756 201612
rect 299296 201560 299348 201612
rect 311992 201764 312044 201816
rect 366916 201764 366968 201816
rect 420184 201764 420236 201816
rect 308404 201696 308456 201748
rect 364892 201696 364944 201748
rect 381544 201696 381596 201748
rect 410156 201696 410208 201748
rect 411168 201696 411220 201748
rect 380072 201628 380124 201680
rect 409236 201628 409288 201680
rect 314936 201560 314988 201612
rect 380256 201560 380308 201612
rect 127624 201492 127676 201544
rect 134340 201492 134392 201544
rect 198556 201492 198608 201544
rect 202880 201492 202932 201544
rect 212448 201492 212500 201544
rect 220084 201492 220136 201544
rect 246488 201492 246540 201544
rect 251456 201492 251508 201544
rect 258080 201424 258132 201476
rect 264888 201492 264940 201544
rect 266544 201492 266596 201544
rect 266636 201492 266688 201544
rect 267280 201492 267332 201544
rect 282276 201492 282328 201544
rect 284944 201492 284996 201544
rect 286232 201492 286284 201544
rect 286968 201492 287020 201544
rect 305000 201492 305052 201544
rect 324044 201492 324096 201544
rect 327080 201492 327132 201544
rect 355324 201492 355376 201544
rect 355968 201492 356020 201544
rect 359648 201492 359700 201544
rect 360108 201492 360160 201544
rect 360568 201492 360620 201544
rect 361396 201492 361448 201544
rect 362316 201492 362368 201544
rect 362776 201492 362828 201544
rect 130568 201220 130620 201272
rect 145564 201220 145616 201272
rect 133512 201152 133564 201204
rect 153384 201152 153436 201204
rect 266452 201152 266504 201204
rect 267648 201152 267700 201204
rect 3884 201084 3936 201136
rect 436560 201084 436612 201136
rect 3608 201016 3660 201068
rect 436468 201016 436520 201068
rect 3424 200948 3476 201000
rect 436376 200948 436428 201000
rect 132408 200880 132460 200932
rect 580264 200880 580316 200932
rect 132224 200812 132276 200864
rect 580448 200812 580500 200864
rect 131396 200744 131448 200796
rect 580356 200744 580408 200796
rect 504180 200404 504232 200456
rect 504456 200404 504508 200456
rect 209872 200200 209924 200252
rect 210286 200200 210338 200252
rect 213920 200200 213972 200252
rect 214610 200200 214662 200252
rect 3240 200132 3292 200184
rect 436652 200132 436704 200184
rect 128544 200064 128596 200116
rect 128912 200064 128964 200116
rect 266452 200064 266504 200116
rect 266728 200064 266780 200116
rect 238760 199860 238812 199912
rect 239496 199860 239548 199912
rect 243084 199860 243136 199912
rect 243820 199860 243872 199912
rect 133604 199792 133656 199844
rect 580264 199792 580316 199844
rect 131396 198296 131448 198348
rect 3424 197344 3476 197396
rect 131396 197344 131448 197396
rect 5356 196256 5408 196308
rect 131396 196256 131448 196308
rect 17224 196052 17276 196104
rect 130476 196052 130528 196104
rect 131764 196095 131816 196104
rect 131764 196061 131773 196095
rect 131773 196061 131807 196095
rect 131807 196061 131816 196095
rect 131764 196052 131816 196061
rect 132868 196095 132920 196104
rect 132868 196061 132877 196095
rect 132877 196061 132911 196095
rect 132911 196061 132920 196095
rect 132868 196052 132920 196061
rect 131396 195984 131448 196036
rect 126428 195916 126480 195968
rect 126612 195916 126664 195968
rect 131764 195959 131816 195968
rect 131764 195925 131773 195959
rect 131773 195925 131807 195959
rect 131807 195925 131816 195959
rect 131764 195916 131816 195925
rect 132868 195959 132920 195968
rect 132868 195925 132877 195959
rect 132877 195925 132911 195959
rect 132911 195925 132920 195959
rect 132868 195916 132920 195925
rect 15844 194556 15896 194608
rect 130476 194556 130528 194608
rect 14464 194420 14516 194472
rect 130476 194420 130528 194472
rect 5264 193128 5316 193180
rect 130384 193128 130436 193180
rect 5448 193060 5500 193112
rect 130476 193060 130528 193112
rect 5172 191768 5224 191820
rect 130476 191768 130528 191820
rect 5080 190408 5132 190460
rect 130476 190408 130528 190460
rect 3516 188980 3568 189032
rect 130384 188980 130436 189032
rect 4988 188912 5040 188964
rect 130476 188912 130528 188964
rect 4896 187620 4948 187672
rect 130476 187620 130528 187672
rect 4804 186260 4856 186312
rect 131212 186260 131264 186312
rect 131212 186124 131264 186176
rect 13084 184832 13136 184884
rect 131212 184832 131264 184884
rect 72424 183472 72476 183524
rect 131212 183472 131264 183524
rect 131212 183336 131264 183388
rect 132868 181432 132920 181484
rect 133328 181432 133380 181484
rect 2872 180752 2924 180804
rect 15844 180752 15896 180804
rect 128912 180795 128964 180804
rect 128912 180761 128921 180795
rect 128921 180761 128955 180795
rect 128955 180761 128964 180795
rect 128912 180752 128964 180761
rect 126428 176604 126480 176656
rect 126612 176604 126664 176656
rect 504456 173884 504508 173936
rect 504640 173884 504692 173936
rect 129004 171096 129056 171148
rect 132960 168580 133012 168632
rect 133328 168580 133380 168632
rect 128912 164228 128964 164280
rect 129004 164228 129056 164280
rect 504180 164160 504232 164212
rect 504364 164160 504416 164212
rect 126520 161440 126572 161492
rect 126612 161440 126664 161492
rect 128912 157428 128964 157480
rect 436836 157360 436888 157412
rect 580172 157360 580224 157412
rect 131212 157335 131264 157344
rect 131212 157301 131221 157335
rect 131221 157301 131255 157335
rect 131255 157301 131264 157335
rect 131212 157292 131264 157301
rect 128820 157224 128872 157276
rect 131120 156272 131172 156324
rect 3516 156068 3568 156120
rect 131304 156068 131356 156120
rect 3240 156000 3292 156052
rect 131120 156000 131172 156052
rect 131304 155932 131356 155984
rect 3608 155864 3660 155916
rect 131120 155864 131172 155916
rect 436100 155184 436152 155236
rect 438124 155184 438176 155236
rect 3332 154232 3384 154284
rect 124220 154368 124272 154420
rect 4068 153144 4120 153196
rect 131120 153144 131172 153196
rect 437388 153144 437440 153196
rect 447784 153144 447836 153196
rect 3976 152940 4028 152992
rect 131304 153119 131356 153128
rect 131304 153085 131313 153119
rect 131313 153085 131347 153119
rect 131347 153085 131356 153119
rect 131304 153076 131356 153085
rect 131212 152872 131264 152924
rect 131304 151895 131356 151904
rect 131304 151861 131313 151895
rect 131313 151861 131347 151895
rect 131347 151861 131356 151895
rect 131304 151852 131356 151861
rect 3792 151716 3844 151768
rect 131120 151716 131172 151768
rect 3700 150356 3752 150408
rect 131120 150356 131172 150408
rect 437388 150356 437440 150408
rect 446404 150356 446456 150408
rect 28264 148996 28316 149048
rect 31024 148928 31076 148980
rect 131120 148928 131172 148980
rect 436100 148996 436152 149048
rect 445024 148996 445076 149048
rect 131120 148588 131172 148640
rect 131212 147679 131264 147688
rect 131212 147645 131221 147679
rect 131221 147645 131255 147679
rect 131255 147645 131264 147679
rect 131212 147636 131264 147645
rect 21364 147568 21416 147620
rect 131120 147568 131172 147620
rect 19984 146208 20036 146260
rect 131120 146208 131172 146260
rect 437388 146140 437440 146192
rect 442264 146140 442316 146192
rect 437020 144848 437072 144900
rect 514024 144848 514076 144900
rect 24768 144644 24820 144696
rect 128176 144712 128228 144764
rect 126244 144372 126296 144424
rect 131120 144372 131172 144424
rect 132868 143556 132920 143608
rect 132776 142171 132828 142180
rect 132776 142137 132785 142171
rect 132785 142137 132819 142171
rect 132819 142137 132828 142171
rect 132776 142128 132828 142137
rect 128820 142103 128872 142112
rect 128820 142069 128829 142103
rect 128829 142069 128863 142103
rect 128863 142069 128872 142103
rect 128820 142060 128872 142069
rect 436100 142060 436152 142112
rect 438216 142060 438268 142112
rect 437388 137912 437440 137964
rect 580540 137912 580592 137964
rect 3332 136552 3384 136604
rect 17224 136552 17276 136604
rect 437020 136552 437072 136604
rect 504456 136552 504508 136604
rect 130660 135532 130712 135584
rect 132316 135532 132368 135584
rect 128820 133875 128872 133884
rect 128820 133841 128829 133875
rect 128829 133841 128863 133875
rect 128863 133841 128872 133875
rect 128820 133832 128872 133841
rect 131120 133832 131172 133884
rect 131304 133832 131356 133884
rect 437388 133832 437440 133884
rect 580632 133832 580684 133884
rect 132316 132404 132368 132456
rect 437388 132404 437440 132456
rect 580724 132404 580776 132456
rect 133144 132336 133196 132388
rect 437388 129684 437440 129736
rect 580816 129684 580868 129736
rect 126060 124108 126112 124160
rect 126428 124108 126480 124160
rect 131120 124108 131172 124160
rect 131396 124108 131448 124160
rect 134064 122383 134116 122392
rect 134064 122349 134073 122383
rect 134073 122349 134107 122383
rect 134107 122349 134116 122383
rect 134064 122340 134116 122349
rect 134064 120776 134116 120828
rect 580908 120776 580960 120828
rect 132408 120708 132460 120760
rect 580356 120708 580408 120760
rect 133972 120640 134024 120692
rect 580264 120640 580316 120692
rect 3332 120572 3384 120624
rect 436284 120572 436336 120624
rect 133144 120300 133196 120352
rect 135168 120300 135220 120352
rect 186596 120232 186648 120284
rect 145012 120139 145064 120148
rect 145012 120105 145021 120139
rect 145021 120105 145055 120139
rect 145055 120105 145064 120139
rect 145012 120096 145064 120105
rect 395114 119756 395166 119808
rect 395988 119756 396040 119808
rect 135168 119348 135220 119400
rect 192116 119348 192168 119400
rect 138296 119280 138348 119332
rect 138848 119280 138900 119332
rect 130752 118940 130804 118992
rect 140780 118940 140832 118992
rect 130936 118872 130988 118924
rect 142252 118872 142304 118924
rect 142528 118872 142580 118924
rect 129556 118804 129608 118856
rect 131028 118736 131080 118788
rect 149060 118736 149112 118788
rect 129648 118668 129700 118720
rect 147772 118668 147824 118720
rect 424784 118668 424836 118720
rect 42708 118600 42760 118652
rect 129740 118600 129792 118652
rect 155316 118600 155368 118652
rect 218428 118600 218480 118652
rect 243544 118600 243596 118652
rect 253296 118600 253348 118652
rect 258264 118600 258316 118652
rect 306012 118600 306064 118652
rect 332876 118600 332928 118652
rect 353116 118600 353168 118652
rect 425336 118600 425388 118652
rect 426348 118600 426400 118652
rect 429844 118600 429896 118652
rect 431776 118600 431828 118652
rect 511264 118600 511316 118652
rect 97908 118532 97960 118584
rect 181076 118532 181128 118584
rect 190368 118532 190420 118584
rect 231308 118532 231360 118584
rect 237196 118532 237248 118584
rect 255320 118532 255372 118584
rect 257344 118532 257396 118584
rect 264336 118532 264388 118584
rect 308496 118532 308548 118584
rect 338396 118532 338448 118584
rect 362316 118532 362368 118584
rect 443000 118532 443052 118584
rect 82728 118464 82780 118516
rect 164516 118464 164568 118516
rect 175924 118464 175976 118516
rect 220268 118464 220320 118516
rect 227720 118464 227772 118516
rect 232504 118464 232556 118516
rect 240232 118464 240284 118516
rect 240968 118464 241020 118516
rect 247776 118464 247828 118516
rect 310888 118464 310940 118516
rect 341432 118464 341484 118516
rect 347596 118464 347648 118516
rect 376024 118464 376076 118516
rect 393596 118464 393648 118516
rect 475384 118464 475436 118516
rect 71504 118396 71556 118448
rect 88340 118396 88392 118448
rect 124128 118396 124180 118448
rect 190460 118396 190512 118448
rect 194508 118396 194560 118448
rect 233240 118396 233292 118448
rect 234528 118396 234580 118448
rect 253940 118396 253992 118448
rect 256608 118396 256660 118448
rect 265532 118396 265584 118448
rect 309692 118396 309744 118448
rect 339592 118396 339644 118448
rect 342168 118396 342220 118448
rect 389824 118396 389876 118448
rect 397276 118396 397328 118448
rect 478144 118396 478196 118448
rect 56508 118328 56560 118380
rect 125784 118328 125836 118380
rect 129280 118328 129332 118380
rect 182916 118328 182968 118380
rect 186044 118328 186096 118380
rect 229468 118328 229520 118380
rect 231768 118328 231820 118380
rect 252744 118328 252796 118380
rect 257988 118328 258040 118380
rect 266360 118328 266412 118380
rect 311532 118328 311584 118380
rect 343916 118328 343968 118380
rect 365996 118328 366048 118380
rect 449900 118328 449952 118380
rect 31668 118260 31720 118312
rect 107568 118260 107620 118312
rect 109040 118260 109092 118312
rect 28908 118192 28960 118244
rect 111708 118192 111760 118244
rect 23388 118124 23440 118176
rect 110328 118124 110380 118176
rect 113088 118260 113140 118312
rect 175648 118260 175700 118312
rect 176016 118260 176068 118312
rect 213828 118260 213880 118312
rect 223672 118260 223724 118312
rect 227628 118260 227680 118312
rect 250260 118260 250312 118312
rect 250536 118260 250588 118312
rect 260840 118260 260892 118312
rect 296168 118260 296220 118312
rect 305644 118260 305696 118312
rect 307208 118260 307260 118312
rect 334624 118260 334676 118312
rect 336648 118260 336700 118312
rect 374644 118260 374696 118312
rect 377036 118260 377088 118312
rect 389916 118260 389968 118312
rect 474004 118260 474056 118312
rect 129188 118192 129240 118244
rect 177396 118192 177448 118244
rect 179328 118192 179380 118244
rect 219992 118192 220044 118244
rect 222200 118192 222252 118244
rect 231124 118192 231176 118244
rect 238024 118192 238076 118244
rect 252100 118192 252152 118244
rect 254676 118192 254728 118244
rect 263692 118192 263744 118244
rect 293776 118192 293828 118244
rect 302884 118192 302936 118244
rect 307668 118192 307720 118244
rect 336924 118192 336976 118244
rect 338488 118192 338540 118244
rect 384212 118192 384264 118244
rect 386236 118192 386288 118244
rect 469864 118192 469916 118244
rect 129096 118124 129148 118176
rect 173900 118124 173952 118176
rect 177304 118124 177356 118176
rect 223948 118124 224000 118176
rect 226248 118124 226300 118176
rect 249800 118124 249852 118176
rect 251088 118124 251140 118176
rect 262496 118124 262548 118176
rect 283932 118124 283984 118176
rect 290096 118124 290148 118176
rect 295616 118124 295668 118176
rect 308404 118124 308456 118176
rect 311716 118124 311768 118176
rect 345204 118124 345256 118176
rect 349436 118124 349488 118176
rect 369676 118124 369728 118176
rect 456800 118124 456852 118176
rect 71688 118056 71740 118108
rect 73804 118056 73856 118108
rect 73988 118056 74040 118108
rect 125692 118056 125744 118108
rect 170036 118056 170088 118108
rect 170404 118056 170456 118108
rect 216680 118056 216732 118108
rect 219256 118056 219308 118108
rect 245936 118056 245988 118108
rect 248328 118056 248380 118108
rect 261300 118056 261352 118108
rect 60648 117988 60700 118040
rect 82728 117988 82780 118040
rect 88340 117988 88392 118040
rect 179420 117988 179472 118040
rect 183468 117988 183520 118040
rect 38476 117920 38528 117972
rect 69664 117920 69716 117972
rect 73988 117920 74040 117972
rect 109040 117920 109092 117972
rect 171876 117920 171928 117972
rect 174544 117920 174596 117972
rect 220084 117988 220136 118040
rect 225788 117988 225840 118040
rect 229008 117988 229060 118040
rect 251272 117988 251324 118040
rect 255228 117988 255280 118040
rect 264980 118056 265032 118108
rect 284576 118056 284628 118108
rect 291384 118056 291436 118108
rect 296628 118056 296680 118108
rect 314844 118056 314896 118108
rect 357992 118056 358044 118108
rect 373356 118056 373408 118108
rect 463700 118056 463752 118108
rect 262128 117988 262180 118040
rect 268016 117988 268068 118040
rect 298652 117988 298704 118040
rect 318984 117988 319036 118040
rect 321928 117988 321980 118040
rect 363512 117988 363564 118040
rect 470600 117988 470652 118040
rect 223488 117920 223540 117972
rect 248512 117920 248564 117972
rect 249708 117920 249760 117972
rect 262220 117920 262272 117972
rect 263508 117920 263560 117972
rect 268660 117920 268712 117972
rect 294328 117920 294380 117972
rect 295248 117920 295300 117972
rect 297456 117920 297508 117972
rect 298008 117920 298060 117972
rect 300492 117920 300544 117972
rect 321744 117920 321796 117972
rect 325424 117920 325476 117972
rect 369124 117920 369176 117972
rect 380716 117920 380768 117972
rect 477500 117920 477552 117972
rect 99196 117852 99248 117904
rect 101220 117852 101272 117904
rect 107568 117852 107620 117904
rect 149888 117852 149940 117904
rect 185676 117852 185728 117904
rect 225144 117852 225196 117904
rect 229192 117852 229244 117904
rect 236184 117852 236236 117904
rect 237288 117852 237340 117904
rect 255780 117852 255832 117904
rect 263416 117852 263468 117904
rect 269212 117852 269264 117904
rect 288900 117852 288952 117904
rect 82728 117784 82780 117836
rect 113088 117784 113140 117836
rect 122748 117784 122800 117836
rect 160836 117784 160888 117836
rect 234712 117784 234764 117836
rect 238668 117784 238720 117836
rect 256700 117784 256752 117836
rect 293132 117852 293184 117904
rect 293868 117852 293920 117904
rect 304816 117852 304868 117904
rect 331312 117852 331364 117904
rect 416780 117852 416832 117904
rect 420828 117852 420880 117904
rect 500224 117852 500276 117904
rect 297364 117784 297416 117836
rect 306656 117784 306708 117836
rect 333980 117784 334032 117836
rect 344008 117784 344060 117836
rect 344928 117784 344980 117836
rect 345848 117784 345900 117836
rect 396724 117784 396776 117836
rect 480904 117784 480956 117836
rect 125784 117716 125836 117768
rect 162860 117716 162912 117768
rect 185584 117716 185636 117768
rect 233884 117716 233936 117768
rect 238852 117716 238904 117768
rect 104992 117648 105044 117700
rect 115204 117648 115256 117700
rect 129372 117648 129424 117700
rect 135260 117648 135312 117700
rect 166356 117648 166408 117700
rect 175280 117648 175332 117700
rect 175464 117648 175516 117700
rect 195980 117648 196032 117700
rect 197268 117648 197320 117700
rect 128820 117580 128872 117632
rect 158996 117580 159048 117632
rect 195888 117580 195940 117632
rect 120724 117512 120776 117564
rect 125692 117512 125744 117564
rect 130384 117512 130436 117564
rect 130844 117512 130896 117564
rect 135260 117512 135312 117564
rect 135444 117512 135496 117564
rect 142988 117512 143040 117564
rect 122104 117444 122156 117496
rect 122748 117444 122800 117496
rect 123484 117444 123536 117496
rect 124128 117444 124180 117496
rect 130568 117444 130620 117496
rect 143724 117512 143776 117564
rect 157340 117512 157392 117564
rect 193864 117512 193916 117564
rect 233148 117648 233200 117700
rect 245476 117716 245528 117768
rect 259460 117716 259512 117768
rect 302148 117716 302200 117768
rect 329288 117716 329340 117768
rect 358176 117716 358228 117768
rect 364064 117716 364116 117768
rect 400864 117716 400916 117768
rect 415308 117716 415360 117768
rect 418160 117716 418212 117768
rect 429660 117716 429712 117768
rect 430488 117716 430540 117768
rect 430948 117716 431000 117768
rect 431868 117716 431920 117768
rect 502984 117716 503036 117768
rect 240048 117648 240100 117700
rect 256976 117648 257028 117700
rect 261484 117648 261536 117700
rect 267740 117648 267792 117700
rect 304172 117648 304224 117700
rect 329840 117648 329892 117700
rect 360476 117648 360528 117700
rect 398104 117648 398156 117700
rect 411904 117648 411956 117700
rect 417424 117648 417476 117700
rect 234988 117580 235040 117632
rect 201408 117512 201460 117564
rect 236828 117580 236880 117632
rect 236644 117512 236696 117564
rect 242256 117580 242308 117632
rect 244188 117580 244240 117632
rect 258816 117580 258868 117632
rect 294972 117580 295024 117632
rect 311900 117580 311952 117632
rect 314568 117580 314620 117632
rect 320824 117580 320876 117632
rect 330484 117580 330536 117632
rect 331036 117580 331088 117632
rect 356796 117580 356848 117632
rect 208308 117444 208360 117496
rect 67548 117376 67600 117428
rect 71044 117376 71096 117428
rect 168380 117376 168432 117428
rect 211068 117376 211120 117428
rect 225604 117376 225656 117428
rect 97264 117308 97316 117360
rect 97908 117308 97960 117360
rect 111708 117308 111760 117360
rect 148048 117308 148100 117360
rect 171784 117308 171836 117360
rect 212908 117308 212960 117360
rect 214564 117308 214616 117360
rect 226984 117308 227036 117360
rect 230388 117444 230440 117496
rect 238024 117444 238076 117496
rect 240416 117376 240468 117428
rect 241428 117512 241480 117564
rect 257620 117512 257672 117564
rect 266268 117512 266320 117564
rect 270500 117512 270552 117564
rect 280068 117512 280120 117564
rect 283012 117512 283064 117564
rect 299848 117512 299900 117564
rect 315304 117512 315356 117564
rect 354956 117512 355008 117564
rect 369216 117512 369268 117564
rect 241704 117444 241756 117496
rect 243544 117376 243596 117428
rect 245568 117444 245620 117496
rect 260012 117444 260064 117496
rect 267648 117444 267700 117496
rect 271052 117444 271104 117496
rect 282736 117444 282788 117496
rect 284944 117444 284996 117496
rect 320088 117444 320140 117496
rect 324964 117444 325016 117496
rect 326344 117444 326396 117496
rect 328092 117444 328144 117496
rect 328276 117444 328328 117496
rect 367836 117444 367888 117496
rect 377404 117444 377456 117496
rect 391112 117580 391164 117632
rect 391756 117580 391808 117632
rect 404268 117580 404320 117632
rect 384396 117512 384448 117564
rect 413284 117512 413336 117564
rect 393964 117444 394016 117496
rect 399668 117444 399720 117496
rect 400036 117444 400088 117496
rect 419264 117512 419316 117564
rect 420184 117512 420236 117564
rect 422944 117648 422996 117700
rect 424324 117648 424376 117700
rect 427728 117648 427780 117700
rect 493324 117648 493376 117700
rect 482284 117580 482336 117632
rect 413744 117444 413796 117496
rect 416044 117444 416096 117496
rect 418620 117444 418672 117496
rect 419448 117444 419500 117496
rect 419908 117444 419960 117496
rect 420828 117444 420880 117496
rect 421748 117444 421800 117496
rect 422208 117444 422260 117496
rect 496084 117512 496136 117564
rect 424140 117444 424192 117496
rect 424968 117444 425020 117496
rect 425428 117444 425480 117496
rect 426348 117444 426400 117496
rect 427268 117444 427320 117496
rect 427728 117444 427780 117496
rect 428464 117444 428516 117496
rect 430304 117444 430356 117496
rect 431224 117444 431276 117496
rect 432788 117444 432840 117496
rect 433248 117444 433300 117496
rect 507124 117444 507176 117496
rect 239404 117308 239456 117360
rect 244280 117308 244332 117360
rect 247224 117376 247276 117428
rect 247684 117376 247736 117428
rect 251456 117376 251508 117428
rect 252468 117376 252520 117428
rect 263140 117376 263192 117428
rect 269764 117376 269816 117428
rect 271880 117376 271932 117428
rect 272524 117376 272576 117428
rect 273536 117376 273588 117428
rect 278412 117376 278464 117428
rect 279148 117376 279200 117428
rect 282092 117376 282144 117428
rect 283564 117376 283616 117428
rect 289452 117376 289504 117428
rect 294604 117376 294656 117428
rect 318248 117376 318300 117428
rect 322204 117376 322256 117428
rect 332968 117376 333020 117428
rect 333888 117376 333940 117428
rect 371516 117376 371568 117428
rect 372528 117376 372580 117428
rect 405188 117376 405240 117428
rect 405648 117376 405700 117428
rect 408224 117376 408276 117428
rect 486424 117376 486476 117428
rect 250444 117308 250496 117360
rect 254584 117308 254636 117360
rect 259368 117308 259420 117360
rect 266820 117308 266872 117360
rect 268384 117308 268436 117360
rect 269856 117308 269908 117360
rect 273168 117308 273220 117360
rect 274180 117308 274232 117360
rect 277860 117308 277912 117360
rect 278872 117308 278924 117360
rect 279056 117308 279108 117360
rect 280344 117308 280396 117360
rect 280896 117308 280948 117360
rect 281356 117308 281408 117360
rect 283380 117308 283432 117360
rect 284208 117308 284260 117360
rect 285220 117308 285272 117360
rect 285588 117308 285640 117360
rect 286416 117308 286468 117360
rect 286968 117308 287020 117360
rect 287612 117308 287664 117360
rect 288348 117308 288400 117360
rect 290004 117308 290056 117360
rect 291108 117308 291160 117360
rect 291936 117308 291988 117360
rect 292488 117308 292540 117360
rect 301136 117308 301188 117360
rect 302148 117308 302200 117360
rect 302976 117308 303028 117360
rect 303528 117308 303580 117360
rect 305368 117308 305420 117360
rect 306288 117308 306340 117360
rect 312728 117308 312780 117360
rect 313188 117308 313240 117360
rect 313924 117308 313976 117360
rect 314568 117308 314620 117360
rect 315212 117308 315264 117360
rect 315856 117308 315908 117360
rect 316408 117308 316460 117360
rect 317328 117308 317380 117360
rect 319444 117308 319496 117360
rect 320088 117308 320140 117360
rect 320732 117308 320784 117360
rect 321376 117308 321428 117360
rect 323768 117308 323820 117360
rect 324228 117308 324280 117360
rect 326252 117308 326304 117360
rect 326988 117308 327040 117360
rect 327448 117308 327500 117360
rect 328368 117308 328420 117360
rect 331680 117308 331732 117360
rect 332508 117308 332560 117360
rect 333520 117308 333572 117360
rect 333796 117308 333848 117360
rect 334808 117308 334860 117360
rect 335268 117308 335320 117360
rect 336004 117308 336056 117360
rect 336648 117308 336700 117360
rect 337200 117308 337252 117360
rect 338028 117308 338080 117360
rect 339040 117308 339092 117360
rect 339408 117308 339460 117360
rect 340328 117308 340380 117360
rect 340788 117308 340840 117360
rect 341524 117308 341576 117360
rect 342168 117308 342220 117360
rect 342720 117308 342772 117360
rect 343548 117308 343600 117360
rect 344560 117308 344612 117360
rect 344836 117308 344888 117360
rect 347044 117308 347096 117360
rect 347688 117308 347740 117360
rect 348240 117308 348292 117360
rect 349068 117308 349120 117360
rect 350080 117308 350132 117360
rect 350448 117308 350500 117360
rect 351276 117308 351328 117360
rect 351828 117308 351880 117360
rect 352564 117308 352616 117360
rect 353208 117308 353260 117360
rect 353760 117308 353812 117360
rect 354588 117308 354640 117360
rect 355600 117308 355652 117360
rect 355968 117308 356020 117360
rect 358084 117308 358136 117360
rect 358636 117308 358688 117360
rect 359280 117308 359332 117360
rect 360108 117308 360160 117360
rect 361120 117308 361172 117360
rect 361488 117308 361540 117360
rect 363604 117308 363656 117360
rect 364248 117308 364300 117360
rect 364800 117308 364852 117360
rect 365628 117308 365680 117360
rect 366640 117308 366692 117360
rect 367008 117308 367060 117360
rect 369032 117308 369084 117360
rect 369768 117308 369820 117360
rect 370320 117308 370372 117360
rect 371148 117308 371200 117360
rect 372160 117308 372212 117360
rect 372436 117308 372488 117360
rect 374552 117308 374604 117360
rect 375196 117308 375248 117360
rect 375840 117308 375892 117360
rect 376668 117308 376720 117360
rect 377680 117308 377732 117360
rect 378048 117308 378100 117360
rect 378876 117308 378928 117360
rect 379428 117308 379480 117360
rect 380072 117308 380124 117360
rect 380808 117308 380860 117360
rect 381360 117308 381412 117360
rect 382188 117308 382240 117360
rect 382556 117308 382608 117360
rect 383568 117308 383620 117360
rect 385592 117308 385644 117360
rect 386328 117308 386380 117360
rect 386788 117308 386840 117360
rect 387616 117308 387668 117360
rect 388076 117308 388128 117360
rect 389088 117308 389140 117360
rect 392308 117308 392360 117360
rect 393136 117308 393188 117360
rect 396632 117308 396684 117360
rect 397368 117308 397420 117360
rect 397828 117308 397880 117360
rect 398748 117308 398800 117360
rect 399116 117308 399168 117360
rect 400128 117308 400180 117360
rect 402152 117308 402204 117360
rect 402796 117308 402848 117360
rect 403348 117308 403400 117360
rect 404268 117308 404320 117360
rect 406384 117308 406436 117360
rect 407028 117308 407080 117360
rect 407672 117308 407724 117360
rect 408408 117308 408460 117360
rect 408868 117308 408920 117360
rect 409696 117308 409748 117360
rect 410708 117308 410760 117360
rect 411168 117308 411220 117360
rect 413192 117308 413244 117360
rect 413928 117308 413980 117360
rect 414388 117308 414440 117360
rect 415308 117308 415360 117360
rect 416228 117308 416280 117360
rect 416688 117308 416740 117360
rect 489184 117308 489236 117360
rect 122840 117240 122892 117292
rect 133788 117240 133840 117292
rect 402244 117240 402296 117292
rect 198740 116560 198792 116612
rect 199476 116560 199528 116612
rect 200120 116560 200172 116612
rect 200672 116560 200724 116612
rect 201500 116560 201552 116612
rect 201868 116560 201920 116612
rect 202972 116560 203024 116612
rect 203708 116560 203760 116612
rect 204260 116560 204312 116612
rect 204904 116560 204956 116612
rect 190736 115948 190788 116000
rect 191012 115948 191064 116000
rect 272248 115948 272300 116000
rect 272432 115948 272484 116000
rect 322388 115948 322440 116000
rect 322572 115948 322624 116000
rect 382924 115948 382976 116000
rect 383108 115948 383160 116000
rect 133788 115880 133840 115932
rect 134524 115880 134576 115932
rect 150808 115880 150860 115932
rect 151360 115880 151412 115932
rect 173992 115880 174044 115932
rect 174360 115880 174412 115932
rect 248328 115880 248380 115932
rect 248420 115880 248472 115932
rect 276020 115880 276072 115932
rect 276112 115880 276164 115932
rect 301688 115880 301740 115932
rect 301964 115880 302016 115932
rect 388720 115880 388772 115932
rect 388904 115880 388956 115932
rect 404084 115880 404136 115932
rect 414848 115880 414900 115932
rect 414940 115880 414992 115932
rect 420552 115923 420604 115932
rect 420552 115889 420561 115923
rect 420561 115889 420595 115923
rect 420595 115889 420604 115923
rect 420552 115880 420604 115889
rect 426072 115880 426124 115932
rect 426256 115880 426308 115932
rect 431500 115923 431552 115932
rect 431500 115889 431509 115923
rect 431509 115889 431543 115923
rect 431543 115889 431552 115923
rect 431500 115880 431552 115889
rect 202880 114520 202932 114572
rect 203156 114520 203208 114572
rect 215392 114520 215444 114572
rect 215944 114520 215996 114572
rect 232228 114520 232280 114572
rect 232596 114520 232648 114572
rect 325700 114563 325752 114572
rect 325700 114529 325709 114563
rect 325709 114529 325743 114563
rect 325743 114529 325752 114563
rect 325700 114520 325752 114529
rect 174360 114452 174412 114504
rect 230388 114495 230440 114504
rect 230388 114461 230397 114495
rect 230397 114461 230431 114495
rect 230431 114461 230440 114495
rect 230388 114452 230440 114461
rect 248420 114452 248472 114504
rect 135260 113840 135312 113892
rect 135720 113840 135772 113892
rect 139400 113840 139452 113892
rect 140044 113840 140096 113892
rect 151820 113840 151872 113892
rect 152280 113840 152332 113892
rect 153200 113840 153252 113892
rect 154120 113840 154172 113892
rect 155960 113840 156012 113892
rect 156604 113840 156656 113892
rect 167000 113840 167052 113892
rect 167644 113840 167696 113892
rect 169852 113840 169904 113892
rect 170680 113840 170732 113892
rect 172520 113840 172572 113892
rect 173072 113840 173124 113892
rect 175372 113840 175424 113892
rect 176200 113840 176252 113892
rect 178040 113840 178092 113892
rect 178592 113840 178644 113892
rect 186412 113840 186464 113892
rect 186596 113840 186648 113892
rect 191932 113840 191984 113892
rect 192668 113840 192720 113892
rect 194692 113840 194744 113892
rect 195152 113840 195204 113892
rect 205640 113840 205692 113892
rect 206192 113840 206244 113892
rect 208492 113840 208544 113892
rect 209228 113840 209280 113892
rect 209872 113840 209924 113892
rect 210424 113840 210476 113892
rect 211160 113840 211212 113892
rect 211712 113840 211764 113892
rect 219532 113840 219584 113892
rect 219716 113840 219768 113892
rect 229192 113840 229244 113892
rect 230020 113840 230072 113892
rect 223672 113092 223724 113144
rect 224500 113092 224552 113144
rect 229192 113092 229244 113144
rect 136732 112480 136784 112532
rect 137560 112480 137612 112532
rect 140780 111868 140832 111920
rect 141240 111868 141292 111920
rect 436928 111732 436980 111784
rect 579804 111732 579856 111784
rect 189080 111528 189132 111580
rect 189632 111528 189684 111580
rect 244464 109080 244516 109132
rect 143632 109012 143684 109064
rect 144184 109012 144236 109064
rect 192024 109012 192076 109064
rect 387524 109012 387576 109064
rect 387708 109012 387760 109064
rect 393044 109012 393096 109064
rect 393228 109012 393280 109064
rect 192208 108944 192260 108996
rect 244464 108944 244516 108996
rect 420552 108987 420604 108996
rect 420552 108953 420561 108987
rect 420561 108953 420595 108987
rect 420595 108953 420604 108987
rect 420552 108944 420604 108953
rect 431684 108944 431736 108996
rect 186136 106292 186188 106344
rect 403900 106335 403952 106344
rect 403900 106301 403909 106335
rect 403909 106301 403943 106335
rect 403943 106301 403952 106335
rect 403900 106292 403952 106301
rect 128912 106267 128964 106276
rect 128912 106233 128921 106267
rect 128921 106233 128955 106267
rect 128955 106233 128964 106267
rect 128912 106224 128964 106233
rect 133972 106224 134024 106276
rect 157524 106267 157576 106276
rect 157524 106233 157533 106267
rect 157533 106233 157567 106267
rect 157567 106233 157576 106267
rect 157524 106224 157576 106233
rect 179512 106267 179564 106276
rect 179512 106233 179521 106267
rect 179521 106233 179555 106267
rect 179555 106233 179564 106267
rect 179512 106224 179564 106233
rect 221004 106267 221056 106276
rect 221004 106233 221013 106267
rect 221013 106233 221047 106267
rect 221047 106233 221056 106267
rect 221004 106224 221056 106233
rect 244464 106224 244516 106276
rect 244556 106224 244608 106276
rect 301964 106267 302016 106276
rect 301964 106233 301973 106267
rect 301973 106233 302007 106267
rect 302007 106233 302016 106267
rect 301964 106224 302016 106233
rect 322664 106267 322716 106276
rect 322664 106233 322673 106267
rect 322673 106233 322707 106267
rect 322707 106233 322716 106267
rect 322664 106224 322716 106233
rect 388720 106224 388772 106276
rect 388812 106224 388864 106276
rect 394424 106267 394476 106276
rect 394424 106233 394433 106267
rect 394433 106233 394467 106267
rect 394467 106233 394476 106267
rect 394424 106224 394476 106233
rect 420552 106224 420604 106276
rect 420644 106224 420696 106276
rect 431592 106224 431644 106276
rect 431684 106224 431736 106276
rect 186228 106156 186280 106208
rect 133972 106088 134024 106140
rect 227904 104932 227956 104984
rect 174176 104907 174228 104916
rect 174176 104873 174185 104907
rect 174185 104873 174219 104907
rect 174219 104873 174228 104907
rect 174176 104864 174228 104873
rect 227812 104864 227864 104916
rect 248328 104907 248380 104916
rect 248328 104873 248337 104907
rect 248337 104873 248371 104907
rect 248371 104873 248380 104907
rect 248328 104864 248380 104873
rect 215392 104839 215444 104848
rect 215392 104805 215401 104839
rect 215401 104805 215435 104839
rect 215435 104805 215444 104839
rect 215392 104796 215444 104805
rect 276112 104839 276164 104848
rect 276112 104805 276121 104839
rect 276121 104805 276155 104839
rect 276155 104805 276164 104839
rect 276112 104796 276164 104805
rect 325700 104839 325752 104848
rect 325700 104805 325709 104839
rect 325709 104805 325743 104839
rect 325743 104805 325752 104839
rect 325700 104796 325752 104805
rect 415032 104839 415084 104848
rect 415032 104805 415041 104839
rect 415041 104805 415075 104839
rect 415075 104805 415084 104839
rect 415032 104796 415084 104805
rect 426256 104839 426308 104848
rect 426256 104805 426265 104839
rect 426265 104805 426299 104839
rect 426299 104805 426308 104839
rect 426256 104796 426308 104805
rect 431592 104839 431644 104848
rect 431592 104805 431601 104839
rect 431601 104805 431635 104839
rect 431635 104805 431644 104839
rect 431592 104796 431644 104805
rect 229192 103504 229244 103556
rect 230388 103547 230440 103556
rect 230388 103513 230397 103547
rect 230397 103513 230431 103547
rect 230431 103513 230440 103547
rect 230388 103504 230440 103513
rect 186228 103479 186280 103488
rect 186228 103445 186237 103479
rect 186237 103445 186271 103479
rect 186271 103445 186280 103479
rect 186228 103436 186280 103445
rect 233332 103479 233384 103488
rect 233332 103445 233341 103479
rect 233341 103445 233375 103479
rect 233375 103445 233384 103479
rect 233332 103436 233384 103445
rect 279792 103436 279844 103488
rect 223672 102119 223724 102128
rect 223672 102085 223681 102119
rect 223681 102085 223715 102119
rect 223715 102085 223724 102119
rect 223672 102076 223724 102085
rect 161388 101396 161440 101448
rect 161756 101396 161808 101448
rect 222292 100691 222344 100700
rect 222292 100657 222301 100691
rect 222301 100657 222335 100691
rect 222335 100657 222344 100691
rect 222292 100648 222344 100657
rect 240232 100079 240284 100088
rect 240232 100045 240241 100079
rect 240241 100045 240275 100079
rect 240275 100045 240284 100079
rect 240232 100036 240284 100045
rect 248420 100036 248472 100088
rect 140964 99424 141016 99476
rect 208768 99424 208820 99476
rect 214196 99424 214248 99476
rect 232228 99424 232280 99476
rect 140872 99356 140924 99408
rect 208584 99356 208636 99408
rect 214104 99356 214156 99408
rect 227812 99356 227864 99408
rect 232136 99356 232188 99408
rect 248512 99356 248564 99408
rect 128912 99331 128964 99340
rect 128912 99297 128921 99331
rect 128921 99297 128955 99331
rect 128955 99297 128964 99331
rect 128912 99288 128964 99297
rect 157616 99288 157668 99340
rect 179512 99331 179564 99340
rect 179512 99297 179521 99331
rect 179521 99297 179555 99331
rect 179555 99297 179564 99331
rect 179512 99288 179564 99297
rect 227904 99288 227956 99340
rect 248420 99288 248472 99340
rect 383292 99424 383344 99476
rect 403900 99356 403952 99408
rect 301964 99331 302016 99340
rect 301964 99297 301973 99331
rect 301973 99297 302007 99331
rect 302007 99297 302016 99331
rect 301964 99288 302016 99297
rect 322664 99331 322716 99340
rect 322664 99297 322673 99331
rect 322673 99297 322707 99331
rect 322707 99297 322716 99331
rect 322664 99288 322716 99297
rect 383200 99288 383252 99340
rect 394424 99331 394476 99340
rect 394424 99297 394433 99331
rect 394433 99297 394467 99331
rect 394467 99297 394476 99331
rect 394424 99288 394476 99297
rect 403992 99288 404044 99340
rect 174176 97180 174228 97232
rect 145012 96679 145064 96688
rect 145012 96645 145021 96679
rect 145021 96645 145055 96679
rect 145055 96645 145064 96679
rect 145012 96636 145064 96645
rect 162952 96636 163004 96688
rect 221004 96679 221056 96688
rect 221004 96645 221013 96679
rect 221013 96645 221047 96679
rect 221047 96645 221056 96679
rect 221004 96636 221056 96645
rect 128912 96568 128964 96620
rect 129004 96568 129056 96620
rect 138020 96611 138072 96620
rect 138020 96577 138029 96611
rect 138029 96577 138063 96611
rect 138063 96577 138072 96611
rect 138020 96568 138072 96577
rect 162860 96568 162912 96620
rect 214104 96568 214156 96620
rect 214288 96568 214340 96620
rect 216772 96611 216824 96620
rect 216772 96577 216781 96611
rect 216781 96577 216815 96611
rect 216815 96577 216824 96611
rect 216772 96568 216824 96577
rect 290556 96611 290608 96620
rect 290556 96577 290565 96611
rect 290565 96577 290599 96611
rect 290599 96577 290608 96611
rect 290556 96568 290608 96577
rect 341064 96568 341116 96620
rect 341340 96568 341392 96620
rect 383200 96568 383252 96620
rect 388720 96568 388772 96620
rect 403992 96568 404044 96620
rect 420736 96568 420788 96620
rect 150624 95344 150676 95396
rect 150808 95344 150860 95396
rect 426256 95319 426308 95328
rect 426256 95285 426265 95319
rect 426265 95285 426299 95319
rect 426299 95285 426308 95319
rect 426256 95276 426308 95285
rect 173900 95251 173952 95260
rect 173900 95217 173909 95251
rect 173909 95217 173943 95251
rect 173943 95217 173952 95251
rect 173900 95208 173952 95217
rect 215392 95251 215444 95260
rect 215392 95217 215401 95251
rect 215401 95217 215435 95251
rect 215435 95217 215444 95251
rect 215392 95208 215444 95217
rect 240324 95208 240376 95260
rect 248328 95251 248380 95260
rect 248328 95217 248337 95251
rect 248337 95217 248371 95251
rect 248371 95217 248380 95251
rect 248328 95208 248380 95217
rect 276112 95251 276164 95260
rect 276112 95217 276121 95251
rect 276121 95217 276155 95251
rect 276155 95217 276164 95251
rect 276112 95208 276164 95217
rect 325700 95251 325752 95260
rect 325700 95217 325709 95251
rect 325709 95217 325743 95251
rect 325743 95217 325752 95251
rect 325700 95208 325752 95217
rect 415216 95208 415268 95260
rect 140872 95183 140924 95192
rect 140872 95149 140881 95183
rect 140881 95149 140915 95183
rect 140915 95149 140924 95183
rect 140872 95140 140924 95149
rect 150624 95183 150676 95192
rect 150624 95149 150633 95183
rect 150633 95149 150667 95183
rect 150667 95149 150676 95183
rect 150624 95140 150676 95149
rect 162860 95183 162912 95192
rect 162860 95149 162869 95183
rect 162869 95149 162903 95183
rect 162903 95149 162912 95183
rect 271972 95183 272024 95192
rect 162860 95140 162912 95149
rect 271972 95149 271981 95183
rect 271981 95149 272015 95183
rect 272015 95149 272024 95183
rect 271972 95140 272024 95149
rect 229192 93916 229244 93968
rect 186320 93848 186372 93900
rect 229284 93848 229336 93900
rect 233424 93848 233476 93900
rect 279700 93891 279752 93900
rect 279700 93857 279709 93891
rect 279709 93857 279743 93891
rect 279743 93857 279752 93891
rect 279700 93848 279752 93857
rect 2780 93304 2832 93356
rect 5356 93304 5408 93356
rect 161388 92964 161440 93016
rect 161664 92964 161716 93016
rect 223764 92488 223816 92540
rect 227904 92463 227956 92472
rect 227904 92429 227913 92463
rect 227913 92429 227947 92463
rect 227947 92429 227956 92463
rect 227904 92420 227956 92429
rect 207204 89768 207256 89820
rect 126060 89700 126112 89752
rect 126244 89700 126296 89752
rect 179420 89700 179472 89752
rect 179604 89700 179656 89752
rect 183652 89700 183704 89752
rect 190644 89700 190696 89752
rect 192300 89700 192352 89752
rect 138112 89632 138164 89684
rect 183744 89564 183796 89616
rect 190736 89564 190788 89616
rect 322572 89700 322624 89752
rect 322756 89700 322808 89752
rect 394332 89700 394384 89752
rect 394516 89700 394568 89752
rect 415216 89768 415268 89820
rect 207204 89632 207256 89684
rect 415124 89632 415176 89684
rect 192392 89564 192444 89616
rect 234804 89564 234856 89616
rect 216864 89496 216916 89548
rect 234804 89428 234856 89480
rect 290556 89403 290608 89412
rect 290556 89369 290565 89403
rect 290565 89369 290599 89403
rect 290599 89369 290608 89403
rect 290556 89360 290608 89369
rect 131212 88272 131264 88324
rect 580172 88272 580224 88324
rect 248604 86980 248656 87032
rect 383108 87023 383160 87032
rect 383108 86989 383117 87023
rect 383117 86989 383151 87023
rect 383151 86989 383160 87023
rect 383108 86980 383160 86989
rect 388628 87023 388680 87032
rect 388628 86989 388637 87023
rect 388637 86989 388671 87023
rect 388671 86989 388680 87023
rect 388628 86980 388680 86989
rect 403900 87023 403952 87032
rect 403900 86989 403909 87023
rect 403909 86989 403943 87023
rect 403943 86989 403952 87023
rect 403900 86980 403952 86989
rect 420644 87023 420696 87032
rect 420644 86989 420653 87023
rect 420653 86989 420687 87023
rect 420687 86989 420696 87023
rect 420644 86980 420696 86989
rect 426256 86980 426308 87032
rect 431592 87023 431644 87032
rect 431592 86989 431601 87023
rect 431601 86989 431635 87023
rect 431635 86989 431644 87023
rect 431592 86980 431644 86989
rect 128728 86912 128780 86964
rect 128912 86912 128964 86964
rect 140964 86844 141016 86896
rect 162952 86844 163004 86896
rect 290556 86955 290608 86964
rect 290556 86921 290565 86955
rect 290565 86921 290599 86955
rect 290599 86921 290608 86955
rect 290556 86912 290608 86921
rect 322664 86955 322716 86964
rect 322664 86921 322673 86955
rect 322673 86921 322707 86955
rect 322707 86921 322716 86955
rect 322664 86912 322716 86921
rect 394424 86955 394476 86964
rect 394424 86921 394433 86955
rect 394433 86921 394467 86955
rect 394467 86921 394476 86955
rect 394424 86912 394476 86921
rect 248788 86844 248840 86896
rect 150716 85552 150768 85604
rect 233332 85552 233384 85604
rect 233516 85552 233568 85604
rect 272064 85552 272116 85604
rect 426164 85595 426216 85604
rect 426164 85561 426173 85595
rect 426173 85561 426207 85595
rect 426207 85561 426216 85595
rect 426164 85552 426216 85561
rect 128728 85484 128780 85536
rect 148140 85484 148192 85536
rect 161664 85484 161716 85536
rect 161756 85484 161808 85536
rect 214104 85527 214156 85536
rect 214104 85493 214113 85527
rect 214113 85493 214147 85527
rect 214147 85493 214156 85527
rect 214104 85484 214156 85493
rect 325700 85527 325752 85536
rect 325700 85493 325709 85527
rect 325709 85493 325743 85527
rect 325743 85493 325752 85527
rect 325700 85484 325752 85493
rect 140964 84167 141016 84176
rect 140964 84133 140973 84167
rect 140973 84133 141007 84167
rect 141007 84133 141016 84167
rect 140964 84124 141016 84133
rect 192392 84124 192444 84176
rect 230388 84167 230440 84176
rect 230388 84133 230397 84167
rect 230397 84133 230431 84167
rect 230431 84133 230440 84167
rect 230388 84124 230440 84133
rect 248788 84124 248840 84176
rect 279700 84167 279752 84176
rect 279700 84133 279709 84167
rect 279709 84133 279743 84167
rect 279743 84133 279752 84167
rect 279700 84124 279752 84133
rect 426164 84124 426216 84176
rect 222568 82832 222620 82884
rect 228088 82832 228140 82884
rect 420276 82084 420328 82136
rect 420644 82084 420696 82136
rect 207296 80835 207348 80844
rect 207296 80801 207305 80835
rect 207305 80801 207339 80835
rect 207339 80801 207348 80835
rect 207296 80792 207348 80801
rect 271880 80724 271932 80776
rect 272156 80724 272208 80776
rect 216864 80155 216916 80164
rect 216864 80121 216873 80155
rect 216873 80121 216907 80155
rect 216907 80121 216916 80155
rect 216864 80112 216916 80121
rect 223764 80112 223816 80164
rect 229284 80112 229336 80164
rect 232136 80155 232188 80164
rect 232136 80121 232145 80155
rect 232145 80121 232179 80155
rect 232179 80121 232188 80155
rect 232136 80112 232188 80121
rect 234804 80112 234856 80164
rect 240324 80112 240376 80164
rect 150532 80044 150584 80096
rect 150716 80044 150768 80096
rect 234712 80044 234764 80096
rect 240232 80044 240284 80096
rect 431592 80044 431644 80096
rect 431776 80044 431828 80096
rect 3240 79976 3292 80028
rect 434996 79976 435048 80028
rect 216864 79951 216916 79960
rect 216864 79917 216873 79951
rect 216873 79917 216907 79951
rect 216907 79917 216916 79951
rect 216864 79908 216916 79917
rect 232136 79951 232188 79960
rect 232136 79917 232145 79951
rect 232145 79917 232179 79951
rect 232179 79917 232188 79951
rect 232136 79908 232188 79917
rect 290556 79951 290608 79960
rect 290556 79917 290565 79951
rect 290565 79917 290599 79951
rect 290599 79917 290608 79951
rect 290556 79908 290608 79917
rect 301872 77324 301924 77376
rect 302056 77324 302108 77376
rect 126244 77256 126296 77308
rect 126336 77256 126388 77308
rect 207296 77299 207348 77308
rect 207296 77265 207305 77299
rect 207305 77265 207339 77299
rect 207339 77265 207348 77299
rect 207296 77256 207348 77265
rect 245752 77256 245804 77308
rect 245936 77256 245988 77308
rect 322756 77256 322808 77308
rect 394516 77256 394568 77308
rect 132132 77188 132184 77240
rect 580172 77188 580224 77240
rect 302056 77120 302108 77172
rect 341340 77163 341392 77172
rect 341340 77129 341349 77163
rect 341349 77129 341383 77163
rect 341383 77129 341392 77163
rect 341340 77120 341392 77129
rect 383200 77163 383252 77172
rect 383200 77129 383209 77163
rect 383209 77129 383243 77163
rect 383243 77129 383252 77163
rect 383200 77120 383252 77129
rect 388720 77163 388772 77172
rect 388720 77129 388729 77163
rect 388729 77129 388763 77163
rect 388763 77129 388772 77163
rect 388720 77120 388772 77129
rect 403992 77163 404044 77172
rect 403992 77129 404001 77163
rect 404001 77129 404035 77163
rect 404035 77129 404044 77163
rect 403992 77120 404044 77129
rect 128636 75939 128688 75948
rect 128636 75905 128645 75939
rect 128645 75905 128679 75939
rect 128679 75905 128688 75939
rect 128636 75896 128688 75905
rect 147956 75939 148008 75948
rect 147956 75905 147965 75939
rect 147965 75905 147999 75939
rect 147999 75905 148008 75939
rect 147956 75896 148008 75905
rect 157340 75896 157392 75948
rect 157708 75896 157760 75948
rect 183744 75896 183796 75948
rect 183836 75896 183888 75948
rect 186228 75896 186280 75948
rect 186320 75896 186372 75948
rect 190552 75896 190604 75948
rect 190644 75896 190696 75948
rect 214104 75939 214156 75948
rect 214104 75905 214113 75939
rect 214113 75905 214147 75939
rect 214147 75905 214156 75939
rect 214104 75896 214156 75905
rect 325700 75939 325752 75948
rect 325700 75905 325709 75939
rect 325709 75905 325743 75939
rect 325743 75905 325752 75939
rect 325700 75896 325752 75905
rect 415032 75896 415084 75948
rect 415124 75896 415176 75948
rect 244280 75871 244332 75880
rect 244280 75837 244289 75871
rect 244289 75837 244323 75871
rect 244323 75837 244332 75871
rect 244280 75828 244332 75837
rect 245752 75871 245804 75880
rect 245752 75837 245761 75871
rect 245761 75837 245795 75871
rect 245795 75837 245804 75871
rect 245752 75828 245804 75837
rect 271880 75871 271932 75880
rect 271880 75837 271889 75871
rect 271889 75837 271923 75871
rect 271923 75837 271932 75871
rect 271880 75828 271932 75837
rect 431592 75871 431644 75880
rect 431592 75837 431601 75871
rect 431601 75837 431635 75871
rect 431635 75837 431644 75871
rect 431592 75828 431644 75837
rect 141056 74536 141108 74588
rect 192208 74579 192260 74588
rect 192208 74545 192217 74579
rect 192217 74545 192251 74579
rect 192251 74545 192260 74579
rect 192208 74536 192260 74545
rect 223672 74579 223724 74588
rect 223672 74545 223681 74579
rect 223681 74545 223715 74579
rect 223715 74545 223724 74579
rect 223672 74536 223724 74545
rect 229192 74579 229244 74588
rect 229192 74545 229201 74579
rect 229201 74545 229235 74579
rect 229235 74545 229244 74579
rect 229192 74536 229244 74545
rect 230388 74579 230440 74588
rect 230388 74545 230397 74579
rect 230397 74545 230431 74579
rect 230431 74545 230440 74579
rect 230388 74536 230440 74545
rect 248420 74579 248472 74588
rect 248420 74545 248429 74579
rect 248429 74545 248463 74579
rect 248463 74545 248472 74579
rect 248420 74536 248472 74545
rect 222384 73176 222436 73228
rect 222476 73176 222528 73228
rect 227904 73176 227956 73228
rect 227996 73176 228048 73228
rect 150716 70456 150768 70508
rect 179696 70456 179748 70508
rect 192208 70456 192260 70508
rect 150624 70320 150676 70372
rect 179604 70320 179656 70372
rect 192116 70320 192168 70372
rect 245844 70320 245896 70372
rect 161756 70252 161808 70304
rect 244372 70252 244424 70304
rect 161756 70116 161808 70168
rect 426072 69683 426124 69692
rect 426072 69649 426081 69683
rect 426081 69649 426115 69683
rect 426115 69649 426124 69683
rect 426072 69640 426124 69649
rect 162952 67736 163004 67788
rect 145012 67600 145064 67652
rect 145104 67600 145156 67652
rect 147956 67600 148008 67652
rect 148048 67600 148100 67652
rect 162952 67600 163004 67652
rect 173992 67600 174044 67652
rect 301964 67643 302016 67652
rect 301964 67609 301973 67643
rect 301973 67609 302007 67643
rect 302007 67609 302016 67643
rect 301964 67600 302016 67609
rect 341432 67600 341484 67652
rect 383292 67600 383344 67652
rect 388812 67600 388864 67652
rect 394424 67600 394476 67652
rect 394516 67600 394568 67652
rect 404084 67600 404136 67652
rect 216864 67575 216916 67584
rect 216864 67541 216873 67575
rect 216873 67541 216907 67575
rect 216907 67541 216916 67575
rect 216864 67532 216916 67541
rect 238944 67575 238996 67584
rect 238944 67541 238953 67575
rect 238953 67541 238987 67575
rect 238987 67541 238996 67575
rect 238944 67532 238996 67541
rect 174084 67464 174136 67516
rect 271972 66240 272024 66292
rect 279792 66240 279844 66292
rect 322664 66240 322716 66292
rect 322756 66240 322808 66292
rect 420460 66240 420512 66292
rect 420552 66240 420604 66292
rect 431592 66283 431644 66292
rect 431592 66249 431601 66283
rect 431601 66249 431635 66283
rect 431635 66249 431644 66283
rect 431592 66240 431644 66249
rect 128820 66215 128872 66224
rect 128820 66181 128829 66215
rect 128829 66181 128863 66215
rect 128863 66181 128872 66215
rect 128820 66172 128872 66181
rect 162952 66215 163004 66224
rect 162952 66181 162961 66215
rect 162961 66181 162995 66215
rect 162995 66181 163004 66215
rect 162952 66172 163004 66181
rect 214104 66172 214156 66224
rect 276112 66172 276164 66224
rect 276296 66172 276348 66224
rect 325700 66172 325752 66224
rect 415032 66215 415084 66224
rect 415032 66181 415041 66215
rect 415041 66181 415075 66215
rect 415075 66181 415084 66215
rect 415032 66172 415084 66181
rect 420460 66104 420512 66156
rect 420644 66104 420696 66156
rect 3332 64812 3384 64864
rect 131672 64812 131724 64864
rect 145012 64812 145064 64864
rect 157340 64855 157392 64864
rect 157340 64821 157349 64855
rect 157349 64821 157383 64855
rect 157383 64821 157392 64855
rect 157340 64812 157392 64821
rect 174084 64812 174136 64864
rect 174268 64812 174320 64864
rect 290464 64855 290516 64864
rect 290464 64821 290473 64855
rect 290473 64821 290507 64855
rect 290507 64821 290516 64855
rect 290464 64812 290516 64821
rect 436836 64812 436888 64864
rect 579804 64812 579856 64864
rect 216864 61047 216916 61056
rect 216864 61013 216873 61047
rect 216873 61013 216907 61047
rect 216907 61013 216916 61047
rect 216864 61004 216916 61013
rect 192116 60800 192168 60852
rect 383292 60800 383344 60852
rect 388812 60800 388864 60852
rect 404084 60800 404136 60852
rect 150532 60664 150584 60716
rect 150716 60664 150768 60716
rect 161572 60664 161624 60716
rect 161756 60664 161808 60716
rect 183652 60664 183704 60716
rect 183836 60664 183888 60716
rect 190644 60664 190696 60716
rect 190828 60664 190880 60716
rect 192116 60664 192168 60716
rect 244372 60664 244424 60716
rect 244556 60664 244608 60716
rect 245844 60664 245896 60716
rect 246028 60664 246080 60716
rect 248420 60664 248472 60716
rect 248604 60664 248656 60716
rect 271972 60664 272024 60716
rect 272156 60664 272208 60716
rect 279884 60664 279936 60716
rect 280068 60664 280120 60716
rect 383200 60664 383252 60716
rect 388720 60664 388772 60716
rect 403992 60664 404044 60716
rect 220728 58624 220780 58676
rect 221004 58624 221056 58676
rect 140872 57944 140924 57996
rect 141056 57944 141108 57996
rect 186228 57944 186280 57996
rect 238944 57987 238996 57996
rect 238944 57953 238953 57987
rect 238953 57953 238987 57987
rect 238987 57953 238996 57987
rect 238944 57944 238996 57953
rect 186320 57876 186372 57928
rect 248236 57876 248288 57928
rect 248328 57876 248380 57928
rect 280068 57919 280120 57928
rect 280068 57885 280077 57919
rect 280077 57885 280111 57919
rect 280111 57885 280120 57919
rect 280068 57876 280120 57885
rect 301780 57919 301832 57928
rect 301780 57885 301789 57919
rect 301789 57885 301823 57919
rect 301823 57885 301832 57919
rect 301780 57876 301832 57885
rect 322756 57876 322808 57928
rect 383200 57919 383252 57928
rect 383200 57885 383209 57919
rect 383209 57885 383243 57919
rect 383243 57885 383252 57919
rect 383200 57876 383252 57885
rect 388720 57919 388772 57928
rect 388720 57885 388729 57919
rect 388729 57885 388763 57919
rect 388763 57885 388772 57919
rect 388720 57876 388772 57885
rect 403992 57919 404044 57928
rect 403992 57885 404001 57919
rect 404001 57885 404035 57919
rect 404035 57885 404044 57919
rect 403992 57876 404044 57885
rect 140872 57851 140924 57860
rect 140872 57817 140881 57851
rect 140881 57817 140915 57851
rect 140915 57817 140924 57851
rect 140872 57808 140924 57817
rect 126244 56652 126296 56704
rect 125968 56584 126020 56636
rect 128912 56584 128964 56636
rect 162952 56627 163004 56636
rect 162952 56593 162961 56627
rect 162961 56593 162995 56627
rect 162995 56593 163004 56627
rect 162952 56584 163004 56593
rect 214104 56584 214156 56636
rect 325516 56627 325568 56636
rect 325516 56593 325525 56627
rect 325525 56593 325559 56627
rect 325559 56593 325568 56627
rect 325516 56584 325568 56593
rect 415032 56627 415084 56636
rect 415032 56593 415041 56627
rect 415041 56593 415075 56627
rect 415075 56593 415084 56627
rect 415032 56584 415084 56593
rect 179420 56559 179472 56568
rect 179420 56525 179429 56559
rect 179429 56525 179463 56559
rect 179463 56525 179472 56559
rect 179420 56516 179472 56525
rect 192116 56559 192168 56568
rect 192116 56525 192125 56559
rect 192125 56525 192159 56559
rect 192159 56525 192168 56559
rect 192116 56516 192168 56525
rect 207204 56516 207256 56568
rect 431592 56516 431644 56568
rect 431776 56516 431828 56568
rect 144920 55267 144972 55276
rect 144920 55233 144929 55267
rect 144929 55233 144963 55267
rect 144963 55233 144972 55267
rect 144920 55224 144972 55233
rect 157432 55224 157484 55276
rect 290556 55224 290608 55276
rect 186320 55156 186372 55208
rect 426072 53116 426124 53168
rect 426256 53116 426308 53168
rect 157432 51756 157484 51808
rect 415032 51280 415084 51332
rect 415216 51280 415268 51332
rect 223672 51144 223724 51196
rect 229192 51144 229244 51196
rect 290556 51144 290608 51196
rect 341524 51187 341576 51196
rect 341524 51153 341533 51187
rect 341533 51153 341567 51187
rect 341567 51153 341576 51187
rect 341524 51144 341576 51153
rect 125968 51119 126020 51128
rect 125968 51085 125977 51119
rect 125977 51085 126011 51119
rect 126011 51085 126020 51119
rect 125968 51076 126020 51085
rect 148048 51076 148100 51128
rect 161756 51076 161808 51128
rect 128912 51008 128964 51060
rect 147956 51008 148008 51060
rect 129004 50940 129056 50992
rect 272156 51076 272208 51128
rect 223672 51008 223724 51060
rect 229192 51008 229244 51060
rect 272064 51008 272116 51060
rect 280068 51051 280120 51060
rect 280068 51017 280077 51051
rect 280077 51017 280111 51051
rect 280111 51017 280120 51051
rect 280068 51008 280120 51017
rect 161756 50872 161808 50924
rect 140964 48288 141016 48340
rect 162860 48288 162912 48340
rect 162952 48288 163004 48340
rect 183836 48288 183888 48340
rect 183928 48288 183980 48340
rect 301872 48288 301924 48340
rect 322664 48331 322716 48340
rect 322664 48297 322673 48331
rect 322673 48297 322707 48331
rect 322707 48297 322716 48331
rect 322664 48288 322716 48297
rect 383292 48288 383344 48340
rect 388812 48288 388864 48340
rect 394424 48288 394476 48340
rect 394516 48288 394568 48340
rect 404084 48288 404136 48340
rect 272064 48152 272116 48204
rect 290372 47039 290424 47048
rect 290372 47005 290381 47039
rect 290381 47005 290415 47039
rect 290415 47005 290424 47039
rect 290372 46996 290424 47005
rect 125968 46971 126020 46980
rect 125968 46937 125977 46971
rect 125977 46937 126011 46971
rect 126011 46937 126020 46971
rect 125968 46928 126020 46937
rect 179512 46928 179564 46980
rect 192116 46971 192168 46980
rect 192116 46937 192125 46971
rect 192125 46937 192159 46971
rect 192159 46937 192168 46971
rect 192116 46928 192168 46937
rect 133328 46903 133380 46912
rect 133328 46869 133337 46903
rect 133337 46869 133371 46903
rect 133371 46869 133380 46903
rect 133328 46860 133380 46869
rect 145012 46860 145064 46912
rect 147956 46860 148008 46912
rect 150808 46860 150860 46912
rect 162952 46903 163004 46912
rect 162952 46869 162961 46903
rect 162961 46869 162995 46903
rect 162995 46869 163004 46903
rect 162952 46860 163004 46869
rect 214104 46903 214156 46912
rect 214104 46869 214113 46903
rect 214113 46869 214147 46903
rect 214147 46869 214156 46903
rect 214104 46860 214156 46869
rect 215392 46903 215444 46912
rect 215392 46869 215401 46903
rect 215401 46869 215435 46903
rect 215435 46869 215444 46903
rect 215392 46860 215444 46869
rect 248328 46903 248380 46912
rect 248328 46869 248337 46903
rect 248337 46869 248371 46903
rect 248371 46869 248380 46903
rect 248328 46860 248380 46869
rect 276112 46860 276164 46912
rect 290372 46860 290424 46912
rect 325700 46903 325752 46912
rect 325700 46869 325709 46903
rect 325709 46869 325743 46903
rect 325743 46869 325752 46903
rect 325700 46860 325752 46869
rect 420460 46860 420512 46912
rect 420644 46860 420696 46912
rect 425980 46903 426032 46912
rect 425980 46869 425989 46903
rect 425989 46869 426023 46903
rect 426023 46869 426032 46903
rect 425980 46860 426032 46869
rect 431500 46860 431552 46912
rect 431592 46860 431644 46912
rect 125968 46792 126020 46844
rect 126152 46792 126204 46844
rect 144920 46792 144972 46844
rect 147864 46792 147916 46844
rect 192116 45883 192168 45892
rect 192116 45849 192125 45883
rect 192125 45849 192159 45883
rect 192159 45849 192168 45883
rect 192116 45840 192168 45849
rect 173992 45568 174044 45620
rect 174268 45568 174320 45620
rect 186228 45611 186280 45620
rect 186228 45577 186237 45611
rect 186237 45577 186271 45611
rect 186271 45577 186280 45611
rect 186228 45568 186280 45577
rect 341524 45611 341576 45620
rect 341524 45577 341533 45611
rect 341533 45577 341567 45611
rect 341567 45577 341576 45611
rect 341524 45568 341576 45577
rect 183928 45500 183980 45552
rect 190736 45500 190788 45552
rect 414940 45543 414992 45552
rect 414940 45509 414949 45543
rect 414949 45509 414983 45543
rect 414983 45509 414992 45543
rect 414940 45500 414992 45509
rect 341524 45432 341576 45484
rect 221004 44140 221056 44192
rect 221188 44140 221240 44192
rect 248696 42032 248748 42084
rect 248880 42032 248932 42084
rect 133604 41352 133656 41404
rect 580172 41352 580224 41404
rect 192208 41284 192260 41336
rect 227904 41284 227956 41336
rect 228180 41284 228232 41336
rect 271880 41327 271932 41336
rect 271880 41293 271889 41327
rect 271889 41293 271923 41327
rect 271923 41293 271932 41327
rect 271880 41284 271932 41293
rect 173992 40715 174044 40724
rect 173992 40681 174001 40715
rect 174001 40681 174035 40715
rect 174035 40681 174044 40715
rect 173992 40672 174044 40681
rect 186320 40672 186372 40724
rect 190644 40715 190696 40724
rect 190644 40681 190653 40715
rect 190653 40681 190687 40715
rect 190687 40681 190696 40715
rect 190644 40672 190696 40681
rect 140872 38632 140924 38684
rect 141056 38632 141108 38684
rect 157616 38675 157668 38684
rect 157616 38641 157625 38675
rect 157625 38641 157659 38675
rect 157659 38641 157668 38675
rect 157616 38632 157668 38641
rect 207480 38675 207532 38684
rect 207480 38641 207489 38675
rect 207489 38641 207523 38675
rect 207523 38641 207532 38675
rect 207480 38632 207532 38641
rect 244280 38632 244332 38684
rect 244556 38632 244608 38684
rect 245752 38632 245804 38684
rect 246028 38632 246080 38684
rect 279884 38632 279936 38684
rect 280068 38632 280120 38684
rect 271880 38607 271932 38616
rect 271880 38573 271889 38607
rect 271889 38573 271923 38607
rect 271923 38573 271932 38607
rect 271880 38564 271932 38573
rect 322756 38564 322808 38616
rect 383200 38607 383252 38616
rect 383200 38573 383209 38607
rect 383209 38573 383243 38607
rect 383243 38573 383252 38607
rect 383200 38564 383252 38573
rect 403992 38607 404044 38616
rect 403992 38573 404001 38607
rect 404001 38573 404035 38607
rect 404035 38573 404044 38607
rect 403992 38564 404044 38573
rect 290648 38539 290700 38548
rect 290648 38505 290657 38539
rect 290657 38505 290691 38539
rect 290691 38505 290700 38539
rect 290648 38496 290700 38505
rect 341432 38267 341484 38276
rect 341432 38233 341441 38267
rect 341441 38233 341475 38267
rect 341475 38233 341484 38267
rect 341432 38224 341484 38233
rect 133512 37272 133564 37324
rect 150624 37315 150676 37324
rect 150624 37281 150633 37315
rect 150633 37281 150667 37315
rect 150667 37281 150676 37315
rect 150624 37272 150676 37281
rect 162952 37315 163004 37324
rect 162952 37281 162961 37315
rect 162961 37281 162995 37315
rect 162995 37281 163004 37315
rect 162952 37272 163004 37281
rect 214104 37315 214156 37324
rect 214104 37281 214113 37315
rect 214113 37281 214147 37315
rect 214147 37281 214156 37315
rect 214104 37272 214156 37281
rect 215392 37315 215444 37324
rect 215392 37281 215401 37315
rect 215401 37281 215435 37315
rect 215435 37281 215444 37315
rect 215392 37272 215444 37281
rect 248328 37315 248380 37324
rect 248328 37281 248337 37315
rect 248337 37281 248371 37315
rect 248371 37281 248380 37315
rect 248328 37272 248380 37281
rect 426072 37272 426124 37324
rect 179420 37247 179472 37256
rect 179420 37213 179429 37247
rect 179429 37213 179463 37247
rect 179463 37213 179472 37247
rect 179420 37204 179472 37213
rect 244280 37247 244332 37256
rect 244280 37213 244289 37247
rect 244289 37213 244323 37247
rect 244323 37213 244332 37247
rect 244280 37204 244332 37213
rect 245752 37247 245804 37256
rect 245752 37213 245761 37247
rect 245761 37213 245795 37247
rect 245795 37213 245804 37247
rect 245752 37204 245804 37213
rect 431592 37247 431644 37256
rect 431592 37213 431601 37247
rect 431601 37213 431635 37247
rect 431635 37213 431644 37247
rect 431592 37204 431644 37213
rect 415032 35912 415084 35964
rect 3424 35844 3476 35896
rect 436192 35844 436244 35896
rect 227904 34416 227956 34468
rect 227996 34416 228048 34468
rect 150624 33804 150676 33856
rect 150808 33804 150860 33856
rect 129004 31764 129056 31816
rect 223672 31832 223724 31884
rect 301964 31832 302016 31884
rect 290648 31764 290700 31816
rect 128912 31696 128964 31748
rect 192208 31739 192260 31748
rect 192208 31705 192217 31739
rect 192217 31705 192251 31739
rect 192251 31705 192260 31739
rect 192208 31696 192260 31705
rect 223580 31696 223632 31748
rect 279884 31696 279936 31748
rect 280068 31696 280120 31748
rect 302056 31696 302108 31748
rect 388720 31696 388772 31748
rect 388904 31696 388956 31748
rect 244372 31628 244424 31680
rect 245844 31628 245896 31680
rect 290648 31628 290700 31680
rect 341432 31628 341484 31680
rect 341524 31628 341576 31680
rect 431684 31628 431736 31680
rect 132408 30268 132460 30320
rect 580172 30268 580224 30320
rect 276112 29087 276164 29096
rect 276112 29053 276121 29087
rect 276121 29053 276155 29087
rect 276155 29053 276164 29087
rect 276112 29044 276164 29053
rect 325700 29087 325752 29096
rect 325700 29053 325709 29087
rect 325709 29053 325743 29087
rect 325743 29053 325752 29087
rect 325700 29044 325752 29053
rect 133328 28976 133380 29028
rect 133512 28976 133564 29028
rect 161756 28976 161808 29028
rect 161848 28976 161900 29028
rect 271972 28976 272024 29028
rect 322664 29019 322716 29028
rect 322664 28985 322673 29019
rect 322673 28985 322707 29019
rect 322707 28985 322716 29019
rect 322664 28976 322716 28985
rect 383292 28976 383344 29028
rect 394424 28976 394476 29028
rect 394516 28976 394568 29028
rect 404084 28976 404136 29028
rect 128912 28908 128964 28960
rect 140964 28908 141016 28960
rect 207480 28951 207532 28960
rect 207480 28917 207489 28951
rect 207489 28917 207523 28951
rect 207523 28917 207532 28951
rect 207480 28908 207532 28917
rect 280068 28908 280120 28960
rect 129004 28840 129056 28892
rect 179512 27616 179564 27668
rect 183744 27659 183796 27668
rect 183744 27625 183753 27659
rect 183753 27625 183787 27659
rect 183787 27625 183796 27659
rect 183744 27616 183796 27625
rect 248512 27616 248564 27668
rect 248696 27616 248748 27668
rect 126060 27548 126112 27600
rect 133328 27591 133380 27600
rect 133328 27557 133337 27591
rect 133337 27557 133371 27591
rect 133371 27557 133380 27591
rect 133328 27548 133380 27557
rect 162952 27591 163004 27600
rect 162952 27557 162961 27591
rect 162961 27557 162995 27591
rect 162995 27557 163004 27591
rect 162952 27548 163004 27557
rect 190644 27548 190696 27600
rect 192208 27591 192260 27600
rect 192208 27557 192217 27591
rect 192217 27557 192251 27591
rect 192251 27557 192260 27591
rect 192208 27548 192260 27557
rect 214104 27591 214156 27600
rect 214104 27557 214113 27591
rect 214113 27557 214147 27591
rect 214147 27557 214156 27591
rect 214104 27548 214156 27557
rect 215392 27591 215444 27600
rect 215392 27557 215401 27591
rect 215401 27557 215435 27591
rect 215435 27557 215444 27591
rect 215392 27548 215444 27557
rect 276112 27591 276164 27600
rect 276112 27557 276121 27591
rect 276121 27557 276155 27591
rect 276155 27557 276164 27591
rect 276112 27548 276164 27557
rect 325700 27591 325752 27600
rect 325700 27557 325709 27591
rect 325709 27557 325743 27591
rect 325743 27557 325752 27591
rect 325700 27548 325752 27557
rect 420460 27591 420512 27600
rect 420460 27557 420469 27591
rect 420469 27557 420503 27591
rect 420503 27557 420512 27591
rect 420460 27548 420512 27557
rect 186228 27115 186280 27124
rect 186228 27081 186237 27115
rect 186237 27081 186271 27115
rect 186271 27081 186280 27115
rect 186228 27072 186280 27081
rect 174084 26256 174136 26308
rect 183744 26231 183796 26240
rect 183744 26197 183753 26231
rect 183753 26197 183787 26231
rect 183787 26197 183796 26231
rect 183744 26188 183796 26197
rect 192208 26231 192260 26240
rect 192208 26197 192217 26231
rect 192217 26197 192251 26231
rect 192251 26197 192260 26231
rect 301872 26231 301924 26240
rect 192208 26188 192260 26197
rect 301872 26197 301881 26231
rect 301881 26197 301915 26231
rect 301915 26197 301924 26231
rect 301872 26188 301924 26197
rect 415032 26231 415084 26240
rect 415032 26197 415041 26231
rect 415041 26197 415075 26231
rect 415075 26197 415084 26231
rect 415032 26188 415084 26197
rect 431684 26188 431736 26240
rect 383384 25279 383436 25288
rect 383384 25245 383393 25279
rect 383393 25245 383427 25279
rect 383427 25245 383436 25279
rect 383384 25236 383436 25245
rect 222384 24896 222436 24948
rect 221004 24828 221056 24880
rect 221188 24828 221240 24880
rect 230388 24760 230440 24812
rect 147864 24148 147916 24200
rect 148048 24148 148100 24200
rect 388720 24148 388772 24200
rect 388904 24148 388956 24200
rect 222292 23511 222344 23520
rect 222292 23477 222301 23511
rect 222301 23477 222335 23511
rect 222335 23477 222344 23511
rect 222292 23468 222344 23477
rect 161756 22763 161808 22772
rect 161756 22729 161765 22763
rect 161765 22729 161799 22763
rect 161799 22729 161808 22763
rect 161756 22720 161808 22729
rect 238944 22219 238996 22228
rect 238944 22185 238953 22219
rect 238953 22185 238987 22219
rect 238987 22185 238996 22219
rect 238944 22176 238996 22185
rect 174084 22108 174136 22160
rect 3148 22040 3200 22092
rect 132224 22040 132276 22092
rect 144920 22040 144972 22092
rect 145104 22040 145156 22092
rect 404084 22108 404136 22160
rect 244372 22040 244424 22092
rect 244556 22040 244608 22092
rect 245844 22040 245896 22092
rect 246028 22040 246080 22092
rect 248420 22040 248472 22092
rect 248604 22040 248656 22092
rect 290740 22040 290792 22092
rect 290924 22040 290976 22092
rect 403992 22040 404044 22092
rect 174084 21972 174136 22024
rect 221004 20068 221056 20120
rect 227996 20000 228048 20052
rect 221004 19932 221056 19984
rect 140872 19431 140924 19440
rect 140872 19397 140881 19431
rect 140881 19397 140915 19431
rect 140915 19397 140924 19431
rect 140872 19388 140924 19397
rect 207204 19388 207256 19440
rect 150624 19320 150676 19372
rect 150716 19320 150768 19372
rect 238944 19363 238996 19372
rect 238944 19329 238953 19363
rect 238953 19329 238987 19363
rect 238987 19329 238996 19363
rect 238944 19320 238996 19329
rect 279976 19363 280028 19372
rect 279976 19329 279985 19363
rect 279985 19329 280019 19363
rect 280019 19329 280028 19363
rect 279976 19320 280028 19329
rect 383384 19363 383436 19372
rect 383384 19329 383393 19363
rect 383393 19329 383427 19363
rect 383427 19329 383436 19363
rect 383384 19320 383436 19329
rect 133328 19295 133380 19304
rect 133328 19261 133337 19295
rect 133337 19261 133371 19295
rect 133371 19261 133380 19295
rect 133328 19252 133380 19261
rect 140872 19295 140924 19304
rect 140872 19261 140881 19295
rect 140881 19261 140915 19295
rect 140915 19261 140924 19295
rect 140872 19252 140924 19261
rect 179696 19295 179748 19304
rect 179696 19261 179705 19295
rect 179705 19261 179739 19295
rect 179739 19261 179748 19295
rect 179696 19252 179748 19261
rect 207296 19252 207348 19304
rect 238668 19252 238720 19304
rect 290924 19295 290976 19304
rect 290924 19261 290933 19295
rect 290933 19261 290967 19295
rect 290967 19261 290976 19295
rect 290924 19252 290976 19261
rect 425980 19252 426032 19304
rect 426072 19252 426124 19304
rect 162952 18003 163004 18012
rect 162952 17969 162961 18003
rect 162961 17969 162995 18003
rect 162995 17969 163004 18003
rect 162952 17960 163004 17969
rect 190460 18003 190512 18012
rect 190460 17969 190469 18003
rect 190469 17969 190503 18003
rect 190503 17969 190512 18003
rect 190460 17960 190512 17969
rect 276112 18003 276164 18012
rect 276112 17969 276121 18003
rect 276121 17969 276155 18003
rect 276155 17969 276164 18003
rect 276112 17960 276164 17969
rect 420552 17960 420604 18012
rect 436744 17892 436796 17944
rect 579804 17892 579856 17944
rect 183836 16600 183888 16652
rect 192208 16643 192260 16652
rect 192208 16609 192217 16643
rect 192217 16609 192251 16643
rect 192251 16609 192260 16643
rect 192208 16600 192260 16609
rect 415032 16643 415084 16652
rect 415032 16609 415041 16643
rect 415041 16609 415075 16643
rect 415075 16609 415084 16643
rect 415032 16600 415084 16609
rect 431500 16643 431552 16652
rect 431500 16609 431509 16643
rect 431509 16609 431543 16643
rect 431543 16609 431552 16643
rect 431500 16600 431552 16609
rect 274824 15895 274876 15904
rect 274824 15861 274833 15895
rect 274833 15861 274867 15895
rect 274867 15861 274876 15895
rect 274824 15852 274876 15861
rect 222292 15172 222344 15224
rect 222384 15104 222436 15156
rect 162952 12452 163004 12504
rect 168472 12452 168524 12504
rect 186228 12452 186280 12504
rect 208400 12452 208452 12504
rect 208584 12452 208636 12504
rect 237288 12520 237340 12572
rect 383292 12563 383344 12572
rect 383292 12529 383301 12563
rect 383301 12529 383335 12563
rect 383335 12529 383344 12563
rect 383292 12520 383344 12529
rect 237196 12452 237248 12504
rect 162860 12384 162912 12436
rect 186044 12384 186096 12436
rect 237104 12384 237156 12436
rect 248328 12452 248380 12504
rect 276112 12452 276164 12504
rect 394332 12452 394384 12504
rect 247960 12384 248012 12436
rect 237196 12316 237248 12368
rect 321744 12384 321796 12436
rect 276480 12316 276532 12368
rect 322756 12316 322808 12368
rect 415032 12452 415084 12504
rect 420552 12452 420604 12504
rect 414940 12384 414992 12436
rect 420460 12384 420512 12436
rect 463700 12384 463752 12436
rect 464344 12384 464396 12436
rect 394424 12316 394476 12368
rect 161756 11883 161808 11892
rect 161756 11849 161765 11883
rect 161765 11849 161799 11883
rect 161799 11849 161808 11883
rect 161756 11840 161808 11849
rect 371056 10684 371108 10736
rect 459652 10684 459704 10736
rect 372344 10616 372396 10668
rect 463240 10616 463292 10668
rect 375196 10548 375248 10600
rect 466828 10548 466880 10600
rect 376576 10480 376628 10532
rect 470324 10480 470376 10532
rect 377956 10412 378008 10464
rect 473360 10412 473412 10464
rect 380808 10344 380860 10396
rect 477684 10344 477736 10396
rect 382096 10276 382148 10328
rect 481088 10276 481140 10328
rect 125968 9707 126020 9716
rect 125968 9673 125977 9707
rect 125977 9673 126011 9707
rect 126011 9673 126020 9707
rect 125968 9664 126020 9673
rect 133144 9664 133196 9716
rect 133328 9664 133380 9716
rect 141056 9664 141108 9716
rect 168380 9707 168432 9716
rect 168380 9673 168389 9707
rect 168389 9673 168423 9707
rect 168423 9673 168432 9707
rect 168380 9664 168432 9673
rect 179788 9664 179840 9716
rect 207204 9707 207256 9716
rect 207204 9673 207213 9707
rect 207213 9673 207247 9707
rect 207247 9673 207256 9707
rect 207204 9664 207256 9673
rect 214196 9664 214248 9716
rect 215484 9664 215536 9716
rect 238392 9707 238444 9716
rect 238392 9673 238401 9707
rect 238401 9673 238435 9707
rect 238435 9673 238444 9707
rect 238392 9664 238444 9673
rect 275284 9664 275336 9716
rect 280436 9664 280488 9716
rect 281264 9664 281316 9716
rect 282920 9664 282972 9716
rect 283380 9664 283432 9716
rect 290924 9707 290976 9716
rect 290924 9673 290933 9707
rect 290933 9673 290967 9707
rect 290967 9673 290976 9707
rect 290924 9664 290976 9673
rect 326252 9664 326304 9716
rect 383292 9707 383344 9716
rect 383292 9673 383301 9707
rect 383301 9673 383335 9707
rect 383335 9673 383344 9707
rect 383292 9664 383344 9673
rect 57612 9596 57664 9648
rect 162860 9596 162912 9648
rect 368388 9596 368440 9648
rect 454868 9596 454920 9648
rect 58808 9528 58860 9580
rect 164332 9528 164384 9580
rect 371148 9528 371200 9580
rect 458456 9528 458508 9580
rect 55220 9460 55272 9512
rect 161756 9460 161808 9512
rect 372436 9460 372488 9512
rect 462044 9460 462096 9512
rect 51632 9392 51684 9444
rect 160192 9392 160244 9444
rect 419448 9392 419500 9444
rect 552388 9392 552440 9444
rect 43352 9324 43404 9376
rect 156052 9324 156104 9376
rect 420460 9324 420512 9376
rect 555976 9324 556028 9376
rect 40960 9256 41012 9308
rect 154672 9256 154724 9308
rect 422116 9256 422168 9308
rect 559564 9256 559616 9308
rect 36176 9188 36228 9240
rect 151820 9188 151872 9240
rect 409512 9188 409564 9240
rect 409788 9188 409840 9240
rect 424968 9188 425020 9240
rect 563152 9188 563204 9240
rect 18328 9120 18380 9172
rect 135444 9120 135496 9172
rect 350356 9120 350408 9172
rect 420368 9120 420420 9172
rect 425980 9120 426032 9172
rect 566740 9120 566792 9172
rect 20720 9052 20772 9104
rect 143632 9052 143684 9104
rect 353208 9052 353260 9104
rect 423956 9052 424008 9104
rect 427636 9052 427688 9104
rect 570236 9052 570288 9104
rect 11244 8984 11296 9036
rect 139492 8984 139544 9036
rect 354496 8984 354548 9036
rect 427544 8984 427596 9036
rect 431500 8984 431552 9036
rect 577412 8984 577464 9036
rect 5264 8916 5316 8968
rect 136824 8916 136876 8968
rect 143264 8916 143316 8968
rect 207204 8916 207256 8968
rect 355876 8916 355928 8968
rect 431132 8916 431184 8968
rect 433156 8916 433208 8968
rect 581000 8916 581052 8968
rect 64788 8848 64840 8900
rect 167092 8848 167144 8900
rect 369768 8848 369820 8900
rect 456064 8848 456116 8900
rect 71872 8780 71924 8832
rect 169852 8780 169904 8832
rect 366916 8780 366968 8832
rect 452476 8780 452528 8832
rect 79048 8712 79100 8764
rect 173992 8712 174044 8764
rect 365536 8712 365588 8764
rect 448980 8712 449032 8764
rect 120632 8644 120684 8696
rect 175464 8644 175516 8696
rect 361396 8644 361448 8696
rect 441804 8644 441856 8696
rect 106372 8576 106424 8628
rect 133144 8576 133196 8628
rect 364248 8576 364300 8628
rect 445392 8576 445444 8628
rect 360016 8508 360068 8560
rect 438216 8508 438268 8560
rect 358636 8440 358688 8492
rect 434628 8440 434680 8492
rect 129280 8304 129332 8356
rect 302056 8304 302108 8356
rect 3424 8236 3476 8288
rect 131764 8236 131816 8288
rect 133788 8236 133840 8288
rect 203064 8236 203116 8288
rect 384948 8236 385000 8288
rect 486976 8236 487028 8288
rect 114744 8168 114796 8220
rect 191932 8168 191984 8220
rect 387616 8168 387668 8220
rect 490564 8168 490616 8220
rect 107568 8100 107620 8152
rect 189172 8100 189224 8152
rect 388904 8100 388956 8152
rect 494152 8100 494204 8152
rect 100484 8032 100536 8084
rect 184940 8032 184992 8084
rect 390468 8032 390520 8084
rect 497740 8032 497792 8084
rect 48136 7964 48188 8016
rect 158812 7964 158864 8016
rect 393136 7964 393188 8016
rect 501236 7964 501288 8016
rect 13636 7896 13688 7948
rect 141056 7896 141108 7948
rect 394332 7896 394384 7948
rect 504824 7896 504876 7948
rect 7656 7828 7708 7880
rect 136732 7828 136784 7880
rect 140872 7828 140924 7880
rect 205640 7828 205692 7880
rect 395896 7828 395948 7880
rect 508412 7828 508464 7880
rect 4068 7760 4120 7812
rect 135260 7760 135312 7812
rect 139676 7760 139728 7812
rect 205732 7760 205784 7812
rect 413928 7760 413980 7812
rect 541716 7760 541768 7812
rect 1676 7692 1728 7744
rect 134064 7692 134116 7744
rect 136088 7692 136140 7744
rect 202972 7692 203024 7744
rect 344744 7692 344796 7744
rect 409696 7692 409748 7744
rect 414940 7692 414992 7744
rect 545304 7692 545356 7744
rect 2872 7624 2924 7676
rect 135352 7624 135404 7676
rect 137284 7624 137336 7676
rect 204352 7624 204404 7676
rect 347688 7624 347740 7676
rect 413284 7624 413336 7676
rect 416596 7624 416648 7676
rect 548892 7624 548944 7676
rect 572 7556 624 7608
rect 133880 7556 133932 7608
rect 134892 7556 134944 7608
rect 202880 7556 202932 7608
rect 348976 7556 349028 7608
rect 416780 7556 416832 7608
rect 417976 7556 418028 7608
rect 430488 7556 430540 7608
rect 573824 7556 573876 7608
rect 121828 7488 121880 7540
rect 196072 7488 196124 7540
rect 383292 7488 383344 7540
rect 126612 7420 126664 7472
rect 198832 7420 198884 7472
rect 367008 7420 367060 7472
rect 451280 7420 451332 7472
rect 127624 7352 127676 7404
rect 77852 7284 77904 7336
rect 117136 7216 117188 7268
rect 84936 7148 84988 7200
rect 125416 7284 125468 7336
rect 197452 7352 197504 7404
rect 365628 7352 365680 7404
rect 447784 7352 447836 7404
rect 477500 7488 477552 7540
rect 478696 7488 478748 7540
rect 483480 7352 483532 7404
rect 129004 7284 129056 7336
rect 200212 7284 200264 7336
rect 362868 7284 362920 7336
rect 444196 7284 444248 7336
rect 127808 7216 127860 7268
rect 198740 7216 198792 7268
rect 361488 7216 361540 7268
rect 440608 7216 440660 7268
rect 95700 7080 95752 7132
rect 129096 7148 129148 7200
rect 131396 7148 131448 7200
rect 201592 7148 201644 7200
rect 360108 7148 360160 7200
rect 437020 7148 437072 7200
rect 129188 7080 129240 7132
rect 130200 7080 130252 7132
rect 200120 7080 200172 7132
rect 358728 7080 358780 7132
rect 435824 7080 435876 7132
rect 132592 7012 132644 7064
rect 201500 7012 201552 7064
rect 416872 7012 416924 7064
rect 227812 6919 227864 6928
rect 227812 6885 227821 6919
rect 227821 6885 227855 6919
rect 227855 6885 227864 6919
rect 227812 6876 227864 6885
rect 230112 6919 230164 6928
rect 230112 6885 230121 6919
rect 230121 6885 230155 6919
rect 230155 6885 230164 6919
rect 230112 6876 230164 6885
rect 94504 6808 94556 6860
rect 182272 6808 182324 6860
rect 317236 6808 317288 6860
rect 356152 6808 356204 6860
rect 391756 6808 391808 6860
rect 498936 6808 498988 6860
rect 93308 6740 93360 6792
rect 180984 6740 181036 6792
rect 326896 6740 326948 6792
rect 374000 6740 374052 6792
rect 393228 6740 393280 6792
rect 502432 6740 502484 6792
rect 90916 6672 90968 6724
rect 180892 6672 180944 6724
rect 328184 6672 328236 6724
rect 377588 6672 377640 6724
rect 394608 6672 394660 6724
rect 506020 6672 506072 6724
rect 86132 6604 86184 6656
rect 178132 6604 178184 6656
rect 331036 6604 331088 6656
rect 381176 6604 381228 6656
rect 397368 6604 397420 6656
rect 509608 6604 509660 6656
rect 82636 6536 82688 6588
rect 175372 6536 175424 6588
rect 332416 6536 332468 6588
rect 384672 6536 384724 6588
rect 398656 6536 398708 6588
rect 513196 6536 513248 6588
rect 8852 6468 8904 6520
rect 103520 6468 103572 6520
rect 105176 6468 105228 6520
rect 187700 6468 187752 6520
rect 336648 6468 336700 6520
rect 391848 6468 391900 6520
rect 399944 6468 399996 6520
rect 516784 6468 516836 6520
rect 75460 6400 75512 6452
rect 172612 6400 172664 6452
rect 333704 6400 333756 6452
rect 388260 6400 388312 6452
rect 402796 6400 402848 6452
rect 520280 6400 520332 6452
rect 68284 6332 68336 6384
rect 168380 6332 168432 6384
rect 337936 6332 337988 6384
rect 395436 6332 395488 6384
rect 404176 6332 404228 6384
rect 523868 6332 523920 6384
rect 61200 6264 61252 6316
rect 164424 6264 164476 6316
rect 342168 6264 342220 6316
rect 402520 6264 402572 6316
rect 408408 6264 408460 6316
rect 531044 6264 531096 6316
rect 54024 6196 54076 6248
rect 161480 6196 161532 6248
rect 339316 6196 339368 6248
rect 399024 6196 399076 6248
rect 405556 6196 405608 6248
rect 527456 6196 527508 6248
rect 44548 6128 44600 6180
rect 155960 6128 156012 6180
rect 157524 6128 157576 6180
rect 214196 6128 214248 6180
rect 343456 6128 343508 6180
rect 406108 6128 406160 6180
rect 409604 6128 409656 6180
rect 534540 6128 534592 6180
rect 101588 6060 101640 6112
rect 186504 6060 186556 6112
rect 318708 6060 318760 6112
rect 358544 6060 358596 6112
rect 388996 6060 389048 6112
rect 495348 6060 495400 6112
rect 98092 5992 98144 6044
rect 183836 5992 183888 6044
rect 317144 5992 317196 6044
rect 354956 5992 355008 6044
rect 387708 5992 387760 6044
rect 491760 5992 491812 6044
rect 108764 5924 108816 5976
rect 189080 5924 189132 5976
rect 315948 5924 316000 5976
rect 352564 5924 352616 5976
rect 383476 5924 383528 5976
rect 484584 5924 484636 5976
rect 112352 5856 112404 5908
rect 191840 5856 191892 5908
rect 315856 5856 315908 5908
rect 351368 5856 351420 5908
rect 386328 5856 386380 5908
rect 488172 5856 488224 5908
rect 113548 5788 113600 5840
rect 192208 5788 192260 5840
rect 379336 5788 379388 5840
rect 476304 5788 476356 5840
rect 115940 5720 115992 5772
rect 193220 5720 193272 5772
rect 382188 5720 382240 5772
rect 479892 5720 479944 5772
rect 119436 5652 119488 5704
rect 194692 5652 194744 5704
rect 378048 5652 378100 5704
rect 472716 5652 472768 5704
rect 123024 5584 123076 5636
rect 197360 5584 197412 5636
rect 373908 5584 373960 5636
rect 465632 5584 465684 5636
rect 150440 5516 150492 5568
rect 211252 5516 211304 5568
rect 376668 5516 376720 5568
rect 469128 5516 469180 5568
rect 73068 5448 73120 5500
rect 171232 5448 171284 5500
rect 171692 5448 171744 5500
rect 211160 5448 211212 5500
rect 335176 5448 335228 5500
rect 390652 5448 390704 5500
rect 415308 5448 415360 5500
rect 544108 5448 544160 5500
rect 69480 5380 69532 5432
rect 169944 5380 169996 5432
rect 187240 5380 187292 5432
rect 229100 5380 229152 5432
rect 339408 5380 339460 5432
rect 397828 5380 397880 5432
rect 416688 5380 416740 5432
rect 547696 5380 547748 5432
rect 65984 5312 66036 5364
rect 167000 5312 167052 5364
rect 170588 5312 170640 5364
rect 221004 5312 221056 5364
rect 340696 5312 340748 5364
rect 401324 5312 401376 5364
rect 418068 5312 418120 5364
rect 551192 5312 551244 5364
rect 62396 5244 62448 5296
rect 165712 5244 165764 5296
rect 167092 5244 167144 5296
rect 219532 5244 219584 5296
rect 343548 5244 343600 5296
rect 404912 5244 404964 5296
rect 420828 5244 420880 5296
rect 554780 5244 554832 5296
rect 37372 5176 37424 5228
rect 153292 5176 153344 5228
rect 163504 5176 163556 5228
rect 218152 5176 218204 5228
rect 344836 5176 344888 5228
rect 408684 5176 408736 5228
rect 422208 5176 422260 5228
rect 558368 5176 558420 5228
rect 33876 5108 33928 5160
rect 150716 5108 150768 5160
rect 158720 5108 158772 5160
rect 215300 5108 215352 5160
rect 346308 5108 346360 5160
rect 412088 5108 412140 5160
rect 426348 5108 426400 5160
rect 565544 5108 565596 5160
rect 29092 5040 29144 5092
rect 148048 5040 148100 5092
rect 155132 5040 155184 5092
rect 213920 5040 213972 5092
rect 349068 5040 349120 5092
rect 415676 5040 415728 5092
rect 423588 5040 423640 5092
rect 561956 5040 562008 5092
rect 26700 4972 26752 5024
rect 147772 4972 147824 5024
rect 152740 4972 152792 5024
rect 212632 4972 212684 5024
rect 219348 4972 219400 5024
rect 246028 4972 246080 5024
rect 350448 4972 350500 5024
rect 419172 4972 419224 5024
rect 427728 4972 427780 5024
rect 569040 4972 569092 5024
rect 21916 4904 21968 4956
rect 145104 4904 145156 4956
rect 149244 4904 149296 4956
rect 209872 4904 209924 4956
rect 215852 4904 215904 4956
rect 244556 4904 244608 4956
rect 310428 4904 310480 4956
rect 341892 4904 341944 4956
rect 351736 4904 351788 4956
rect 422760 4904 422812 4956
rect 429108 4904 429160 4956
rect 572628 4904 572680 4956
rect 12440 4836 12492 4888
rect 139400 4836 139452 4888
rect 142068 4836 142120 4888
rect 207020 4836 207072 4888
rect 212264 4836 212316 4888
rect 242992 4836 243044 4888
rect 314568 4836 314620 4888
rect 349068 4836 349120 4888
rect 354588 4836 354640 4888
rect 426348 4836 426400 4888
rect 431868 4836 431920 4888
rect 576216 4836 576268 4888
rect 17224 4768 17276 4820
rect 142252 4768 142304 4820
rect 145656 4768 145708 4820
rect 208400 4768 208452 4820
rect 208676 4768 208728 4820
rect 240140 4768 240192 4820
rect 313096 4768 313148 4820
rect 347872 4768 347924 4820
rect 355968 4768 356020 4820
rect 429936 4768 429988 4820
rect 433248 4768 433300 4820
rect 579804 4768 579856 4820
rect 76656 4700 76708 4752
rect 172520 4700 172572 4752
rect 203800 4700 203852 4752
rect 237472 4700 237524 4752
rect 338028 4700 338080 4752
rect 394240 4700 394292 4752
rect 412548 4700 412600 4752
rect 540520 4700 540572 4752
rect 80244 4632 80296 4684
rect 175556 4632 175608 4684
rect 205088 4632 205140 4684
rect 238944 4632 238996 4684
rect 333796 4632 333848 4684
rect 387064 4632 387116 4684
rect 411168 4632 411220 4684
rect 536932 4632 536984 4684
rect 83832 4564 83884 4616
rect 176752 4564 176804 4616
rect 204168 4564 204220 4616
rect 234620 4564 234672 4616
rect 332508 4564 332560 4616
rect 383568 4564 383620 4616
rect 409788 4564 409840 4616
rect 533436 4564 533488 4616
rect 87328 4496 87380 4548
rect 178040 4496 178092 4548
rect 329748 4496 329800 4548
rect 379980 4496 380032 4548
rect 406936 4496 406988 4548
rect 529848 4496 529900 4548
rect 49332 4428 49384 4480
rect 130384 4428 130436 4480
rect 138480 4428 138532 4480
rect 204260 4428 204312 4480
rect 328276 4428 328328 4480
rect 376392 4428 376444 4480
rect 405648 4428 405700 4480
rect 526260 4428 526312 4480
rect 52828 4360 52880 4412
rect 122104 4360 122156 4412
rect 124220 4360 124272 4412
rect 125968 4360 126020 4412
rect 63592 4292 63644 4344
rect 128820 4292 128872 4344
rect 70676 4224 70728 4276
rect 120724 4224 120776 4276
rect 123484 4224 123536 4276
rect 109960 4156 110012 4208
rect 46940 4088 46992 4140
rect 39764 4020 39816 4072
rect 153200 4088 153252 4140
rect 156328 4088 156380 4140
rect 214012 4360 214064 4412
rect 326988 4360 327040 4412
rect 372804 4360 372856 4412
rect 401508 4360 401560 4412
rect 519084 4360 519136 4412
rect 165620 4292 165672 4344
rect 215576 4292 215628 4344
rect 324136 4292 324188 4344
rect 369216 4292 369268 4344
rect 404268 4292 404320 4344
rect 522672 4292 522724 4344
rect 168288 4224 168340 4276
rect 208492 4224 208544 4276
rect 322572 4224 322624 4276
rect 365720 4224 365772 4276
rect 400036 4224 400088 4276
rect 515588 4224 515640 4276
rect 321376 4156 321428 4208
rect 362132 4156 362184 4208
rect 398748 4156 398800 4208
rect 512000 4156 512052 4208
rect 171784 4088 171836 4140
rect 174544 4088 174596 4140
rect 177764 4088 177816 4140
rect 185676 4088 185728 4140
rect 189632 4088 189684 4140
rect 190368 4088 190420 4140
rect 190828 4088 190880 4140
rect 157340 4020 157392 4072
rect 34980 3952 35032 4004
rect 151912 3952 151964 4004
rect 161112 3952 161164 4004
rect 170404 4020 170456 4072
rect 174176 4020 174228 4072
rect 185584 4020 185636 4072
rect 188436 4020 188488 4072
rect 218152 4020 218204 4072
rect 219256 4020 219308 4072
rect 222936 4020 222988 4072
rect 223488 4020 223540 4072
rect 226524 4088 226576 4140
rect 227628 4088 227680 4140
rect 227720 4088 227772 4140
rect 229008 4088 229060 4140
rect 231308 4088 231360 4140
rect 231768 4088 231820 4140
rect 232504 4088 232556 4140
rect 233148 4088 233200 4140
rect 233700 4088 233752 4140
rect 234528 4088 234580 4140
rect 236000 4088 236052 4140
rect 237196 4088 237248 4140
rect 239588 4088 239640 4140
rect 240048 4088 240100 4140
rect 240784 4088 240836 4140
rect 241428 4088 241480 4140
rect 243176 4088 243228 4140
rect 244188 4088 244240 4140
rect 251456 4088 251508 4140
rect 252468 4088 252520 4140
rect 265808 4088 265860 4140
rect 266268 4088 266320 4140
rect 268108 4088 268160 4140
rect 269764 4088 269816 4140
rect 271696 4088 271748 4140
rect 272524 4088 272576 4140
rect 274088 4088 274140 4140
rect 274548 4088 274600 4140
rect 280068 4088 280120 4140
rect 282460 4088 282512 4140
rect 284944 4088 284996 4140
rect 288348 4088 288400 4140
rect 292396 4088 292448 4140
rect 307392 4088 307444 4140
rect 315304 4088 315356 4140
rect 315856 4088 315908 4140
rect 321468 4088 321520 4140
rect 231952 4020 232004 4072
rect 241980 4020 242032 4072
rect 243544 4020 243596 4072
rect 283564 4020 283616 4072
rect 287152 4020 287204 4072
rect 297916 4020 297968 4072
rect 298008 4020 298060 4072
rect 316960 4020 317012 4072
rect 324228 4020 324280 4072
rect 168196 3952 168248 4004
rect 176016 3952 176068 4004
rect 183744 3952 183796 4004
rect 227812 3952 227864 4004
rect 269304 3952 269356 4004
rect 272156 3952 272208 4004
rect 32680 3884 32732 3936
rect 150624 3884 150676 3936
rect 164700 3884 164752 3936
rect 175924 3884 175976 3936
rect 180156 3884 180208 3936
rect 226432 3884 226484 3936
rect 236644 3884 236696 3936
rect 285588 3884 285640 3936
rect 293132 3952 293184 4004
rect 318064 3952 318116 4004
rect 322848 3952 322900 4004
rect 358084 4088 358136 4140
rect 360936 4088 360988 4140
rect 363604 4088 363656 4140
rect 364524 4088 364576 4140
rect 391756 4088 391808 4140
rect 500132 4088 500184 4140
rect 500224 4088 500276 4140
rect 507124 4088 507176 4140
rect 571432 4088 571484 4140
rect 368020 4020 368072 4072
rect 395988 4020 396040 4072
rect 507216 4020 507268 4072
rect 511264 4020 511316 4072
rect 578608 4020 578660 4072
rect 363328 3952 363380 4004
rect 400128 3952 400180 4004
rect 514392 3952 514444 4004
rect 288256 3884 288308 3936
rect 297916 3884 297968 3936
rect 302148 3884 302200 3936
rect 324044 3884 324096 3936
rect 326344 3884 326396 3936
rect 370412 3884 370464 3936
rect 374644 3884 374696 3936
rect 25504 3816 25556 3868
rect 146392 3816 146444 3868
rect 153936 3816 153988 3868
rect 171508 3816 171560 3868
rect 176568 3816 176620 3868
rect 24308 3748 24360 3800
rect 146300 3748 146352 3800
rect 151544 3748 151596 3800
rect 171692 3748 171744 3800
rect 172980 3748 173032 3800
rect 222384 3816 222436 3868
rect 233424 3816 233476 3868
rect 286968 3816 287020 3868
rect 295524 3816 295576 3868
rect 299388 3816 299440 3868
rect 320456 3816 320508 3868
rect 328368 3816 328420 3868
rect 375196 3816 375248 3868
rect 402888 3884 402940 3936
rect 521476 3884 521528 3936
rect 393044 3816 393096 3868
rect 230572 3748 230624 3800
rect 234804 3748 234856 3800
rect 250444 3748 250496 3800
rect 288072 3748 288124 3800
rect 299112 3748 299164 3800
rect 302056 3748 302108 3800
rect 325240 3748 325292 3800
rect 326160 3748 326212 3800
rect 334624 3748 334676 3800
rect 335912 3748 335964 3800
rect 19524 3680 19576 3732
rect 143540 3680 143592 3732
rect 146852 3680 146904 3732
rect 168288 3680 168340 3732
rect 169392 3680 169444 3732
rect 220820 3680 220872 3732
rect 221740 3680 221792 3732
rect 240692 3680 240744 3732
rect 286876 3680 286928 3732
rect 296720 3680 296772 3732
rect 303528 3680 303580 3732
rect 327632 3680 327684 3732
rect 333888 3680 333940 3732
rect 385868 3748 385920 3800
rect 389824 3748 389876 3800
rect 403716 3748 403768 3800
rect 407028 3816 407080 3868
rect 528652 3816 528704 3868
rect 409512 3748 409564 3800
rect 535736 3748 535788 3800
rect 382372 3680 382424 3732
rect 384304 3680 384356 3732
rect 396632 3680 396684 3732
rect 396724 3680 396776 3732
rect 410892 3680 410944 3732
rect 418160 3680 418212 3732
rect 542912 3680 542964 3732
rect 14832 3612 14884 3664
rect 140780 3612 140832 3664
rect 165896 3612 165948 3664
rect 219624 3612 219676 3664
rect 224132 3612 224184 3664
rect 228916 3612 228968 3664
rect 247684 3612 247736 3664
rect 284208 3612 284260 3664
rect 289544 3612 289596 3664
rect 290924 3612 290976 3664
rect 303804 3612 303856 3664
rect 306288 3612 306340 3664
rect 332416 3612 332468 3664
rect 335268 3612 335320 3664
rect 389456 3612 389508 3664
rect 393964 3612 394016 3664
rect 413192 3612 413244 3664
rect 420184 3612 420236 3664
rect 553584 3612 553636 3664
rect 16028 3544 16080 3596
rect 142344 3544 142396 3596
rect 162308 3544 162360 3596
rect 216864 3544 216916 3596
rect 223580 3544 223632 3596
rect 248604 3544 248656 3596
rect 291108 3544 291160 3596
rect 302608 3544 302660 3596
rect 303436 3544 303488 3596
rect 328828 3544 328880 3596
rect 331128 3544 331180 3596
rect 341616 3544 341668 3596
rect 343088 3544 343140 3596
rect 366916 3544 366968 3596
rect 398104 3544 398156 3596
rect 408316 3544 408368 3596
rect 408500 3544 408552 3596
rect 427636 3544 427688 3596
rect 560760 3544 560812 3596
rect 10048 3476 10100 3528
rect 138020 3476 138072 3528
rect 159916 3476 159968 3528
rect 165620 3476 165672 3528
rect 175372 3476 175424 3528
rect 177304 3476 177356 3528
rect 196808 3476 196860 3528
rect 197268 3476 197320 3528
rect 200396 3476 200448 3528
rect 201408 3476 201460 3528
rect 207480 3476 207532 3528
rect 208308 3476 208360 3528
rect 209872 3476 209924 3528
rect 211068 3476 211120 3528
rect 257436 3476 257488 3528
rect 257988 3476 258040 3528
rect 259828 3476 259880 3528
rect 261484 3476 261536 3528
rect 262220 3476 262272 3528
rect 263508 3476 263560 3528
rect 291016 3476 291068 3528
rect 305000 3476 305052 3528
rect 305644 3476 305696 3528
rect 306288 3476 306340 3528
rect 309048 3476 309100 3528
rect 339500 3476 339552 3528
rect 344928 3476 344980 3528
rect 407304 3476 407356 3528
rect 417884 3476 417936 3528
rect 6460 3408 6512 3460
rect 136916 3408 136968 3460
rect 144460 3408 144512 3460
rect 208584 3408 208636 3460
rect 214564 3408 214616 3460
rect 217048 3408 217100 3460
rect 243636 3408 243688 3460
rect 270500 3408 270552 3460
rect 273352 3408 273404 3460
rect 285496 3408 285548 3460
rect 294328 3408 294380 3460
rect 295248 3408 295300 3460
rect 310980 3408 311032 3460
rect 313188 3408 313240 3460
rect 346676 3408 346728 3460
rect 351828 3408 351880 3460
rect 421564 3476 421616 3528
rect 427820 3476 427872 3528
rect 439412 3476 439464 3528
rect 567844 3476 567896 3528
rect 418344 3408 418396 3460
rect 432328 3408 432380 3460
rect 442172 3408 442224 3460
rect 582196 3408 582248 3460
rect 27896 3340 27948 3392
rect 28908 3340 28960 3392
rect 50528 3340 50580 3392
rect 158904 3340 158956 3392
rect 194416 3340 194468 3392
rect 225328 3340 225380 3392
rect 226248 3340 226300 3392
rect 250352 3340 250404 3392
rect 251088 3340 251140 3392
rect 293868 3340 293920 3392
rect 308588 3340 308640 3392
rect 320088 3340 320140 3392
rect 359740 3340 359792 3392
rect 389088 3340 389140 3392
rect 492956 3340 493008 3392
rect 496084 3340 496136 3392
rect 42156 3272 42208 3324
rect 42708 3272 42760 3324
rect 45744 3272 45796 3324
rect 143724 3272 143776 3324
rect 182548 3272 182600 3324
rect 183468 3272 183520 3324
rect 193220 3272 193272 3324
rect 194508 3272 194560 3324
rect 232136 3272 232188 3324
rect 244372 3272 244424 3324
rect 245476 3272 245528 3324
rect 249156 3272 249208 3324
rect 249708 3272 249760 3324
rect 253848 3272 253900 3324
rect 257344 3272 257396 3324
rect 267004 3272 267056 3324
rect 267648 3272 267700 3324
rect 292488 3272 292540 3324
rect 306196 3272 306248 3324
rect 306288 3272 306340 3324
rect 314568 3272 314620 3324
rect 317328 3272 317380 3324
rect 353760 3272 353812 3324
rect 358176 3272 358228 3324
rect 378784 3272 378836 3324
rect 383476 3272 383528 3324
rect 482284 3272 482336 3324
rect 486424 3272 486476 3324
rect 60004 3204 60056 3256
rect 60648 3204 60700 3256
rect 73804 3204 73856 3256
rect 74264 3204 74316 3256
rect 81440 3204 81492 3256
rect 82728 3204 82780 3256
rect 89720 3204 89772 3256
rect 179880 3204 179932 3256
rect 181352 3204 181404 3256
rect 211068 3204 211120 3256
rect 220544 3204 220596 3256
rect 238024 3204 238076 3256
rect 246764 3204 246816 3256
rect 250536 3204 250588 3256
rect 261024 3204 261076 3256
rect 262128 3204 262180 3256
rect 281448 3204 281500 3256
rect 285956 3204 286008 3256
rect 294604 3204 294656 3256
rect 301412 3204 301464 3256
rect 315856 3204 315908 3256
rect 321652 3204 321704 3256
rect 322204 3204 322256 3256
rect 357348 3204 357400 3256
rect 379428 3204 379480 3256
rect 475108 3204 475160 3256
rect 475384 3204 475436 3256
rect 493324 3272 493376 3324
rect 502984 3272 503036 3324
rect 564348 3340 564400 3392
rect 557172 3272 557224 3324
rect 503628 3204 503680 3256
rect 550088 3204 550140 3256
rect 92112 3068 92164 3120
rect 97264 3136 97316 3188
rect 98000 3136 98052 3188
rect 99288 3136 99340 3188
rect 96896 3068 96948 3120
rect 183560 3136 183612 3188
rect 184848 3136 184900 3188
rect 103980 3068 104032 3120
rect 186596 3068 186648 3120
rect 192024 3136 192076 3188
rect 203892 3136 203944 3188
rect 233884 3136 233936 3188
rect 281356 3136 281408 3188
rect 284760 3136 284812 3188
rect 297364 3136 297416 3188
rect 300308 3136 300360 3188
rect 302884 3136 302936 3188
rect 309784 3136 309836 3188
rect 320824 3136 320876 3188
rect 350264 3136 350316 3188
rect 375288 3136 375340 3188
rect 467932 3136 467984 3188
rect 474004 3136 474056 3188
rect 496544 3136 496596 3188
rect 546500 3136 546552 3188
rect 193864 3068 193916 3120
rect 202696 3068 202748 3120
rect 231124 3068 231176 3120
rect 258632 3068 258684 3120
rect 259368 3068 259420 3120
rect 264612 3068 264664 3120
rect 268384 3068 268436 3120
rect 372528 3068 372580 3120
rect 460848 3068 460900 3120
rect 469864 3068 469916 3120
rect 489368 3068 489420 3120
rect 111156 3000 111208 3052
rect 190736 3000 190788 3052
rect 199200 3000 199252 3052
rect 225604 3000 225656 3052
rect 252652 3000 252704 3052
rect 254584 3000 254636 3052
rect 377404 3000 377456 3052
rect 453672 3000 453724 3052
rect 489184 3000 489236 3052
rect 539324 3068 539376 3120
rect 532240 3000 532292 3052
rect 118240 2932 118292 2984
rect 194784 2932 194836 2984
rect 198004 2932 198056 2984
rect 204168 2932 204220 2984
rect 206284 2932 206336 2984
rect 232412 2932 232464 2984
rect 308404 2932 308456 2984
rect 313372 2932 313424 2984
rect 369124 2932 369176 2984
rect 371608 2932 371660 2984
rect 376024 2932 376076 2984
rect 414480 2932 414532 2984
rect 416044 2932 416096 2984
rect 418160 2932 418212 2984
rect 424324 2932 424376 2984
rect 201500 2864 201552 2916
rect 203800 2864 203852 2916
rect 214656 2864 214708 2916
rect 239404 2864 239456 2916
rect 369400 2864 369452 2916
rect 428740 2864 428792 2916
rect 429844 2864 429896 2916
rect 478144 2932 478196 2984
rect 482192 2932 482244 2984
rect 510804 2932 510856 2984
rect 485780 2864 485832 2916
rect 148048 2796 148100 2848
rect 209964 2796 210016 2848
rect 340788 2796 340840 2848
rect 400220 2796 400272 2848
rect 402244 2796 402296 2848
rect 446588 2796 446640 2848
rect 480904 2796 480956 2848
rect 525064 2864 525116 2916
rect 517888 2796 517940 2848
rect 23112 552 23164 604
rect 23388 552 23440 604
rect 178960 552 179012 604
rect 179328 552 179380 604
rect 272892 552 272944 604
rect 273168 552 273220 604
rect 290096 552 290148 604
rect 290740 552 290792 604
rect 291384 552 291436 604
rect 291936 552 291988 604
rect 318984 552 319036 604
rect 319260 552 319312 604
rect 326436 595 326488 604
rect 326436 561 326445 595
rect 326445 561 326479 595
rect 326479 561 326488 595
rect 326436 552 326488 561
rect 332876 552 332928 604
rect 333612 552 333664 604
rect 336924 552 336976 604
rect 337108 552 337160 604
rect 343916 552 343968 604
rect 344284 552 344336 604
rect 425152 552 425204 604
rect 425336 552 425388 604
rect 456800 552 456852 604
rect 457260 552 457312 604
rect 470600 552 470652 604
rect 471520 552 471572 604
rect 473360 552 473412 604
rect 473912 552 473964 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700398 8156 703520
rect 8116 700392 8168 700398
rect 8116 700334 8168 700340
rect 13084 700392 13136 700398
rect 13084 700334 13136 700340
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 4802 653576 4858 653585
rect 4802 653511 4858 653520
rect 3422 624880 3478 624889
rect 3422 624815 3478 624824
rect 3436 623830 3464 624815
rect 3424 623824 3476 623830
rect 3424 623766 3476 623772
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 610026 3464 610399
rect 3424 610020 3476 610026
rect 3424 609962 3476 609968
rect 4066 596048 4122 596057
rect 4066 595983 4122 595992
rect 4080 594862 4108 595983
rect 4068 594856 4120 594862
rect 4068 594798 4120 594804
rect 3422 567352 3478 567361
rect 3422 567287 3478 567296
rect 3146 553072 3202 553081
rect 3146 553007 3202 553016
rect 3160 552090 3188 553007
rect 3148 552084 3200 552090
rect 3148 552026 3200 552032
rect 3330 495544 3386 495553
rect 3330 495479 3332 495488
rect 3384 495479 3386 495488
rect 3332 495450 3384 495456
rect 3054 452432 3110 452441
rect 3054 452367 3110 452376
rect 3068 451382 3096 452367
rect 3056 451376 3108 451382
rect 3056 451318 3108 451324
rect 2778 366208 2834 366217
rect 2778 366143 2834 366152
rect 2792 365770 2820 366143
rect 2780 365764 2832 365770
rect 2780 365706 2832 365712
rect 2962 337512 3018 337521
rect 2962 337447 3018 337456
rect 2976 336802 3004 337447
rect 2964 336796 3016 336802
rect 2964 336738 3016 336744
rect 3330 294400 3386 294409
rect 3330 294335 3386 294344
rect 3344 294030 3372 294335
rect 3332 294024 3384 294030
rect 3332 293966 3384 293972
rect 2778 265704 2834 265713
rect 2778 265639 2834 265648
rect 2792 264994 2820 265639
rect 2780 264988 2832 264994
rect 2780 264930 2832 264936
rect 3330 251288 3386 251297
rect 3330 251223 3332 251232
rect 3384 251223 3386 251232
rect 3332 251194 3384 251200
rect 3330 237008 3386 237017
rect 3330 236943 3386 236952
rect 2962 222592 3018 222601
rect 2962 222527 3018 222536
rect 2976 222222 3004 222527
rect 2964 222216 3016 222222
rect 2964 222158 3016 222164
rect 2962 208176 3018 208185
rect 2962 208111 3018 208120
rect 2976 207058 3004 208111
rect 2964 207052 3016 207058
rect 2964 206994 3016 207000
rect 3240 200184 3292 200190
rect 3240 200126 3292 200132
rect 2872 180804 2924 180810
rect 2872 180746 2924 180752
rect 2884 179489 2912 180746
rect 2870 179480 2926 179489
rect 2870 179415 2926 179424
rect 3252 165073 3280 200126
rect 3238 165064 3294 165073
rect 3238 164999 3294 165008
rect 3240 156052 3292 156058
rect 3240 155994 3292 156000
rect 3252 150793 3280 155994
rect 3344 154290 3372 236943
rect 3436 201006 3464 567287
rect 3514 538656 3570 538665
rect 3514 538591 3570 538600
rect 3424 201000 3476 201006
rect 3424 200942 3476 200948
rect 3424 197396 3476 197402
rect 3424 197338 3476 197344
rect 3332 154284 3384 154290
rect 3332 154226 3384 154232
rect 3238 150784 3294 150793
rect 3238 150719 3294 150728
rect 3332 136604 3384 136610
rect 3332 136546 3384 136552
rect 3344 136377 3372 136546
rect 3330 136368 3386 136377
rect 3330 136303 3386 136312
rect 3330 122088 3386 122097
rect 3330 122023 3386 122032
rect 3344 120630 3372 122023
rect 3332 120624 3384 120630
rect 3332 120566 3384 120572
rect 2780 93356 2832 93362
rect 2780 93298 2832 93304
rect 2792 93265 2820 93298
rect 2778 93256 2834 93265
rect 2778 93191 2834 93200
rect 3240 80028 3292 80034
rect 3240 79970 3292 79976
rect 3252 78985 3280 79970
rect 3238 78976 3294 78985
rect 3238 78911 3294 78920
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 3436 50153 3464 197338
rect 3528 189038 3556 538591
rect 3606 509960 3662 509969
rect 3606 509895 3662 509904
rect 3620 201074 3648 509895
rect 4066 481128 4122 481137
rect 4066 481063 4122 481072
rect 4080 480690 4108 481063
rect 4068 480684 4120 480690
rect 4068 480626 4120 480632
rect 3698 438016 3754 438025
rect 3698 437951 3754 437960
rect 3608 201068 3660 201074
rect 3608 201010 3660 201016
rect 3606 193896 3662 193905
rect 3606 193831 3662 193840
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3516 156120 3568 156126
rect 3516 156062 3568 156068
rect 3528 107681 3556 156062
rect 3620 155922 3648 193831
rect 3608 155916 3660 155922
rect 3608 155858 3660 155864
rect 3712 150414 3740 437951
rect 4066 423736 4122 423745
rect 4066 423671 4068 423680
rect 4120 423671 4122 423680
rect 4068 423642 4120 423648
rect 3882 395040 3938 395049
rect 3882 394975 3938 394984
rect 3790 380624 3846 380633
rect 3790 380559 3846 380568
rect 3804 151774 3832 380559
rect 3896 201142 3924 394975
rect 3974 323096 4030 323105
rect 3974 323031 4030 323040
rect 3884 201136 3936 201142
rect 3884 201078 3936 201084
rect 3988 152998 4016 323031
rect 4066 308816 4122 308825
rect 4066 308751 4122 308760
rect 4080 307834 4108 308751
rect 4068 307828 4120 307834
rect 4068 307770 4120 307776
rect 4066 280120 4122 280129
rect 4066 280055 4122 280064
rect 4080 153202 4108 280055
rect 4816 186318 4844 653511
rect 4896 594856 4948 594862
rect 4896 594798 4948 594804
rect 4908 187678 4936 594798
rect 4988 480684 5040 480690
rect 4988 480626 5040 480632
rect 5000 188970 5028 480626
rect 5080 423700 5132 423706
rect 5080 423642 5132 423648
rect 5092 190466 5120 423642
rect 5172 365764 5224 365770
rect 5172 365706 5224 365712
rect 5184 191826 5212 365706
rect 5264 307828 5316 307834
rect 5264 307770 5316 307776
rect 5276 193186 5304 307770
rect 5448 264988 5500 264994
rect 5448 264930 5500 264936
rect 5356 196308 5408 196314
rect 5356 196250 5408 196256
rect 5264 193180 5316 193186
rect 5264 193122 5316 193128
rect 5172 191820 5224 191826
rect 5172 191762 5224 191768
rect 5080 190460 5132 190466
rect 5080 190402 5132 190408
rect 4988 188964 5040 188970
rect 4988 188906 5040 188912
rect 4896 187672 4948 187678
rect 4896 187614 4948 187620
rect 4804 186312 4856 186318
rect 4804 186254 4856 186260
rect 4068 153196 4120 153202
rect 4068 153138 4120 153144
rect 3976 152992 4028 152998
rect 3976 152934 4028 152940
rect 3792 151768 3844 151774
rect 3792 151710 3844 151716
rect 3700 150408 3752 150414
rect 3700 150350 3752 150356
rect 3514 107672 3570 107681
rect 3514 107607 3570 107616
rect 5368 93362 5396 196250
rect 5460 193118 5488 264930
rect 5448 193112 5500 193118
rect 5448 193054 5500 193060
rect 13096 184890 13124 700334
rect 24320 699718 24348 703520
rect 40512 700330 40540 703520
rect 40500 700324 40552 700330
rect 40500 700266 40552 700272
rect 72988 699718 73016 703520
rect 89180 700398 89208 703520
rect 105464 700466 105492 703520
rect 133972 701004 134024 701010
rect 133972 700946 134024 700952
rect 133788 700936 133840 700942
rect 133788 700878 133840 700884
rect 132500 700868 132552 700874
rect 132500 700810 132552 700816
rect 131120 700732 131172 700738
rect 131120 700674 131172 700680
rect 105452 700460 105504 700466
rect 105452 700402 105504 700408
rect 89168 700392 89220 700398
rect 89168 700334 89220 700340
rect 126244 700392 126296 700398
rect 126244 700334 126296 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 72424 699712 72476 699718
rect 72424 699654 72476 699660
rect 72976 699712 73028 699718
rect 72976 699654 73028 699660
rect 19984 667956 20036 667962
rect 19984 667898 20036 667904
rect 14464 222216 14516 222222
rect 14464 222158 14516 222164
rect 14476 194478 14504 222158
rect 17224 196104 17276 196110
rect 17224 196046 17276 196052
rect 15844 194608 15896 194614
rect 15844 194550 15896 194556
rect 14464 194472 14516 194478
rect 14464 194414 14516 194420
rect 13084 184884 13136 184890
rect 13084 184826 13136 184832
rect 15856 180810 15884 194550
rect 15844 180804 15896 180810
rect 15844 180746 15896 180752
rect 17236 136610 17264 196046
rect 19996 146266 20024 667898
rect 21364 610020 21416 610026
rect 21364 609962 21416 609968
rect 21376 147626 21404 609962
rect 21364 147620 21416 147626
rect 21364 147562 21416 147568
rect 19984 146260 20036 146266
rect 19984 146202 20036 146208
rect 24780 144702 24808 699654
rect 28264 552084 28316 552090
rect 28264 552026 28316 552032
rect 28276 149054 28304 552026
rect 70308 524476 70360 524482
rect 70308 524418 70360 524424
rect 70216 500268 70268 500274
rect 70216 500210 70268 500216
rect 31024 495508 31076 495514
rect 31024 495450 31076 495456
rect 28264 149048 28316 149054
rect 28264 148990 28316 148996
rect 31036 148986 31064 495450
rect 70124 407856 70176 407862
rect 70124 407798 70176 407804
rect 69940 396772 69992 396778
rect 69940 396714 69992 396720
rect 69664 390584 69716 390590
rect 69664 390526 69716 390532
rect 31024 148980 31076 148986
rect 31024 148922 31076 148928
rect 24768 144696 24820 144702
rect 24768 144638 24820 144644
rect 17224 136604 17276 136610
rect 17224 136546 17276 136552
rect 42708 118652 42760 118658
rect 42708 118594 42760 118600
rect 31668 118312 31720 118318
rect 31668 118254 31720 118260
rect 28908 118244 28960 118250
rect 28908 118186 28960 118192
rect 23388 118176 23440 118182
rect 23388 118118 23440 118124
rect 5356 93356 5408 93362
rect 5356 93298 5408 93304
rect 3422 50144 3478 50153
rect 3422 50079 3478 50088
rect 3424 35896 3476 35902
rect 3422 35864 3424 35873
rect 3476 35864 3478 35873
rect 3422 35799 3478 35808
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 3160 21457 3188 22034
rect 3146 21448 3202 21457
rect 3146 21383 3202 21392
rect 18328 9172 18380 9178
rect 18328 9114 18380 9120
rect 11244 9036 11296 9042
rect 11244 8978 11296 8984
rect 5264 8968 5316 8974
rect 5264 8910 5316 8916
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 1676 7744 1728 7750
rect 1676 7686 1728 7692
rect 572 7608 624 7614
rect 572 7550 624 7556
rect 584 480 612 7550
rect 1688 480 1716 7686
rect 2872 7676 2924 7682
rect 2872 7618 2924 7624
rect 2884 480 2912 7618
rect 3436 7177 3464 8230
rect 4068 7812 4120 7818
rect 4068 7754 4120 7760
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 4080 480 4108 7754
rect 5276 480 5304 8910
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 6460 3460 6512 3466
rect 6460 3402 6512 3408
rect 6472 480 6500 3402
rect 7668 480 7696 7822
rect 8852 6520 8904 6526
rect 8852 6462 8904 6468
rect 8864 480 8892 6462
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 10060 480 10088 3470
rect 11256 480 11284 8978
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 12440 4888 12492 4894
rect 12440 4830 12492 4836
rect 12452 480 12480 4830
rect 13648 480 13676 7890
rect 17224 4820 17276 4826
rect 17224 4762 17276 4768
rect 14832 3664 14884 3670
rect 14832 3606 14884 3612
rect 14844 480 14872 3606
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 16040 480 16068 3538
rect 17236 480 17264 4762
rect 18340 480 18368 9114
rect 20720 9104 20772 9110
rect 20720 9046 20772 9052
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19536 480 19564 3674
rect 20732 480 20760 9046
rect 21916 4956 21968 4962
rect 21916 4898 21968 4904
rect 21928 480 21956 4898
rect 23400 610 23428 118118
rect 26700 5024 26752 5030
rect 26700 4966 26752 4972
rect 25504 3868 25556 3874
rect 25504 3810 25556 3816
rect 24308 3800 24360 3806
rect 24308 3742 24360 3748
rect 23112 604 23164 610
rect 23112 546 23164 552
rect 23388 604 23440 610
rect 23388 546 23440 552
rect 23124 480 23152 546
rect 24320 480 24348 3742
rect 25516 480 25544 3810
rect 26712 480 26740 4966
rect 28920 3398 28948 118186
rect 29092 5092 29144 5098
rect 29092 5034 29144 5040
rect 27896 3392 27948 3398
rect 27896 3334 27948 3340
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 27908 480 27936 3334
rect 29104 480 29132 5034
rect 30286 4856 30342 4865
rect 30286 4791 30342 4800
rect 30300 480 30328 4791
rect 31680 3482 31708 118254
rect 38476 117972 38528 117978
rect 38476 117914 38528 117920
rect 36176 9240 36228 9246
rect 36176 9182 36228 9188
rect 33876 5160 33928 5166
rect 33876 5102 33928 5108
rect 32680 3936 32732 3942
rect 32680 3878 32732 3884
rect 31496 3454 31708 3482
rect 31496 480 31524 3454
rect 32692 480 32720 3878
rect 33888 480 33916 5102
rect 34980 4004 35032 4010
rect 34980 3946 35032 3952
rect 34992 480 35020 3946
rect 36188 480 36216 9182
rect 37372 5228 37424 5234
rect 37372 5170 37424 5176
rect 37384 480 37412 5170
rect 38488 626 38516 117914
rect 40960 9308 41012 9314
rect 40960 9250 41012 9256
rect 39764 4072 39816 4078
rect 39764 4014 39816 4020
rect 38488 598 38608 626
rect 38580 480 38608 598
rect 39776 480 39804 4014
rect 40972 480 41000 9250
rect 42720 3330 42748 118594
rect 69676 118561 69704 390526
rect 69952 385257 69980 396714
rect 70032 395684 70084 395690
rect 70032 395626 70084 395632
rect 69938 385248 69994 385257
rect 69938 385183 69994 385192
rect 70044 362953 70072 395626
rect 70136 370297 70164 407798
rect 70228 377913 70256 500210
rect 70214 377904 70270 377913
rect 70214 377839 70270 377848
rect 70122 370288 70178 370297
rect 70122 370223 70178 370232
rect 70030 362944 70086 362953
rect 70030 362879 70086 362888
rect 70214 355600 70270 355609
rect 70214 355535 70270 355544
rect 70228 342009 70256 355535
rect 70320 348265 70348 524418
rect 71596 407788 71648 407794
rect 71596 407730 71648 407736
rect 71608 392601 71636 407730
rect 71688 398880 71740 398886
rect 71688 398822 71740 398828
rect 71594 392592 71650 392601
rect 71594 392527 71650 392536
rect 71608 390590 71636 392527
rect 71596 390584 71648 390590
rect 71596 390526 71648 390532
rect 71042 377904 71098 377913
rect 71042 377839 71098 377848
rect 70306 348256 70362 348265
rect 70306 348191 70362 348200
rect 70214 342000 70270 342009
rect 70214 341935 70270 341944
rect 69662 118552 69718 118561
rect 69662 118487 69718 118496
rect 56508 118380 56560 118386
rect 56508 118322 56560 118328
rect 55220 9512 55272 9518
rect 55220 9454 55272 9460
rect 51632 9444 51684 9450
rect 51632 9386 51684 9392
rect 43352 9376 43404 9382
rect 43352 9318 43404 9324
rect 42156 3324 42208 3330
rect 42156 3266 42208 3272
rect 42708 3324 42760 3330
rect 42708 3266 42760 3272
rect 42168 480 42196 3266
rect 43364 480 43392 9318
rect 48136 8016 48188 8022
rect 48136 7958 48188 7964
rect 44548 6180 44600 6186
rect 44548 6122 44600 6128
rect 44560 480 44588 6122
rect 46940 4140 46992 4146
rect 46940 4082 46992 4088
rect 45744 3324 45796 3330
rect 45744 3266 45796 3272
rect 45756 480 45784 3266
rect 46952 480 46980 4082
rect 48148 480 48176 7958
rect 49332 4480 49384 4486
rect 49332 4422 49384 4428
rect 49344 480 49372 4422
rect 50528 3392 50580 3398
rect 50528 3334 50580 3340
rect 50540 480 50568 3334
rect 51644 480 51672 9386
rect 54024 6248 54076 6254
rect 54024 6190 54076 6196
rect 52828 4412 52880 4418
rect 52828 4354 52880 4360
rect 52840 480 52868 4354
rect 54036 480 54064 6190
rect 55232 480 55260 9454
rect 56520 626 56548 118322
rect 60648 118040 60700 118046
rect 60648 117982 60700 117988
rect 57612 9648 57664 9654
rect 57612 9590 57664 9596
rect 56428 598 56548 626
rect 56428 480 56456 598
rect 57624 480 57652 9590
rect 58808 9580 58860 9586
rect 58808 9522 58860 9528
rect 58820 480 58848 9522
rect 60660 3262 60688 117982
rect 69676 117978 69704 118487
rect 69664 117972 69716 117978
rect 69664 117914 69716 117920
rect 71056 117434 71084 377839
rect 71594 370288 71650 370297
rect 71594 370223 71650 370232
rect 71502 348256 71558 348265
rect 71502 348191 71558 348200
rect 71516 118454 71544 348191
rect 71504 118448 71556 118454
rect 71504 118390 71556 118396
rect 71608 117881 71636 370223
rect 71700 118114 71728 398822
rect 72436 183530 72464 699654
rect 85396 583364 85448 583370
rect 85396 583306 85448 583312
rect 84106 545864 84162 545873
rect 84106 545799 84162 545808
rect 84014 541512 84070 541521
rect 84014 541447 84070 541456
rect 83922 528728 83978 528737
rect 83922 528663 83978 528672
rect 82818 524920 82874 524929
rect 82818 524855 82874 524864
rect 82832 524482 82860 524855
rect 82820 524476 82872 524482
rect 82820 524418 82872 524424
rect 83936 497554 83964 528663
rect 83924 497548 83976 497554
rect 83924 497490 83976 497496
rect 75828 398132 75880 398138
rect 75828 398074 75880 398080
rect 75840 396250 75868 398074
rect 80796 397860 80848 397866
rect 80796 397802 80848 397808
rect 80808 396250 80836 397802
rect 75532 396222 75868 396250
rect 80500 396222 80836 396250
rect 84028 395894 84056 541447
rect 84016 395888 84068 395894
rect 84016 395830 84068 395836
rect 84120 395758 84148 545799
rect 85302 533080 85358 533089
rect 85302 533015 85358 533024
rect 85316 521286 85344 533015
rect 85408 525609 85436 583306
rect 85580 583296 85632 583302
rect 85580 583238 85632 583244
rect 85488 549908 85540 549914
rect 85488 549850 85540 549856
rect 85394 525600 85450 525609
rect 85394 525535 85450 525544
rect 85304 521280 85356 521286
rect 85304 521222 85356 521228
rect 85500 398886 85528 549850
rect 85592 537781 85620 583238
rect 122748 578604 122800 578610
rect 122748 578546 122800 578552
rect 115388 578468 115440 578474
rect 115388 578410 115440 578416
rect 115204 578332 115256 578338
rect 115204 578274 115256 578280
rect 110328 575544 110380 575550
rect 110328 575486 110380 575492
rect 110340 554810 110368 575486
rect 109408 554804 109460 554810
rect 109408 554746 109460 554752
rect 110328 554804 110380 554810
rect 110328 554746 110380 554752
rect 92112 553988 92164 553994
rect 92112 553930 92164 553936
rect 89168 553920 89220 553926
rect 89168 553862 89220 553868
rect 89180 551820 89208 553862
rect 92124 551820 92152 553930
rect 95056 553784 95108 553790
rect 95056 553726 95108 553732
rect 95068 551820 95096 553726
rect 100760 553716 100812 553722
rect 100760 553658 100812 553664
rect 97816 553512 97868 553518
rect 97816 553454 97868 553460
rect 97828 551820 97856 553454
rect 100772 551820 100800 553658
rect 106464 553648 106516 553654
rect 106464 553590 106516 553596
rect 103704 553580 103756 553586
rect 103704 553522 103756 553528
rect 103716 551820 103744 553522
rect 106476 551820 106504 553590
rect 109420 551820 109448 554746
rect 115112 553852 115164 553858
rect 115112 553794 115164 553800
rect 112352 553444 112404 553450
rect 112352 553386 112404 553392
rect 112364 551820 112392 553386
rect 115124 551820 115152 553794
rect 86406 549944 86462 549953
rect 86406 549879 86408 549888
rect 86460 549879 86462 549888
rect 86408 549850 86460 549856
rect 85578 537772 85634 537781
rect 85578 537707 85634 537716
rect 85592 407794 85620 537707
rect 86604 518770 86632 520132
rect 89364 518906 89392 520132
rect 89352 518900 89404 518906
rect 89352 518842 89404 518848
rect 86592 518764 86644 518770
rect 86592 518706 86644 518712
rect 92308 518226 92336 520132
rect 92296 518220 92348 518226
rect 92296 518162 92348 518168
rect 95252 500274 95280 520132
rect 98012 518430 98040 520132
rect 98000 518424 98052 518430
rect 98000 518366 98052 518372
rect 100956 518294 100984 520132
rect 103532 520118 103914 520146
rect 100944 518288 100996 518294
rect 100944 518230 100996 518236
rect 96528 500948 96580 500954
rect 96528 500890 96580 500896
rect 96540 500274 96568 500890
rect 103532 500886 103560 520118
rect 106660 518362 106688 520132
rect 109604 518838 109632 520132
rect 111812 520118 112562 520146
rect 109592 518832 109644 518838
rect 109592 518774 109644 518780
rect 106648 518356 106700 518362
rect 106648 518298 106700 518304
rect 103520 500880 103572 500886
rect 103520 500822 103572 500828
rect 104808 500880 104860 500886
rect 104808 500822 104860 500828
rect 95240 500268 95292 500274
rect 95240 500210 95292 500216
rect 96528 500268 96580 500274
rect 96528 500210 96580 500216
rect 104820 407862 104848 500822
rect 111708 497956 111760 497962
rect 111708 497898 111760 497904
rect 108948 497616 109000 497622
rect 108948 497558 109000 497564
rect 104808 407856 104860 407862
rect 104808 407798 104860 407804
rect 85580 407788 85632 407794
rect 85580 407730 85632 407736
rect 85488 398880 85540 398886
rect 85488 398822 85540 398828
rect 85500 398750 85528 398822
rect 85488 398744 85540 398750
rect 85488 398686 85540 398692
rect 90272 398744 90324 398750
rect 90272 398686 90324 398692
rect 85948 398200 86000 398206
rect 85948 398142 86000 398148
rect 85960 396250 85988 398142
rect 85652 396222 85988 396250
rect 90284 396250 90312 398686
rect 100668 398268 100720 398274
rect 100668 398210 100720 398216
rect 95884 397588 95936 397594
rect 95884 397530 95936 397536
rect 95896 396250 95924 397530
rect 100680 396250 100708 398210
rect 106004 397656 106056 397662
rect 106004 397598 106056 397604
rect 106016 396250 106044 397598
rect 90284 396222 90620 396250
rect 95588 396222 95924 396250
rect 100556 396222 100708 396250
rect 105708 396222 106044 396250
rect 84108 395752 84160 395758
rect 84108 395694 84160 395700
rect 108960 395690 108988 497558
rect 111720 397730 111748 497898
rect 111812 497486 111840 520118
rect 115216 518838 115244 578274
rect 115296 553988 115348 553994
rect 115296 553930 115348 553936
rect 113824 518832 113876 518838
rect 113824 518774 113876 518780
rect 115204 518832 115256 518838
rect 115204 518774 115256 518780
rect 111800 497480 111852 497486
rect 111800 497422 111852 497428
rect 113836 398274 113864 518774
rect 115308 497962 115336 553930
rect 115400 549914 115428 578410
rect 119344 578400 119396 578406
rect 119344 578342 119396 578348
rect 115940 554804 115992 554810
rect 115940 554746 115992 554752
rect 115388 549908 115440 549914
rect 115388 549850 115440 549856
rect 115296 497956 115348 497962
rect 115296 497898 115348 497904
rect 113824 398268 113876 398274
rect 113824 398210 113876 398216
rect 115952 398138 115980 554746
rect 116032 553444 116084 553450
rect 116032 553386 116084 553392
rect 116044 498098 116072 553386
rect 118054 546544 118110 546553
rect 118054 546479 118110 546488
rect 117318 537432 117374 537441
rect 117318 537367 117374 537376
rect 117332 536858 117360 537367
rect 117320 536852 117372 536858
rect 117320 536794 117372 536800
rect 117318 533352 117374 533361
rect 117318 533287 117374 533296
rect 117332 532778 117360 533287
rect 117320 532772 117372 532778
rect 117320 532714 117372 532720
rect 117964 529916 118016 529922
rect 117964 529858 118016 529864
rect 117976 529553 118004 529858
rect 117962 529544 118018 529553
rect 117962 529479 118018 529488
rect 117318 525192 117374 525201
rect 117318 525127 117374 525136
rect 117332 525094 117360 525127
rect 117320 525088 117372 525094
rect 117320 525030 117372 525036
rect 117318 521112 117374 521121
rect 117318 521047 117374 521056
rect 117332 520946 117360 521047
rect 117320 520940 117372 520946
rect 117320 520882 117372 520888
rect 116032 498092 116084 498098
rect 116032 498034 116084 498040
rect 116044 497622 116072 498034
rect 116032 497616 116084 497622
rect 116032 497558 116084 497564
rect 117320 398812 117372 398818
rect 117320 398754 117372 398760
rect 117332 398206 117360 398754
rect 117320 398200 117372 398206
rect 117320 398142 117372 398148
rect 115940 398132 115992 398138
rect 115940 398074 115992 398080
rect 115848 397792 115900 397798
rect 115848 397734 115900 397740
rect 110972 397724 111024 397730
rect 110972 397666 111024 397672
rect 111708 397724 111760 397730
rect 111708 397666 111760 397672
rect 110984 396250 111012 397666
rect 115860 396250 115888 397734
rect 117976 396778 118004 529479
rect 118068 497622 118096 546479
rect 118238 542464 118294 542473
rect 118238 542399 118294 542408
rect 118252 534070 118280 542399
rect 118240 534064 118292 534070
rect 118240 534006 118292 534012
rect 118516 534064 118568 534070
rect 118516 534006 118568 534012
rect 118528 524550 118556 534006
rect 119356 529922 119384 578342
rect 120724 553784 120776 553790
rect 120724 553726 120776 553732
rect 119344 529916 119396 529922
rect 119344 529858 119396 529864
rect 118516 524544 118568 524550
rect 118516 524486 118568 524492
rect 118424 524408 118476 524414
rect 118424 524350 118476 524356
rect 118436 521665 118464 524350
rect 118238 521656 118294 521665
rect 118238 521591 118294 521600
rect 118422 521656 118478 521665
rect 118422 521591 118478 521600
rect 118252 512038 118280 521591
rect 118240 512032 118292 512038
rect 118240 511974 118292 511980
rect 118516 512032 118568 512038
rect 118516 511974 118568 511980
rect 118528 502382 118556 511974
rect 118332 502376 118384 502382
rect 118516 502376 118568 502382
rect 118384 502324 118464 502330
rect 118332 502318 118464 502324
rect 118516 502318 118568 502324
rect 118344 502302 118464 502318
rect 118436 498137 118464 502302
rect 118422 498128 118478 498137
rect 118422 498063 118478 498072
rect 118056 497616 118108 497622
rect 118056 497558 118108 497564
rect 118436 492674 118464 498063
rect 120736 498030 120764 553726
rect 122760 518974 122788 578546
rect 122748 518968 122800 518974
rect 122748 518910 122800 518916
rect 120724 498024 120776 498030
rect 120724 497966 120776 497972
rect 121368 498024 121420 498030
rect 121368 497966 121420 497972
rect 118436 492658 118556 492674
rect 118332 492652 118384 492658
rect 118436 492652 118568 492658
rect 118436 492646 118516 492652
rect 118332 492594 118384 492600
rect 118516 492594 118568 492600
rect 118344 483041 118372 492594
rect 118330 483032 118386 483041
rect 118330 482967 118386 482976
rect 118606 483032 118662 483041
rect 118606 482967 118662 482976
rect 118620 476082 118648 482967
rect 118436 476054 118648 476082
rect 118436 466546 118464 476054
rect 118424 466540 118476 466546
rect 118424 466482 118476 466488
rect 118332 466404 118384 466410
rect 118332 466346 118384 466352
rect 118344 463690 118372 466346
rect 118056 463684 118108 463690
rect 118056 463626 118108 463632
rect 118332 463684 118384 463690
rect 118332 463626 118384 463632
rect 118068 454073 118096 463626
rect 118054 454064 118110 454073
rect 118054 453999 118110 454008
rect 118238 454064 118294 454073
rect 118238 453999 118294 454008
rect 118252 447166 118280 453999
rect 118240 447160 118292 447166
rect 118240 447102 118292 447108
rect 118332 447092 118384 447098
rect 118332 447034 118384 447040
rect 118344 444378 118372 447034
rect 118056 444372 118108 444378
rect 118056 444314 118108 444320
rect 118332 444372 118384 444378
rect 118332 444314 118384 444320
rect 118068 434761 118096 444314
rect 118054 434752 118110 434761
rect 118054 434687 118110 434696
rect 118238 434752 118294 434761
rect 118238 434687 118294 434696
rect 118252 427854 118280 434687
rect 118240 427848 118292 427854
rect 118240 427790 118292 427796
rect 118332 427780 118384 427786
rect 118332 427722 118384 427728
rect 118344 418146 118372 427722
rect 118344 418118 118464 418146
rect 118436 415410 118464 418118
rect 118424 415404 118476 415410
rect 118424 415346 118476 415352
rect 118516 405748 118568 405754
rect 118516 405690 118568 405696
rect 118528 398834 118556 405690
rect 121380 398886 121408 497966
rect 125876 497480 125928 497486
rect 125876 497422 125928 497428
rect 120908 398880 120960 398886
rect 118528 398818 118648 398834
rect 120908 398822 120960 398828
rect 121368 398880 121420 398886
rect 121368 398822 121420 398828
rect 125692 398880 125744 398886
rect 125692 398822 125744 398828
rect 118528 398812 118660 398818
rect 118528 398806 118608 398812
rect 118608 398754 118660 398760
rect 118620 398723 118648 398754
rect 117964 396772 118016 396778
rect 117964 396714 118016 396720
rect 120920 396250 120948 398822
rect 125600 397520 125652 397526
rect 125600 397462 125652 397468
rect 125612 396250 125640 397462
rect 110676 396222 111012 396250
rect 115644 396222 115888 396250
rect 120612 396222 120948 396250
rect 125580 396222 125640 396250
rect 108948 395684 109000 395690
rect 108948 395626 109000 395632
rect 111708 340264 111760 340270
rect 111708 340206 111760 340212
rect 110328 340196 110380 340202
rect 110328 340138 110380 340144
rect 72588 340054 72924 340082
rect 77556 340054 77892 340082
rect 82524 340054 82768 340082
rect 87492 340054 87828 340082
rect 92460 340054 92796 340082
rect 97612 340054 97948 340082
rect 102580 340054 102916 340082
rect 107548 340054 107608 340082
rect 72896 337618 72924 340054
rect 72884 337612 72936 337618
rect 72884 337554 72936 337560
rect 77864 337482 77892 340054
rect 77852 337476 77904 337482
rect 77852 337418 77904 337424
rect 82740 336734 82768 340054
rect 87800 337414 87828 340054
rect 92768 337754 92796 340054
rect 97920 338026 97948 340054
rect 97908 338020 97960 338026
rect 97908 337962 97960 337968
rect 92756 337748 92808 337754
rect 92756 337690 92808 337696
rect 93768 337748 93820 337754
rect 93768 337690 93820 337696
rect 87788 337408 87840 337414
rect 87788 337350 87840 337356
rect 82728 336728 82780 336734
rect 82728 336670 82780 336676
rect 72424 183524 72476 183530
rect 72424 183466 72476 183472
rect 82740 118522 82768 336670
rect 93780 202162 93808 337690
rect 93768 202156 93820 202162
rect 93768 202098 93820 202104
rect 97920 118590 97948 337962
rect 102888 337754 102916 340054
rect 107580 338094 107608 340054
rect 107568 338088 107620 338094
rect 107568 338030 107620 338036
rect 102876 337748 102928 337754
rect 102876 337690 102928 337696
rect 103428 337748 103480 337754
rect 103428 337690 103480 337696
rect 99288 337476 99340 337482
rect 99288 337418 99340 337424
rect 99300 118697 99328 337418
rect 103440 202230 103468 337690
rect 103428 202224 103480 202230
rect 103428 202166 103480 202172
rect 99286 118688 99342 118697
rect 99286 118623 99342 118632
rect 97908 118584 97960 118590
rect 97908 118526 97960 118532
rect 82728 118516 82780 118522
rect 82728 118458 82780 118464
rect 71688 118108 71740 118114
rect 71688 118050 71740 118056
rect 73804 118108 73856 118114
rect 73804 118050 73856 118056
rect 73988 118108 74040 118114
rect 73988 118050 74040 118056
rect 71594 117872 71650 117881
rect 71594 117807 71650 117816
rect 67548 117428 67600 117434
rect 67548 117370 67600 117376
rect 71044 117428 71096 117434
rect 71044 117370 71096 117376
rect 64788 8900 64840 8906
rect 64788 8842 64840 8848
rect 61200 6316 61252 6322
rect 61200 6258 61252 6264
rect 60004 3256 60056 3262
rect 60004 3198 60056 3204
rect 60648 3256 60700 3262
rect 60648 3198 60700 3204
rect 60016 480 60044 3198
rect 61212 480 61240 6258
rect 62396 5296 62448 5302
rect 62396 5238 62448 5244
rect 62408 480 62436 5238
rect 63592 4344 63644 4350
rect 63592 4286 63644 4292
rect 63604 480 63632 4286
rect 64800 480 64828 8842
rect 65984 5364 66036 5370
rect 65984 5306 66036 5312
rect 65996 480 66024 5306
rect 67560 3482 67588 117370
rect 71872 8832 71924 8838
rect 71872 8774 71924 8780
rect 68284 6384 68336 6390
rect 68284 6326 68336 6332
rect 67192 3454 67588 3482
rect 67192 480 67220 3454
rect 68296 480 68324 6326
rect 69480 5432 69532 5438
rect 69480 5374 69532 5380
rect 69492 480 69520 5374
rect 70676 4276 70728 4282
rect 70676 4218 70728 4224
rect 70688 480 70716 4218
rect 71884 480 71912 8774
rect 73068 5500 73120 5506
rect 73068 5442 73120 5448
rect 73080 480 73108 5442
rect 73816 3262 73844 118050
rect 74000 117978 74028 118050
rect 82740 118046 82768 118458
rect 88340 118448 88392 118454
rect 88340 118390 88392 118396
rect 88352 118046 88380 118390
rect 82728 118040 82780 118046
rect 82728 117982 82780 117988
rect 88340 118040 88392 118046
rect 88340 117982 88392 117988
rect 73988 117972 74040 117978
rect 73988 117914 74040 117920
rect 79966 117872 80022 117881
rect 79966 117807 80022 117816
rect 82728 117836 82780 117842
rect 79980 117722 80008 117807
rect 82728 117778 82780 117784
rect 80150 117736 80206 117745
rect 79980 117694 80150 117722
rect 80150 117671 80206 117680
rect 79048 8764 79100 8770
rect 79048 8706 79100 8712
rect 77852 7336 77904 7342
rect 77852 7278 77904 7284
rect 75460 6452 75512 6458
rect 75460 6394 75512 6400
rect 73804 3256 73856 3262
rect 73804 3198 73856 3204
rect 74264 3256 74316 3262
rect 74264 3198 74316 3204
rect 74276 480 74304 3198
rect 75472 480 75500 6394
rect 76656 4752 76708 4758
rect 76656 4694 76708 4700
rect 76668 480 76696 4694
rect 77864 480 77892 7278
rect 79060 480 79088 8706
rect 82636 6588 82688 6594
rect 82636 6530 82688 6536
rect 80244 4684 80296 4690
rect 80244 4626 80296 4632
rect 80256 480 80284 4626
rect 81440 3256 81492 3262
rect 81440 3198 81492 3204
rect 81452 480 81480 3198
rect 82648 480 82676 6530
rect 82740 3262 82768 117778
rect 84936 7200 84988 7206
rect 84936 7142 84988 7148
rect 83832 4616 83884 4622
rect 83832 4558 83884 4564
rect 82728 3256 82780 3262
rect 82728 3198 82780 3204
rect 83844 480 83872 4558
rect 84948 480 84976 7142
rect 86132 6656 86184 6662
rect 86132 6598 86184 6604
rect 86144 480 86172 6598
rect 87328 4548 87380 4554
rect 87328 4490 87380 4496
rect 87340 480 87368 4490
rect 88352 3482 88380 117982
rect 89810 117872 89866 117881
rect 89640 117830 89810 117858
rect 89640 117745 89668 117830
rect 89810 117807 89866 117816
rect 89626 117736 89682 117745
rect 89626 117671 89682 117680
rect 97920 117366 97948 118526
rect 99196 117904 99248 117910
rect 99194 117872 99196 117881
rect 99248 117872 99250 117881
rect 99194 117807 99250 117816
rect 97264 117360 97316 117366
rect 97264 117302 97316 117308
rect 97908 117360 97960 117366
rect 99300 117337 99328 118623
rect 107580 118318 107608 338030
rect 110340 118425 110368 340138
rect 110326 118416 110382 118425
rect 110326 118351 110382 118360
rect 107568 118312 107620 118318
rect 107568 118254 107620 118260
rect 109040 118312 109092 118318
rect 109040 118254 109092 118260
rect 107580 117910 107608 118254
rect 109052 117978 109080 118254
rect 110340 118182 110368 118351
rect 111720 118250 111748 340206
rect 112516 340054 112852 340082
rect 117668 340054 118004 340082
rect 122636 340054 122788 340082
rect 112824 337958 112852 340054
rect 112812 337952 112864 337958
rect 112812 337894 112864 337900
rect 113088 337952 113140 337958
rect 113088 337894 113140 337900
rect 113100 118318 113128 337894
rect 117976 337550 118004 340054
rect 122760 337890 122788 340054
rect 122748 337884 122800 337890
rect 122748 337826 122800 337832
rect 117964 337544 118016 337550
rect 117964 337486 118016 337492
rect 113088 118312 113140 118318
rect 113088 118254 113140 118260
rect 111708 118244 111760 118250
rect 111708 118186 111760 118192
rect 110328 118176 110380 118182
rect 110328 118118 110380 118124
rect 109040 117972 109092 117978
rect 109040 117914 109092 117920
rect 101220 117904 101272 117910
rect 101218 117872 101220 117881
rect 107568 117904 107620 117910
rect 101272 117872 101274 117881
rect 101218 117807 101274 117816
rect 103518 117872 103574 117881
rect 107568 117846 107620 117852
rect 103518 117807 103574 117816
rect 97908 117302 97960 117308
rect 97998 117328 98054 117337
rect 95700 7132 95752 7138
rect 95700 7074 95752 7080
rect 94504 6860 94556 6866
rect 94504 6802 94556 6808
rect 93308 6792 93360 6798
rect 93308 6734 93360 6740
rect 90916 6724 90968 6730
rect 90916 6666 90968 6672
rect 88352 3454 88564 3482
rect 88536 480 88564 3454
rect 89720 3256 89772 3262
rect 89720 3198 89772 3204
rect 89732 480 89760 3198
rect 90928 480 90956 6666
rect 92112 3120 92164 3126
rect 92112 3062 92164 3068
rect 92124 480 92152 3062
rect 93320 480 93348 6734
rect 94516 480 94544 6802
rect 95712 480 95740 7074
rect 97276 3194 97304 117302
rect 97998 117263 98054 117272
rect 99286 117328 99342 117337
rect 99286 117263 99342 117272
rect 98012 3194 98040 117263
rect 100484 8084 100536 8090
rect 100484 8026 100536 8032
rect 98092 6044 98144 6050
rect 98092 5986 98144 5992
rect 97264 3188 97316 3194
rect 97264 3130 97316 3136
rect 98000 3188 98052 3194
rect 98000 3130 98052 3136
rect 96896 3120 96948 3126
rect 96896 3062 96948 3068
rect 96908 480 96936 3062
rect 98104 480 98132 5986
rect 99288 3188 99340 3194
rect 99288 3130 99340 3136
rect 99300 480 99328 3130
rect 100496 480 100524 8026
rect 103532 6526 103560 117807
rect 104990 117736 105046 117745
rect 104990 117671 104992 117680
rect 105044 117671 105046 117680
rect 104992 117642 105044 117648
rect 111720 117366 111748 118186
rect 113100 117842 113128 118254
rect 115202 117872 115258 117881
rect 113088 117836 113140 117842
rect 122760 117842 122788 337826
rect 124128 337544 124180 337550
rect 124128 337486 124180 337492
rect 124140 118454 124168 337486
rect 124220 154420 124272 154426
rect 124220 154362 124272 154368
rect 124232 154057 124260 154362
rect 124218 154048 124274 154057
rect 124218 153983 124274 153992
rect 124128 118448 124180 118454
rect 124128 118390 124180 118396
rect 122838 117872 122894 117881
rect 115202 117807 115258 117816
rect 122748 117836 122800 117842
rect 113088 117778 113140 117784
rect 115216 117706 115244 117807
rect 122838 117807 122894 117816
rect 122748 117778 122800 117784
rect 115204 117700 115256 117706
rect 115204 117642 115256 117648
rect 120724 117564 120776 117570
rect 120724 117506 120776 117512
rect 111708 117360 111760 117366
rect 111708 117302 111760 117308
rect 120632 8696 120684 8702
rect 120632 8638 120684 8644
rect 106372 8628 106424 8634
rect 106372 8570 106424 8576
rect 103520 6520 103572 6526
rect 103520 6462 103572 6468
rect 105176 6520 105228 6526
rect 105176 6462 105228 6468
rect 102782 6216 102838 6225
rect 102782 6151 102838 6160
rect 101588 6112 101640 6118
rect 101588 6054 101640 6060
rect 101600 480 101628 6054
rect 102796 480 102824 6151
rect 103980 3120 104032 3126
rect 103980 3062 104032 3068
rect 103992 480 104020 3062
rect 105188 480 105216 6462
rect 106384 480 106412 8570
rect 114744 8220 114796 8226
rect 114744 8162 114796 8168
rect 107568 8152 107620 8158
rect 107568 8094 107620 8100
rect 107580 480 107608 8094
rect 108764 5976 108816 5982
rect 108764 5918 108816 5924
rect 108776 480 108804 5918
rect 112352 5908 112404 5914
rect 112352 5850 112404 5856
rect 109960 4208 110012 4214
rect 109960 4150 110012 4156
rect 109972 480 110000 4150
rect 111156 3052 111208 3058
rect 111156 2994 111208 3000
rect 111168 480 111196 2994
rect 112364 480 112392 5850
rect 113548 5840 113600 5846
rect 113548 5782 113600 5788
rect 113560 480 113588 5782
rect 114756 480 114784 8162
rect 117136 7268 117188 7274
rect 117136 7210 117188 7216
rect 115940 5772 115992 5778
rect 115940 5714 115992 5720
rect 115952 480 115980 5714
rect 117148 480 117176 7210
rect 119436 5704 119488 5710
rect 119436 5646 119488 5652
rect 118240 2984 118292 2990
rect 118240 2926 118292 2932
rect 118252 480 118280 2926
rect 119448 480 119476 5646
rect 120644 480 120672 8638
rect 120736 4282 120764 117506
rect 122760 117502 122788 117778
rect 122104 117496 122156 117502
rect 122104 117438 122156 117444
rect 122748 117496 122800 117502
rect 122748 117438 122800 117444
rect 121828 7540 121880 7546
rect 121828 7482 121880 7488
rect 120724 4276 120776 4282
rect 120724 4218 120776 4224
rect 121840 480 121868 7482
rect 122116 4418 122144 117438
rect 122852 117298 122880 117807
rect 124140 117502 124168 118390
rect 125704 118114 125732 398822
rect 125784 395684 125836 395690
rect 125784 395626 125836 395632
rect 125796 118386 125824 395626
rect 125888 336734 125916 497422
rect 126152 397860 126204 397866
rect 126152 397802 126204 397808
rect 126164 383722 126192 397802
rect 126152 383716 126204 383722
rect 126152 383658 126204 383664
rect 126152 374060 126204 374066
rect 126152 374002 126204 374008
rect 126164 364410 126192 374002
rect 126152 364404 126204 364410
rect 126152 364346 126204 364352
rect 126152 354748 126204 354754
rect 126152 354690 126204 354696
rect 126164 345098 126192 354690
rect 126152 345092 126204 345098
rect 126152 345034 126204 345040
rect 125876 336728 125928 336734
rect 125876 336670 125928 336676
rect 126152 335368 126204 335374
rect 126152 335310 126204 335316
rect 126164 325718 126192 335310
rect 126152 325712 126204 325718
rect 126152 325654 126204 325660
rect 126152 316056 126204 316062
rect 126152 315998 126204 316004
rect 126164 296750 126192 315998
rect 126152 296744 126204 296750
rect 126152 296686 126204 296692
rect 126060 292528 126112 292534
rect 126060 292470 126112 292476
rect 126072 282826 126100 292470
rect 126072 282798 126192 282826
rect 126164 280158 126192 282798
rect 126152 280152 126204 280158
rect 126152 280094 126204 280100
rect 126060 270564 126112 270570
rect 126060 270506 126112 270512
rect 126072 263514 126100 270506
rect 126072 263486 126192 263514
rect 126164 260846 126192 263486
rect 126152 260840 126204 260846
rect 126152 260782 126204 260788
rect 126060 251320 126112 251326
rect 126060 251262 126112 251268
rect 126072 244202 126100 251262
rect 126072 244174 126192 244202
rect 126164 234666 126192 244174
rect 126152 234660 126204 234666
rect 126152 234602 126204 234608
rect 126152 224936 126204 224942
rect 126152 224878 126204 224884
rect 126164 215370 126192 224878
rect 126072 215342 126192 215370
rect 126072 202910 126100 215342
rect 126060 202904 126112 202910
rect 126060 202846 126112 202852
rect 126256 144430 126284 700334
rect 129280 583500 129332 583506
rect 129280 583442 129332 583448
rect 126336 583432 126388 583438
rect 126336 583374 126388 583380
rect 126348 397866 126376 583374
rect 129004 578808 129056 578814
rect 129004 578750 129056 578756
rect 128360 553852 128412 553858
rect 128360 553794 128412 553800
rect 127716 518832 127768 518838
rect 127716 518774 127768 518780
rect 126980 518220 127032 518226
rect 126980 518162 127032 518168
rect 126336 397860 126388 397866
rect 126336 397802 126388 397808
rect 126428 397792 126480 397798
rect 126428 397734 126480 397740
rect 126336 383716 126388 383722
rect 126336 383658 126388 383664
rect 126348 374134 126376 383658
rect 126336 374128 126388 374134
rect 126336 374070 126388 374076
rect 126336 364404 126388 364410
rect 126336 364346 126388 364352
rect 126348 354822 126376 364346
rect 126336 354816 126388 354822
rect 126336 354758 126388 354764
rect 126336 345092 126388 345098
rect 126336 345034 126388 345040
rect 126348 335374 126376 345034
rect 126336 335368 126388 335374
rect 126336 335310 126388 335316
rect 126336 325712 126388 325718
rect 126336 325654 126388 325660
rect 126348 316062 126376 325654
rect 126336 316056 126388 316062
rect 126336 315998 126388 316004
rect 126336 296744 126388 296750
rect 126336 296686 126388 296692
rect 126348 292534 126376 296686
rect 126336 292528 126388 292534
rect 126336 292470 126388 292476
rect 126336 234660 126388 234666
rect 126336 234602 126388 234608
rect 126348 224942 126376 234602
rect 126336 224936 126388 224942
rect 126336 224878 126388 224884
rect 126440 205698 126468 397734
rect 126520 396772 126572 396778
rect 126520 396714 126572 396720
rect 126532 384334 126560 396714
rect 126520 384328 126572 384334
rect 126520 384270 126572 384276
rect 126992 338026 127020 518162
rect 127072 497548 127124 497554
rect 127072 497490 127124 497496
rect 126980 338020 127032 338026
rect 126980 337962 127032 337968
rect 127084 337958 127112 497490
rect 127164 398132 127216 398138
rect 127164 398074 127216 398080
rect 127176 340814 127204 398074
rect 127256 397724 127308 397730
rect 127256 397666 127308 397672
rect 127268 340882 127296 397666
rect 127624 397656 127676 397662
rect 127624 397598 127676 397604
rect 127256 340876 127308 340882
rect 127256 340818 127308 340824
rect 127164 340808 127216 340814
rect 127164 340750 127216 340756
rect 127176 340202 127204 340750
rect 127268 340270 127296 340818
rect 127256 340264 127308 340270
rect 127256 340206 127308 340212
rect 127164 340196 127216 340202
rect 127164 340138 127216 340144
rect 127072 337952 127124 337958
rect 127072 337894 127124 337900
rect 126428 205692 126480 205698
rect 126428 205634 126480 205640
rect 126428 205556 126480 205562
rect 126428 205498 126480 205504
rect 126440 201618 126468 205498
rect 126612 202904 126664 202910
rect 126612 202846 126664 202852
rect 126428 201612 126480 201618
rect 126428 201554 126480 201560
rect 126624 201498 126652 202846
rect 127636 201550 127664 397598
rect 127728 340746 127756 518774
rect 128372 358329 128400 553794
rect 128912 521688 128964 521694
rect 128912 521630 128964 521636
rect 128452 520940 128504 520946
rect 128452 520882 128504 520888
rect 128464 373289 128492 520882
rect 128924 514706 128952 521630
rect 129016 520946 129044 578750
rect 129188 578264 129240 578270
rect 129188 578206 129240 578212
rect 129096 553716 129148 553722
rect 129096 553658 129148 553664
rect 129004 520940 129056 520946
rect 129004 520882 129056 520888
rect 128740 514678 128952 514706
rect 128740 512009 128768 514678
rect 128542 512000 128598 512009
rect 128542 511935 128598 511944
rect 128726 512000 128782 512009
rect 128726 511935 128782 511944
rect 128556 502382 128584 511935
rect 128544 502376 128596 502382
rect 128544 502318 128596 502324
rect 128820 502376 128872 502382
rect 128820 502318 128872 502324
rect 128832 495394 128860 502318
rect 129108 498166 129136 553658
rect 129200 525094 129228 578206
rect 129292 553858 129320 583442
rect 129646 582448 129702 582457
rect 129646 582383 129702 582392
rect 129556 563100 129608 563106
rect 129556 563042 129608 563048
rect 129280 553852 129332 553858
rect 129280 553794 129332 553800
rect 129188 525088 129240 525094
rect 129188 525030 129240 525036
rect 129200 521694 129228 525030
rect 129188 521688 129240 521694
rect 129188 521630 129240 521636
rect 129096 498160 129148 498166
rect 129096 498102 129148 498108
rect 128740 495366 128860 495394
rect 128740 492658 128768 495366
rect 128544 492652 128596 492658
rect 128544 492594 128596 492600
rect 128728 492652 128780 492658
rect 128728 492594 128780 492600
rect 128556 483041 128584 492594
rect 128542 483032 128598 483041
rect 128542 482967 128598 482976
rect 128818 483032 128874 483041
rect 128818 482967 128874 482976
rect 128832 476082 128860 482967
rect 128740 476054 128860 476082
rect 128740 468466 128768 476054
rect 128556 468438 128768 468466
rect 128556 463729 128584 468438
rect 128542 463720 128598 463729
rect 128542 463655 128598 463664
rect 128818 463720 128874 463729
rect 128818 463655 128874 463664
rect 128832 456770 128860 463655
rect 128740 456742 128860 456770
rect 128740 449154 128768 456742
rect 128556 449126 128768 449154
rect 128556 444417 128584 449126
rect 128542 444408 128598 444417
rect 128542 444343 128598 444352
rect 128818 444408 128874 444417
rect 128818 444343 128874 444352
rect 128832 437458 128860 444343
rect 128740 437430 128860 437458
rect 128740 429842 128768 437430
rect 128556 429814 128768 429842
rect 128556 425105 128584 429814
rect 128542 425096 128598 425105
rect 128542 425031 128598 425040
rect 128818 425096 128874 425105
rect 128818 425031 128874 425040
rect 128832 418146 128860 425031
rect 128648 418118 128860 418146
rect 128648 415410 128676 418118
rect 128636 415404 128688 415410
rect 128636 415346 128688 415352
rect 128544 405748 128596 405754
rect 128544 405690 128596 405696
rect 128556 404326 128584 405690
rect 128544 404320 128596 404326
rect 128544 404262 128596 404268
rect 128636 394732 128688 394738
rect 128636 394674 128688 394680
rect 128648 394618 128676 394674
rect 128648 394590 128768 394618
rect 128740 388521 128768 394590
rect 128726 388512 128782 388521
rect 128726 388447 128728 388456
rect 128780 388447 128782 388456
rect 128728 388418 128780 388424
rect 128740 388387 128768 388418
rect 129108 380633 129136 498102
rect 129464 398268 129516 398274
rect 129464 398210 129516 398216
rect 129476 397458 129504 398210
rect 129464 397452 129516 397458
rect 129464 397394 129516 397400
rect 129094 380624 129150 380633
rect 129094 380559 129150 380568
rect 128912 376780 128964 376786
rect 128912 376722 128964 376728
rect 128450 373280 128506 373289
rect 128450 373215 128506 373224
rect 128924 369866 128952 376722
rect 128924 369838 129044 369866
rect 129016 360210 129044 369838
rect 128832 360182 129044 360210
rect 128832 360074 128860 360182
rect 128832 360046 128952 360074
rect 128358 358320 128414 358329
rect 128358 358255 128414 358264
rect 128924 341034 128952 360046
rect 129004 351212 129056 351218
rect 129004 351154 129056 351160
rect 129016 350985 129044 351154
rect 129002 350976 129058 350985
rect 129002 350911 129058 350920
rect 129002 343632 129058 343641
rect 129002 343567 129058 343576
rect 129016 342922 129044 343567
rect 129004 342916 129056 342922
rect 129004 342858 129056 342864
rect 128924 341006 129044 341034
rect 127716 340740 127768 340746
rect 127716 340682 127768 340688
rect 127728 337890 127756 340682
rect 129016 338162 129044 341006
rect 128912 338156 128964 338162
rect 128912 338098 128964 338104
rect 129004 338156 129056 338162
rect 129004 338098 129056 338104
rect 127716 337884 127768 337890
rect 127716 337826 127768 337832
rect 128268 337408 128320 337414
rect 128268 337350 128320 337356
rect 126440 201470 126652 201498
rect 127624 201544 127676 201550
rect 127624 201486 127676 201492
rect 126440 195974 126468 201470
rect 126428 195968 126480 195974
rect 126428 195910 126480 195916
rect 126612 195968 126664 195974
rect 126612 195910 126664 195916
rect 126624 191808 126652 195910
rect 126624 191780 126836 191808
rect 126808 182209 126836 191780
rect 126518 182200 126574 182209
rect 126518 182135 126574 182144
rect 126794 182200 126850 182209
rect 126794 182135 126850 182144
rect 126532 176746 126560 182135
rect 126440 176718 126560 176746
rect 126440 176662 126468 176718
rect 126428 176656 126480 176662
rect 126428 176598 126480 176604
rect 126612 176656 126664 176662
rect 126612 176598 126664 176604
rect 126624 161498 126652 176598
rect 126520 161492 126572 161498
rect 126520 161434 126572 161440
rect 126612 161492 126664 161498
rect 126612 161434 126664 161440
rect 126532 157570 126560 161434
rect 126440 157542 126560 157570
rect 126440 153241 126468 157542
rect 126426 153232 126482 153241
rect 126426 153167 126482 153176
rect 126702 153096 126758 153105
rect 126702 153031 126758 153040
rect 126244 144424 126296 144430
rect 126244 144366 126296 144372
rect 126716 143585 126744 153031
rect 128176 144764 128228 144770
rect 128176 144706 128228 144712
rect 128188 144537 128216 144706
rect 128174 144528 128230 144537
rect 128174 144463 128230 144472
rect 126518 143576 126574 143585
rect 126518 143511 126574 143520
rect 126702 143576 126758 143585
rect 126702 143511 126758 143520
rect 126532 138666 126560 143511
rect 126440 138638 126560 138666
rect 126440 124166 126468 138638
rect 126060 124160 126112 124166
rect 126060 124102 126112 124108
rect 126428 124160 126480 124166
rect 126428 124102 126480 124108
rect 125784 118380 125836 118386
rect 125784 118322 125836 118328
rect 125692 118108 125744 118114
rect 125692 118050 125744 118056
rect 125704 117570 125732 118050
rect 125796 117774 125824 118322
rect 125784 117768 125836 117774
rect 125784 117710 125836 117716
rect 126072 117609 126100 124102
rect 128280 118289 128308 337350
rect 128924 331242 128952 338098
rect 128924 331214 129044 331242
rect 129016 328438 129044 331214
rect 129004 328432 129056 328438
rect 129004 328374 129056 328380
rect 128820 318912 128872 318918
rect 128872 318860 128952 318866
rect 128820 318854 128952 318860
rect 128832 318838 128952 318854
rect 128924 317422 128952 318838
rect 128912 317416 128964 317422
rect 128912 317358 128964 317364
rect 128636 307828 128688 307834
rect 128636 307770 128688 307776
rect 128648 302122 128676 307770
rect 128636 302116 128688 302122
rect 128636 302058 128688 302064
rect 128912 302116 128964 302122
rect 128912 302058 128964 302064
rect 128924 299441 128952 302058
rect 128910 299432 128966 299441
rect 128910 299367 128966 299376
rect 128818 289912 128874 289921
rect 128818 289847 128874 289856
rect 128832 289814 128860 289847
rect 128820 289808 128872 289814
rect 128820 289750 128872 289756
rect 128912 280220 128964 280226
rect 128912 280162 128964 280168
rect 128924 280129 128952 280162
rect 128910 280120 128966 280129
rect 128910 280055 128966 280064
rect 129002 279984 129058 279993
rect 129002 279919 129058 279928
rect 129016 270586 129044 279919
rect 128924 270558 129044 270586
rect 128924 263634 128952 270558
rect 128912 263628 128964 263634
rect 128912 263570 128964 263576
rect 128912 260908 128964 260914
rect 128912 260850 128964 260856
rect 128924 260778 128952 260850
rect 128728 260772 128780 260778
rect 128728 260714 128780 260720
rect 128912 260772 128964 260778
rect 128912 260714 128964 260720
rect 128740 253892 128768 260714
rect 128740 253864 128860 253892
rect 128832 244254 128860 253864
rect 128820 244248 128872 244254
rect 128820 244190 128872 244196
rect 129004 244248 129056 244254
rect 129004 244190 129056 244196
rect 129016 236774 129044 244190
rect 129004 236768 129056 236774
rect 129004 236710 129056 236716
rect 129004 231940 129056 231946
rect 129004 231882 129056 231888
rect 129016 222222 129044 231882
rect 128636 222216 128688 222222
rect 128636 222158 128688 222164
rect 129004 222216 129056 222222
rect 129004 222158 129056 222164
rect 128648 215218 128676 222158
rect 128636 215212 128688 215218
rect 128636 215154 128688 215160
rect 129004 215212 129056 215218
rect 129004 215154 129056 215160
rect 129016 202978 129044 215154
rect 129004 202972 129056 202978
rect 129004 202914 129056 202920
rect 128912 202836 128964 202842
rect 128912 202778 128964 202784
rect 128924 200122 128952 202778
rect 128544 200116 128596 200122
rect 128544 200058 128596 200064
rect 128912 200116 128964 200122
rect 128912 200058 128964 200064
rect 128556 190505 128584 200058
rect 128542 190496 128598 190505
rect 128542 190431 128598 190440
rect 128726 190496 128782 190505
rect 128726 190431 128782 190440
rect 128740 186300 128768 190431
rect 128740 186272 128860 186300
rect 128832 182186 128860 186272
rect 128832 182158 128952 182186
rect 128924 180810 128952 182158
rect 128912 180804 128964 180810
rect 128912 180746 128964 180752
rect 129004 171148 129056 171154
rect 129004 171090 129056 171096
rect 129016 164286 129044 171090
rect 128912 164280 128964 164286
rect 128912 164222 128964 164228
rect 129004 164280 129056 164286
rect 129004 164222 129056 164228
rect 128924 157486 128952 164222
rect 128912 157480 128964 157486
rect 128912 157422 128964 157428
rect 128820 157276 128872 157282
rect 128820 157218 128872 157224
rect 128832 142118 128860 157218
rect 128820 142112 128872 142118
rect 128820 142054 128872 142060
rect 128820 133884 128872 133890
rect 128820 133826 128872 133832
rect 128266 118280 128322 118289
rect 128266 118215 128322 118224
rect 126058 117600 126114 117609
rect 125692 117564 125744 117570
rect 126058 117535 126114 117544
rect 125692 117506 125744 117512
rect 123484 117496 123536 117502
rect 123484 117438 123536 117444
rect 124128 117496 124180 117502
rect 124128 117438 124180 117444
rect 122840 117292 122892 117298
rect 122840 117234 122892 117240
rect 123024 5636 123076 5642
rect 123024 5578 123076 5584
rect 122104 4412 122156 4418
rect 122104 4354 122156 4360
rect 123036 480 123064 5578
rect 123496 4282 123524 117438
rect 126072 109018 126100 117535
rect 128280 117337 128308 118215
rect 128832 117638 128860 133826
rect 129108 118182 129136 380559
rect 129186 373280 129242 373289
rect 129186 373215 129242 373224
rect 129200 118250 129228 373215
rect 129370 365936 129426 365945
rect 129370 365871 129426 365880
rect 129384 365702 129412 365871
rect 129372 365696 129424 365702
rect 129372 365638 129424 365644
rect 129278 358320 129334 358329
rect 129278 358255 129334 358264
rect 129292 118386 129320 358255
rect 129280 118380 129332 118386
rect 129280 118322 129332 118328
rect 129188 118244 129240 118250
rect 129188 118186 129240 118192
rect 129096 118176 129148 118182
rect 129096 118118 129148 118124
rect 128820 117632 128872 117638
rect 128820 117574 128872 117580
rect 127622 117328 127678 117337
rect 127622 117263 127678 117272
rect 128266 117328 128322 117337
rect 128266 117263 128322 117272
rect 126072 108990 126192 109018
rect 126164 101402 126192 108990
rect 126164 101374 126284 101402
rect 126256 89758 126284 101374
rect 126060 89752 126112 89758
rect 126244 89752 126296 89758
rect 126112 89700 126244 89706
rect 126060 89694 126296 89700
rect 126072 89678 126284 89694
rect 126256 77314 126284 89678
rect 126244 77308 126296 77314
rect 126244 77250 126296 77256
rect 126336 77308 126388 77314
rect 126336 77250 126388 77256
rect 126348 72434 126376 77250
rect 126256 72406 126376 72434
rect 126256 56710 126284 72406
rect 126244 56704 126296 56710
rect 126244 56646 126296 56652
rect 125968 56636 126020 56642
rect 125968 56578 126020 56584
rect 125980 51134 126008 56578
rect 125968 51128 126020 51134
rect 125968 51070 126020 51076
rect 125968 46980 126020 46986
rect 125968 46922 126020 46928
rect 125980 46850 126008 46922
rect 125968 46844 126020 46850
rect 125968 46786 126020 46792
rect 126152 46844 126204 46850
rect 126152 46786 126204 46792
rect 126164 41392 126192 46786
rect 126072 41364 126192 41392
rect 126072 27606 126100 41364
rect 126060 27600 126112 27606
rect 126060 27542 126112 27548
rect 125968 9716 126020 9722
rect 125968 9658 126020 9664
rect 125416 7336 125468 7342
rect 125416 7278 125468 7284
rect 124220 4412 124272 4418
rect 124220 4354 124272 4360
rect 123484 4276 123536 4282
rect 123484 4218 123536 4224
rect 124232 480 124260 4354
rect 125428 480 125456 7278
rect 125980 4418 126008 9658
rect 126612 7472 126664 7478
rect 126612 7414 126664 7420
rect 125968 4412 126020 4418
rect 125968 4354 126020 4360
rect 126624 480 126652 7414
rect 127636 7410 127664 117263
rect 128832 109018 128860 117574
rect 128832 108990 128952 109018
rect 128924 106282 128952 108990
rect 128912 106276 128964 106282
rect 128912 106218 128964 106224
rect 128912 99340 128964 99346
rect 128912 99282 128964 99288
rect 128924 96642 128952 99282
rect 128924 96626 129044 96642
rect 128912 96620 129056 96626
rect 128964 96614 129004 96620
rect 128912 96562 128964 96568
rect 129004 96562 129056 96568
rect 128924 86970 128952 96562
rect 129016 96531 129044 96562
rect 128728 86964 128780 86970
rect 128728 86906 128780 86912
rect 128912 86964 128964 86970
rect 128912 86906 128964 86912
rect 128740 85542 128768 86906
rect 128728 85536 128780 85542
rect 128728 85478 128780 85484
rect 128636 75948 128688 75954
rect 128636 75890 128688 75896
rect 128648 67697 128676 75890
rect 128634 67688 128690 67697
rect 128634 67623 128690 67632
rect 128818 67688 128874 67697
rect 128818 67623 128874 67632
rect 128832 66230 128860 67623
rect 128820 66224 128872 66230
rect 128820 66166 128872 66172
rect 128912 56636 128964 56642
rect 128912 56578 128964 56584
rect 128924 51066 128952 56578
rect 128912 51060 128964 51066
rect 128912 51002 128964 51008
rect 129004 50992 129056 50998
rect 129004 50934 129056 50940
rect 129016 31822 129044 50934
rect 129004 31816 129056 31822
rect 129004 31758 129056 31764
rect 128912 31748 128964 31754
rect 128912 31690 128964 31696
rect 128924 28966 128952 31690
rect 128912 28960 128964 28966
rect 128912 28902 128964 28908
rect 129004 28892 129056 28898
rect 129004 28834 129056 28840
rect 129016 12594 129044 28834
rect 128924 12566 129044 12594
rect 128924 12458 128952 12566
rect 128832 12430 128952 12458
rect 127624 7404 127676 7410
rect 127624 7346 127676 7352
rect 127808 7268 127860 7274
rect 127808 7210 127860 7216
rect 127820 480 127848 7210
rect 128832 4350 128860 12430
rect 129004 7336 129056 7342
rect 129004 7278 129056 7284
rect 128820 4344 128872 4350
rect 128820 4286 128872 4292
rect 129016 480 129044 7278
rect 129108 7206 129136 118118
rect 129096 7200 129148 7206
rect 129096 7142 129148 7148
rect 129200 7138 129228 118186
rect 129292 8362 129320 118322
rect 129384 117706 129412 365638
rect 129476 117745 129504 397394
rect 129568 118862 129596 563042
rect 129556 118856 129608 118862
rect 129556 118798 129608 118804
rect 129660 118726 129688 582383
rect 130384 578740 130436 578746
rect 130384 578682 130436 578688
rect 130396 518906 130424 578682
rect 129832 518900 129884 518906
rect 129832 518842 129884 518848
rect 130384 518900 130436 518906
rect 130384 518842 130436 518848
rect 129740 398812 129792 398818
rect 129740 398754 129792 398760
rect 129752 398342 129780 398754
rect 129740 398336 129792 398342
rect 129740 398278 129792 398284
rect 129648 118720 129700 118726
rect 129648 118662 129700 118668
rect 129752 118658 129780 398278
rect 129844 351218 129872 518842
rect 131026 500304 131082 500313
rect 131026 500239 131082 500248
rect 130934 500168 130990 500177
rect 130934 500103 130990 500112
rect 130384 407176 130436 407182
rect 130384 407118 130436 407124
rect 130396 398342 130424 407118
rect 130384 398336 130436 398342
rect 130384 398278 130436 398284
rect 129832 351212 129884 351218
rect 129832 351154 129884 351160
rect 130384 351212 130436 351218
rect 130384 351154 130436 351160
rect 130292 342100 130344 342106
rect 130292 342042 130344 342048
rect 130304 342009 130332 342042
rect 130290 342000 130346 342009
rect 130290 341935 130346 341944
rect 130396 340678 130424 351154
rect 130660 342916 130712 342922
rect 130660 342858 130712 342864
rect 130384 340672 130436 340678
rect 130384 340614 130436 340620
rect 130396 339726 130424 340614
rect 130384 339720 130436 339726
rect 130384 339662 130436 339668
rect 130568 201272 130620 201278
rect 130568 201214 130620 201220
rect 130474 196208 130530 196217
rect 130474 196143 130530 196152
rect 130488 196110 130516 196143
rect 130476 196104 130528 196110
rect 130476 196046 130528 196052
rect 130474 194712 130530 194721
rect 130474 194647 130530 194656
rect 130488 194614 130516 194647
rect 130476 194608 130528 194614
rect 130476 194550 130528 194556
rect 130476 194472 130528 194478
rect 130474 194440 130476 194449
rect 130528 194440 130530 194449
rect 130474 194375 130530 194384
rect 130384 193180 130436 193186
rect 130384 193122 130436 193128
rect 130396 192545 130424 193122
rect 130476 193112 130528 193118
rect 130474 193080 130476 193089
rect 130528 193080 130530 193089
rect 130474 193015 130530 193024
rect 130382 192536 130438 192545
rect 130382 192471 130438 192480
rect 130476 191820 130528 191826
rect 130476 191762 130528 191768
rect 130488 191457 130516 191762
rect 130474 191448 130530 191457
rect 130474 191383 130530 191392
rect 130476 190460 130528 190466
rect 130476 190402 130528 190408
rect 130488 190369 130516 190402
rect 130474 190360 130530 190369
rect 130474 190295 130530 190304
rect 130384 189032 130436 189038
rect 130384 188974 130436 188980
rect 130396 188329 130424 188974
rect 130476 188964 130528 188970
rect 130476 188906 130528 188912
rect 130488 188873 130516 188906
rect 130474 188864 130530 188873
rect 130474 188799 130530 188808
rect 130382 188320 130438 188329
rect 130382 188255 130438 188264
rect 130476 187672 130528 187678
rect 130476 187614 130528 187620
rect 130488 187241 130516 187614
rect 130474 187232 130530 187241
rect 130474 187167 130530 187176
rect 129740 118652 129792 118658
rect 129740 118594 129792 118600
rect 129462 117736 129518 117745
rect 129372 117700 129424 117706
rect 129462 117671 129518 117680
rect 129372 117642 129424 117648
rect 130384 117564 130436 117570
rect 130384 117506 130436 117512
rect 129280 8356 129332 8362
rect 129280 8298 129332 8304
rect 129188 7132 129240 7138
rect 129188 7074 129240 7080
rect 130200 7132 130252 7138
rect 130200 7074 130252 7080
rect 130212 480 130240 7074
rect 130396 4486 130424 117506
rect 130580 117502 130608 201214
rect 130672 135590 130700 342858
rect 130752 340196 130804 340202
rect 130752 340138 130804 340144
rect 130660 135584 130712 135590
rect 130660 135526 130712 135532
rect 130764 118998 130792 340138
rect 130844 339720 130896 339726
rect 130844 339662 130896 339668
rect 130752 118992 130804 118998
rect 130752 118934 130804 118940
rect 130856 117570 130884 339662
rect 130948 118930 130976 500103
rect 130936 118924 130988 118930
rect 130936 118866 130988 118872
rect 131040 118794 131068 500239
rect 131132 156330 131160 700674
rect 131212 700596 131264 700602
rect 131212 700538 131264 700544
rect 131224 186318 131252 700538
rect 132316 700528 132368 700534
rect 132316 700470 132368 700476
rect 132132 498228 132184 498234
rect 132132 498170 132184 498176
rect 131948 341692 132000 341698
rect 131948 341634 132000 341640
rect 131672 341556 131724 341562
rect 131672 341498 131724 341504
rect 131580 263628 131632 263634
rect 131580 263570 131632 263576
rect 131304 227792 131356 227798
rect 131304 227734 131356 227740
rect 131212 186312 131264 186318
rect 131212 186254 131264 186260
rect 131212 186176 131264 186182
rect 131212 186118 131264 186124
rect 131224 185609 131252 186118
rect 131210 185600 131266 185609
rect 131210 185535 131266 185544
rect 131212 184884 131264 184890
rect 131212 184826 131264 184832
rect 131224 184521 131252 184826
rect 131210 184512 131266 184521
rect 131210 184447 131266 184456
rect 131210 183560 131266 183569
rect 131210 183495 131212 183504
rect 131264 183495 131266 183504
rect 131212 183466 131264 183472
rect 131212 183388 131264 183394
rect 131212 183330 131264 183336
rect 131224 178265 131252 183330
rect 131210 178256 131266 178265
rect 131210 178191 131266 178200
rect 131316 164529 131344 227734
rect 131488 216708 131540 216714
rect 131488 216650 131540 216656
rect 131396 200796 131448 200802
rect 131396 200738 131448 200744
rect 131408 198354 131436 200738
rect 131396 198348 131448 198354
rect 131396 198290 131448 198296
rect 131394 198248 131450 198257
rect 131394 198183 131450 198192
rect 131408 197402 131436 198183
rect 131396 197396 131448 197402
rect 131396 197338 131448 197344
rect 131394 197160 131450 197169
rect 131394 197095 131450 197104
rect 131408 196314 131436 197095
rect 131396 196308 131448 196314
rect 131396 196250 131448 196256
rect 131396 196036 131448 196042
rect 131396 195978 131448 195984
rect 131302 164520 131358 164529
rect 131302 164455 131358 164464
rect 131210 161392 131266 161401
rect 131210 161327 131266 161336
rect 131224 157350 131252 161327
rect 131212 157344 131264 157350
rect 131212 157286 131264 157292
rect 131302 157176 131358 157185
rect 131302 157111 131358 157120
rect 131120 156324 131172 156330
rect 131120 156266 131172 156272
rect 131118 156224 131174 156233
rect 131118 156159 131174 156168
rect 131132 156058 131160 156159
rect 131316 156126 131344 157111
rect 131304 156120 131356 156126
rect 131304 156062 131356 156068
rect 131120 156052 131172 156058
rect 131120 155994 131172 156000
rect 131304 155984 131356 155990
rect 131304 155926 131356 155932
rect 131120 155916 131172 155922
rect 131120 155858 131172 155864
rect 131132 155145 131160 155858
rect 131118 155136 131174 155145
rect 131118 155071 131174 155080
rect 131120 153196 131172 153202
rect 131120 153138 131172 153144
rect 131132 152969 131160 153138
rect 131316 153134 131344 155926
rect 131304 153128 131356 153134
rect 131304 153070 131356 153076
rect 131118 152960 131174 152969
rect 131118 152895 131174 152904
rect 131212 152924 131264 152930
rect 131212 152866 131264 152872
rect 131224 152017 131252 152866
rect 131210 152008 131266 152017
rect 131210 151943 131266 151952
rect 131304 151904 131356 151910
rect 131304 151846 131356 151852
rect 131120 151768 131172 151774
rect 131120 151710 131172 151716
rect 131132 150929 131160 151710
rect 131118 150920 131174 150929
rect 131118 150855 131174 150864
rect 131120 150408 131172 150414
rect 131120 150350 131172 150356
rect 131132 149841 131160 150350
rect 131118 149832 131174 149841
rect 131118 149767 131174 149776
rect 131120 148980 131172 148986
rect 131120 148922 131172 148928
rect 131132 148753 131160 148922
rect 131118 148744 131174 148753
rect 131118 148679 131174 148688
rect 131120 148640 131172 148646
rect 131120 148582 131172 148588
rect 131132 147801 131160 148582
rect 131118 147792 131174 147801
rect 131118 147727 131174 147736
rect 131212 147688 131264 147694
rect 131212 147630 131264 147636
rect 131120 147620 131172 147626
rect 131120 147562 131172 147568
rect 131132 146713 131160 147562
rect 131118 146704 131174 146713
rect 131118 146639 131174 146648
rect 131120 146260 131172 146266
rect 131120 146202 131172 146208
rect 131132 145625 131160 146202
rect 131118 145616 131174 145625
rect 131118 145551 131174 145560
rect 131120 144424 131172 144430
rect 131120 144366 131172 144372
rect 131132 143585 131160 144366
rect 131118 143576 131174 143585
rect 131118 143511 131174 143520
rect 131224 137714 131252 147630
rect 131316 139369 131344 151846
rect 131302 139360 131358 139369
rect 131302 139295 131358 139304
rect 131132 137686 131252 137714
rect 131132 133890 131160 137686
rect 131120 133884 131172 133890
rect 131120 133826 131172 133832
rect 131304 133884 131356 133890
rect 131304 133826 131356 133832
rect 131316 124273 131344 133826
rect 131408 132025 131436 195978
rect 131394 132016 131450 132025
rect 131394 131951 131450 131960
rect 131500 124545 131528 216650
rect 131592 125633 131620 263570
rect 131684 167793 131712 341498
rect 131856 310548 131908 310554
rect 131856 310490 131908 310496
rect 131762 199336 131818 199345
rect 131762 199271 131818 199280
rect 131776 196110 131804 199271
rect 131764 196104 131816 196110
rect 131764 196046 131816 196052
rect 131764 195968 131816 195974
rect 131764 195910 131816 195916
rect 131670 167784 131726 167793
rect 131670 167719 131726 167728
rect 131670 158264 131726 158273
rect 131670 158199 131726 158208
rect 131578 125624 131634 125633
rect 131578 125559 131634 125568
rect 131486 124536 131542 124545
rect 131486 124471 131542 124480
rect 131118 124264 131174 124273
rect 131118 124199 131174 124208
rect 131302 124264 131358 124273
rect 131302 124199 131358 124208
rect 131132 124166 131160 124199
rect 131120 124160 131172 124166
rect 131120 124102 131172 124108
rect 131396 124160 131448 124166
rect 131396 124102 131448 124108
rect 131028 118788 131080 118794
rect 131028 118730 131080 118736
rect 130844 117564 130896 117570
rect 130844 117506 130896 117512
rect 130568 117496 130620 117502
rect 130568 117438 130620 117444
rect 131408 96665 131436 124102
rect 131210 96656 131266 96665
rect 131210 96591 131266 96600
rect 131394 96656 131450 96665
rect 131394 96591 131450 96600
rect 131224 88330 131252 96591
rect 131212 88324 131264 88330
rect 131212 88266 131264 88272
rect 131684 64870 131712 158199
rect 131672 64864 131724 64870
rect 131672 64806 131724 64812
rect 131776 8294 131804 195910
rect 131868 126721 131896 310490
rect 131960 128761 131988 341634
rect 132040 341624 132092 341630
rect 132040 341566 132092 341572
rect 131946 128752 132002 128761
rect 131946 128687 132002 128696
rect 132052 127809 132080 341566
rect 132144 130937 132172 498170
rect 132224 200864 132276 200870
rect 132224 200806 132276 200812
rect 132236 170921 132264 200806
rect 132222 170912 132278 170921
rect 132222 170847 132278 170856
rect 132222 159352 132278 159361
rect 132222 159287 132278 159296
rect 132130 130928 132186 130937
rect 132130 130863 132186 130872
rect 132038 127800 132094 127809
rect 132038 127735 132094 127744
rect 131854 126712 131910 126721
rect 131854 126647 131910 126656
rect 132130 121408 132186 121417
rect 132130 121343 132186 121352
rect 132144 77246 132172 121343
rect 132132 77240 132184 77246
rect 132132 77182 132184 77188
rect 132236 22098 132264 159287
rect 132328 138281 132356 700470
rect 132512 342038 132540 700810
rect 133696 700800 133748 700806
rect 133696 700742 133748 700748
rect 132592 700392 132644 700398
rect 132592 700334 132644 700340
rect 132500 342032 132552 342038
rect 132500 341974 132552 341980
rect 132500 341896 132552 341902
rect 132500 341838 132552 341844
rect 132408 200932 132460 200938
rect 132408 200874 132460 200880
rect 132420 172009 132448 200874
rect 132512 179353 132540 341838
rect 132498 179344 132554 179353
rect 132498 179279 132554 179288
rect 132604 177177 132632 700334
rect 133420 700256 133472 700262
rect 133420 700198 133472 700204
rect 133328 699712 133380 699718
rect 133328 699654 133380 699660
rect 133144 462392 133196 462398
rect 133144 462334 133196 462340
rect 132960 415472 133012 415478
rect 132960 415414 133012 415420
rect 132868 405748 132920 405754
rect 132868 405690 132920 405696
rect 132880 398834 132908 405690
rect 132696 398818 132908 398834
rect 132684 398812 132920 398818
rect 132736 398806 132868 398812
rect 132684 398754 132736 398760
rect 132868 398754 132920 398760
rect 132696 398723 132724 398754
rect 132880 389298 132908 398754
rect 132868 389292 132920 389298
rect 132868 389234 132920 389240
rect 132868 389156 132920 389162
rect 132868 389098 132920 389104
rect 132880 376854 132908 389098
rect 132776 376848 132828 376854
rect 132696 376796 132776 376802
rect 132696 376790 132828 376796
rect 132868 376848 132920 376854
rect 132868 376790 132920 376796
rect 132696 376774 132816 376790
rect 132696 375358 132724 376774
rect 132684 375352 132736 375358
rect 132684 375294 132736 375300
rect 132776 366988 132828 366994
rect 132776 366930 132828 366936
rect 132788 360262 132816 366930
rect 132972 366926 133000 415414
rect 133052 398132 133104 398138
rect 133052 398074 133104 398080
rect 133064 397594 133092 398074
rect 133052 397588 133104 397594
rect 133052 397530 133104 397536
rect 133064 367062 133092 397530
rect 133156 367062 133184 462334
rect 133236 451308 133288 451314
rect 133236 451250 133288 451256
rect 133052 367056 133104 367062
rect 133052 366998 133104 367004
rect 133144 367056 133196 367062
rect 133144 366998 133196 367004
rect 132960 366920 133012 366926
rect 132960 366862 133012 366868
rect 133052 366852 133104 366858
rect 133052 366794 133104 366800
rect 132960 366784 133012 366790
rect 132960 366726 133012 366732
rect 132776 360256 132828 360262
rect 132776 360198 132828 360204
rect 132776 360120 132828 360126
rect 132776 360062 132828 360068
rect 132788 357354 132816 360062
rect 132788 357326 132908 357354
rect 132880 347818 132908 357326
rect 132684 347812 132736 347818
rect 132684 347754 132736 347760
rect 132868 347812 132920 347818
rect 132868 347754 132920 347760
rect 132696 342106 132724 347754
rect 132684 342100 132736 342106
rect 132684 342042 132736 342048
rect 132868 340604 132920 340610
rect 132868 340546 132920 340552
rect 132880 333282 132908 340546
rect 132972 338026 133000 366726
rect 133064 338026 133092 366794
rect 133144 358692 133196 358698
rect 133144 358634 133196 358640
rect 133156 338026 133184 358634
rect 132960 338020 133012 338026
rect 132960 337962 133012 337968
rect 133052 338020 133104 338026
rect 133052 337962 133104 337968
rect 133144 338020 133196 338026
rect 133144 337962 133196 337968
rect 132960 337884 133012 337890
rect 132960 337826 133012 337832
rect 133052 337884 133104 337890
rect 133052 337826 133104 337832
rect 132696 333254 132908 333282
rect 132696 329338 132724 333254
rect 132696 329310 132816 329338
rect 132788 321722 132816 329310
rect 132696 321694 132816 321722
rect 132696 308310 132724 321694
rect 132776 321632 132828 321638
rect 132776 321574 132828 321580
rect 132684 308304 132736 308310
rect 132684 308246 132736 308252
rect 132684 296132 132736 296138
rect 132684 296074 132736 296080
rect 132696 288998 132724 296074
rect 132684 288992 132736 288998
rect 132684 288934 132736 288940
rect 132684 274712 132736 274718
rect 132684 274654 132736 274660
rect 132590 177168 132646 177177
rect 132590 177103 132646 177112
rect 132406 172000 132462 172009
rect 132406 171935 132462 171944
rect 132696 165617 132724 274654
rect 132788 166705 132816 321574
rect 132868 308304 132920 308310
rect 132868 308246 132920 308252
rect 132880 296138 132908 308246
rect 132868 296132 132920 296138
rect 132868 296074 132920 296080
rect 132868 288992 132920 288998
rect 132868 288934 132920 288940
rect 132880 278118 132908 288934
rect 132868 278112 132920 278118
rect 132868 278054 132920 278060
rect 132868 268456 132920 268462
rect 132868 268398 132920 268404
rect 132880 258806 132908 268398
rect 132868 258800 132920 258806
rect 132868 258742 132920 258748
rect 132868 249144 132920 249150
rect 132868 249086 132920 249092
rect 132880 239494 132908 249086
rect 132868 239488 132920 239494
rect 132868 239430 132920 239436
rect 132868 229764 132920 229770
rect 132868 229706 132920 229712
rect 132880 220114 132908 229706
rect 132868 220108 132920 220114
rect 132868 220050 132920 220056
rect 132868 210452 132920 210458
rect 132868 210394 132920 210400
rect 132880 196110 132908 210394
rect 132868 196104 132920 196110
rect 132868 196046 132920 196052
rect 132868 195968 132920 195974
rect 132868 195910 132920 195916
rect 132880 181490 132908 195910
rect 132868 181484 132920 181490
rect 132868 181426 132920 181432
rect 132972 168745 133000 337826
rect 132958 168736 133014 168745
rect 132958 168671 133014 168680
rect 132960 168632 133012 168638
rect 132960 168574 133012 168580
rect 132774 166696 132830 166705
rect 132774 166631 132830 166640
rect 132682 165608 132738 165617
rect 132682 165543 132738 165552
rect 132406 162480 132462 162489
rect 132406 162415 132462 162424
rect 132314 138272 132370 138281
rect 132314 138207 132370 138216
rect 132316 135584 132368 135590
rect 132316 135526 132368 135532
rect 132328 132462 132356 135526
rect 132316 132456 132368 132462
rect 132316 132398 132368 132404
rect 132420 120766 132448 162415
rect 132972 153218 133000 168574
rect 132880 153190 133000 153218
rect 132880 143614 132908 153190
rect 132868 143608 132920 143614
rect 132868 143550 132920 143556
rect 132776 142180 132828 142186
rect 132776 142122 132828 142128
rect 132788 132410 132816 142122
rect 132696 132382 132816 132410
rect 132696 125474 132724 132382
rect 132696 125446 132908 125474
rect 132408 120760 132460 120766
rect 132408 120702 132460 120708
rect 132406 120456 132462 120465
rect 132406 120391 132462 120400
rect 132420 30326 132448 120391
rect 132880 118153 132908 125446
rect 132866 118144 132922 118153
rect 132866 118079 132922 118088
rect 133064 118017 133092 337826
rect 133144 333328 133196 333334
rect 133144 333270 133196 333276
rect 133156 169833 133184 333270
rect 133142 169824 133198 169833
rect 133142 169759 133198 169768
rect 133144 132388 133196 132394
rect 133144 132330 133196 132336
rect 133156 120358 133184 132330
rect 133248 129849 133276 451250
rect 133340 182481 133368 699654
rect 133326 182472 133382 182481
rect 133326 182407 133382 182416
rect 133328 181484 133380 181490
rect 133328 181426 133380 181432
rect 133340 168638 133368 181426
rect 133432 181393 133460 700198
rect 133512 278112 133564 278118
rect 133512 278054 133564 278060
rect 133524 268462 133552 278054
rect 133512 268456 133564 268462
rect 133512 268398 133564 268404
rect 133512 258800 133564 258806
rect 133512 258742 133564 258748
rect 133524 249150 133552 258742
rect 133512 249144 133564 249150
rect 133512 249086 133564 249092
rect 133512 239488 133564 239494
rect 133512 239430 133564 239436
rect 133524 229770 133552 239430
rect 133512 229764 133564 229770
rect 133512 229706 133564 229712
rect 133512 220108 133564 220114
rect 133512 220050 133564 220056
rect 133524 210458 133552 220050
rect 133512 210452 133564 210458
rect 133512 210394 133564 210400
rect 133512 201204 133564 201210
rect 133512 201146 133564 201152
rect 133418 181384 133474 181393
rect 133418 181319 133474 181328
rect 133328 168632 133380 168638
rect 133328 168574 133380 168580
rect 133524 142497 133552 201146
rect 133604 199844 133656 199850
rect 133604 199786 133656 199792
rect 133616 163577 133644 199786
rect 133602 163568 133658 163577
rect 133602 163503 133658 163512
rect 133602 160440 133658 160449
rect 133602 160375 133658 160384
rect 133510 142488 133566 142497
rect 133510 142423 133566 142432
rect 133234 129840 133290 129849
rect 133234 129775 133290 129784
rect 133144 120352 133196 120358
rect 133144 120294 133196 120300
rect 133326 118144 133382 118153
rect 133326 118079 133382 118088
rect 133050 118008 133106 118017
rect 133050 117943 133106 117952
rect 133340 60738 133368 118079
rect 133248 60710 133368 60738
rect 133248 60602 133276 60710
rect 133248 60574 133368 60602
rect 133340 46918 133368 60574
rect 133328 46912 133380 46918
rect 133328 46854 133380 46860
rect 133616 41410 133644 160375
rect 133708 141409 133736 700742
rect 133694 141400 133750 141409
rect 133694 141335 133750 141344
rect 133800 140457 133828 700878
rect 133984 180713 134012 700946
rect 137848 699718 137876 703520
rect 154132 703474 154160 703520
rect 154132 703446 154252 703474
rect 137836 699712 137888 699718
rect 137836 699654 137888 699660
rect 154224 698290 154252 703446
rect 170324 700670 170352 703520
rect 170312 700664 170364 700670
rect 170312 700606 170364 700612
rect 202800 700262 202828 703520
rect 218992 700806 219020 703520
rect 235184 700806 235212 703520
rect 267660 701010 267688 703520
rect 267648 701004 267700 701010
rect 267648 700946 267700 700952
rect 283852 700942 283880 703520
rect 300136 700942 300164 703520
rect 283840 700936 283892 700942
rect 283840 700878 283892 700884
rect 300124 700936 300176 700942
rect 300124 700878 300176 700884
rect 332520 700874 332548 703520
rect 332508 700868 332560 700874
rect 332508 700810 332560 700816
rect 218980 700800 219032 700806
rect 218980 700742 219032 700748
rect 235172 700800 235224 700806
rect 235172 700742 235224 700748
rect 348804 700738 348832 703520
rect 364996 700738 365024 703520
rect 348792 700732 348844 700738
rect 348792 700674 348844 700680
rect 364984 700732 365036 700738
rect 364984 700674 365036 700680
rect 397472 700602 397500 703520
rect 397460 700596 397512 700602
rect 397460 700538 397512 700544
rect 413664 700534 413692 703520
rect 413652 700528 413704 700534
rect 413652 700470 413704 700476
rect 202788 700256 202840 700262
rect 202788 700198 202840 700204
rect 429856 699718 429884 703520
rect 434076 700936 434128 700942
rect 434076 700878 434128 700884
rect 433984 700732 434036 700738
rect 433984 700674 434036 700680
rect 429844 699712 429896 699718
rect 429844 699654 429896 699660
rect 433892 699712 433944 699718
rect 433892 699654 433944 699660
rect 153568 698284 153620 698290
rect 153568 698226 153620 698232
rect 154212 698284 154264 698290
rect 154212 698226 154264 698232
rect 147588 697128 147640 697134
rect 147586 697096 147588 697105
rect 147640 697096 147642 697105
rect 147586 697031 147642 697040
rect 153580 688786 153608 698226
rect 154486 697232 154542 697241
rect 154486 697167 154542 697176
rect 173806 697232 173862 697241
rect 173806 697167 173862 697176
rect 193126 697232 193182 697241
rect 193126 697167 193182 697176
rect 212446 697232 212502 697241
rect 212446 697167 212502 697176
rect 231766 697232 231822 697241
rect 231766 697167 231822 697176
rect 251086 697232 251142 697241
rect 251086 697167 251142 697176
rect 270406 697232 270462 697241
rect 270406 697167 270462 697176
rect 289726 697232 289782 697241
rect 289726 697167 289782 697176
rect 309046 697232 309102 697241
rect 309046 697167 309102 697176
rect 328366 697232 328422 697241
rect 328366 697167 328422 697176
rect 154500 697134 154528 697167
rect 173820 697134 173848 697167
rect 193140 697134 193168 697167
rect 212460 697134 212488 697167
rect 231780 697134 231808 697167
rect 251100 697134 251128 697167
rect 270420 697134 270448 697167
rect 289740 697134 289768 697167
rect 309060 697134 309088 697167
rect 328380 697134 328408 697167
rect 154488 697128 154540 697134
rect 166908 697128 166960 697134
rect 154488 697070 154540 697076
rect 166906 697096 166908 697105
rect 173808 697128 173860 697134
rect 166960 697096 166962 697105
rect 186228 697128 186280 697134
rect 173808 697070 173860 697076
rect 186226 697096 186228 697105
rect 193128 697128 193180 697134
rect 186280 697096 186282 697105
rect 166906 697031 166962 697040
rect 205548 697128 205600 697134
rect 193128 697070 193180 697076
rect 205546 697096 205548 697105
rect 212448 697128 212500 697134
rect 205600 697096 205602 697105
rect 186226 697031 186282 697040
rect 224868 697128 224920 697134
rect 212448 697070 212500 697076
rect 224866 697096 224868 697105
rect 231768 697128 231820 697134
rect 224920 697096 224922 697105
rect 205546 697031 205602 697040
rect 244188 697128 244240 697134
rect 231768 697070 231820 697076
rect 244186 697096 244188 697105
rect 251088 697128 251140 697134
rect 244240 697096 244242 697105
rect 224866 697031 224922 697040
rect 263508 697128 263560 697134
rect 251088 697070 251140 697076
rect 263506 697096 263508 697105
rect 270408 697128 270460 697134
rect 263560 697096 263562 697105
rect 244186 697031 244242 697040
rect 282828 697128 282880 697134
rect 270408 697070 270460 697076
rect 282826 697096 282828 697105
rect 289728 697128 289780 697134
rect 282880 697096 282882 697105
rect 263506 697031 263562 697040
rect 302148 697128 302200 697134
rect 289728 697070 289780 697076
rect 302146 697096 302148 697105
rect 309048 697128 309100 697134
rect 302200 697096 302202 697105
rect 282826 697031 282882 697040
rect 321468 697128 321520 697134
rect 309048 697070 309100 697076
rect 321466 697096 321468 697105
rect 328368 697128 328420 697134
rect 321520 697096 321522 697105
rect 302146 697031 302202 697040
rect 328368 697070 328420 697076
rect 321466 697031 321522 697040
rect 153580 688758 153700 688786
rect 147770 686352 147826 686361
rect 147600 686310 147770 686338
rect 135258 686216 135314 686225
rect 135258 686151 135260 686160
rect 135312 686151 135314 686160
rect 142896 686180 142948 686186
rect 135260 686122 135312 686128
rect 142896 686122 142948 686128
rect 142908 685953 142936 686122
rect 147600 686089 147628 686310
rect 147770 686287 147826 686296
rect 147586 686080 147642 686089
rect 147586 686015 147642 686024
rect 153672 685982 153700 688758
rect 169022 686488 169078 686497
rect 169022 686423 169078 686432
rect 154578 686352 154634 686361
rect 154578 686287 154580 686296
rect 154632 686287 154634 686296
rect 159456 686316 159508 686322
rect 154580 686258 154632 686264
rect 159456 686258 159508 686264
rect 159468 686225 159496 686258
rect 169036 686225 169064 686423
rect 159454 686216 159510 686225
rect 159454 686151 159510 686160
rect 169022 686216 169078 686225
rect 169022 686151 169078 686160
rect 153292 685976 153344 685982
rect 142894 685944 142950 685953
rect 153292 685918 153344 685924
rect 153660 685976 153712 685982
rect 153660 685918 153712 685924
rect 142894 685879 142950 685888
rect 153304 684486 153332 685918
rect 153292 684480 153344 684486
rect 153292 684422 153344 684428
rect 153660 666596 153712 666602
rect 153660 666538 153712 666544
rect 153672 659682 153700 666538
rect 153488 659654 153700 659682
rect 153488 656878 153516 659654
rect 153476 656872 153528 656878
rect 153476 656814 153528 656820
rect 169022 650584 169078 650593
rect 169022 650519 169078 650528
rect 147770 650448 147826 650457
rect 147600 650406 147770 650434
rect 135258 650312 135314 650321
rect 135258 650247 135260 650256
rect 135312 650247 135314 650256
rect 142896 650276 142948 650282
rect 135260 650218 135312 650224
rect 142896 650218 142948 650224
rect 142908 650049 142936 650218
rect 147600 650185 147628 650406
rect 147770 650383 147826 650392
rect 154578 650448 154634 650457
rect 154578 650383 154580 650392
rect 154632 650383 154634 650392
rect 159456 650412 159508 650418
rect 154580 650354 154632 650360
rect 159456 650354 159508 650360
rect 159468 650321 159496 650354
rect 169036 650321 169064 650519
rect 159454 650312 159510 650321
rect 159454 650247 159510 650256
rect 169022 650312 169078 650321
rect 169022 650247 169078 650256
rect 147586 650176 147642 650185
rect 147586 650111 147642 650120
rect 142894 650040 142950 650049
rect 142894 649975 142950 649984
rect 153568 647284 153620 647290
rect 153568 647226 153620 647232
rect 153580 637702 153608 647226
rect 157062 639296 157118 639305
rect 157246 639296 157302 639305
rect 157118 639254 157246 639282
rect 157062 639231 157118 639240
rect 157246 639231 157302 639240
rect 171046 639296 171102 639305
rect 171046 639231 171102 639240
rect 171060 638897 171088 639231
rect 171046 638888 171102 638897
rect 171046 638823 171102 638832
rect 153292 637696 153344 637702
rect 153568 637696 153620 637702
rect 153344 637644 153424 637650
rect 153292 637638 153424 637644
rect 153568 637638 153620 637644
rect 153304 637622 153424 637638
rect 153396 630766 153424 637622
rect 153384 630760 153436 630766
rect 153384 630702 153436 630708
rect 153568 630556 153620 630562
rect 153568 630498 153620 630504
rect 153580 626550 153608 630498
rect 153568 626544 153620 626550
rect 153568 626486 153620 626492
rect 153752 626544 153804 626550
rect 153752 626486 153804 626492
rect 153764 611250 153792 626486
rect 153568 611244 153620 611250
rect 153568 611186 153620 611192
rect 153752 611244 153804 611250
rect 153752 611186 153804 611192
rect 153580 599010 153608 611186
rect 157062 603392 157118 603401
rect 157246 603392 157302 603401
rect 157118 603350 157246 603378
rect 157062 603327 157118 603336
rect 157246 603327 157302 603336
rect 171046 603392 171102 603401
rect 171046 603327 171102 603336
rect 171060 602993 171088 603327
rect 171046 602984 171102 602993
rect 171046 602919 171102 602928
rect 153384 599004 153436 599010
rect 153384 598946 153436 598952
rect 153568 599004 153620 599010
rect 153568 598946 153620 598952
rect 153396 598913 153424 598946
rect 153382 598904 153438 598913
rect 153382 598839 153438 598848
rect 153566 598904 153622 598913
rect 153566 598839 153622 598848
rect 153580 592006 153608 598839
rect 157062 592376 157118 592385
rect 157246 592376 157302 592385
rect 157118 592334 157246 592362
rect 157062 592311 157118 592320
rect 157246 592311 157302 592320
rect 171046 592376 171102 592385
rect 171046 592311 171102 592320
rect 153292 592000 153344 592006
rect 153292 591942 153344 591948
rect 153568 592000 153620 592006
rect 171060 591977 171088 592311
rect 153568 591942 153620 591948
rect 171046 591968 171102 591977
rect 153304 582434 153332 591942
rect 171046 591903 171102 591912
rect 175924 583704 175976 583710
rect 175924 583646 175976 583652
rect 302792 583704 302844 583710
rect 302792 583646 302844 583652
rect 153304 582406 153424 582434
rect 153396 579630 153424 582406
rect 153384 579624 153436 579630
rect 153384 579566 153436 579572
rect 153476 569968 153528 569974
rect 153476 569910 153528 569916
rect 153488 563174 153516 569910
rect 153476 563168 153528 563174
rect 153476 563110 153528 563116
rect 153292 563032 153344 563038
rect 153292 562974 153344 562980
rect 153304 560250 153332 562974
rect 153292 560244 153344 560250
rect 153292 560186 153344 560192
rect 162124 553920 162176 553926
rect 162124 553862 162176 553868
rect 140044 553648 140096 553654
rect 140044 553590 140096 553596
rect 134064 337612 134116 337618
rect 134064 337554 134116 337560
rect 133970 180704 134026 180713
rect 133970 180639 134026 180648
rect 133786 140448 133842 140457
rect 133786 140383 133842 140392
rect 133970 123040 134026 123049
rect 133970 122975 134026 122984
rect 133984 120698 134012 122975
rect 134076 122398 134104 337554
rect 140056 202298 140084 553590
rect 151084 553580 151136 553586
rect 151084 553522 151136 553528
rect 146944 536852 146996 536858
rect 146944 536794 146996 536800
rect 144184 518424 144236 518430
rect 144184 518366 144236 518372
rect 144196 497894 144224 518366
rect 144184 497888 144236 497894
rect 144184 497830 144236 497836
rect 144196 397526 144224 497830
rect 144184 397520 144236 397526
rect 144184 397462 144236 397468
rect 140780 384328 140832 384334
rect 140780 384270 140832 384276
rect 140792 340610 140820 384270
rect 144196 357406 144224 397462
rect 144184 357400 144236 357406
rect 144184 357342 144236 357348
rect 145564 357400 145616 357406
rect 145564 357342 145616 357348
rect 140780 340604 140832 340610
rect 140780 340546 140832 340552
rect 140792 340202 140820 340546
rect 145576 340542 145604 357342
rect 145564 340536 145616 340542
rect 145564 340478 145616 340484
rect 140780 340196 140832 340202
rect 140780 340138 140832 340144
rect 140044 202292 140096 202298
rect 140044 202234 140096 202240
rect 142528 202224 142580 202230
rect 142528 202166 142580 202172
rect 134708 202156 134760 202162
rect 134708 202098 134760 202104
rect 134156 201612 134208 201618
rect 134156 201554 134208 201560
rect 134168 200002 134196 201554
rect 134340 201544 134392 201550
rect 134340 201486 134392 201492
rect 134352 200002 134380 201486
rect 134720 200002 134748 202098
rect 142540 200002 142568 202166
rect 145576 201278 145604 340478
rect 146956 202162 146984 536794
rect 151096 202230 151124 553522
rect 157984 553512 158036 553518
rect 157984 553454 158036 553460
rect 153476 550656 153528 550662
rect 153476 550598 153528 550604
rect 153488 543658 153516 550598
rect 153292 543652 153344 543658
rect 153292 543594 153344 543600
rect 153476 543652 153528 543658
rect 153476 543594 153528 543600
rect 153304 534070 153332 543594
rect 153292 534064 153344 534070
rect 153292 534006 153344 534012
rect 153476 534064 153528 534070
rect 153476 534006 153528 534012
rect 153488 531321 153516 534006
rect 153474 531312 153530 531321
rect 153474 531247 153530 531256
rect 153750 531312 153806 531321
rect 153750 531247 153806 531256
rect 153764 521694 153792 531247
rect 153568 521688 153620 521694
rect 153568 521630 153620 521636
rect 153752 521688 153804 521694
rect 153752 521630 153804 521636
rect 153580 514706 153608 521630
rect 153844 518356 153896 518362
rect 153844 518298 153896 518304
rect 153488 514678 153608 514706
rect 153488 511986 153516 514678
rect 153396 511958 153516 511986
rect 153396 505170 153424 511958
rect 153384 505164 153436 505170
rect 153384 505106 153436 505112
rect 153384 502376 153436 502382
rect 153384 502318 153436 502324
rect 153396 495446 153424 502318
rect 153384 495440 153436 495446
rect 153384 495382 153436 495388
rect 153568 495440 153620 495446
rect 153568 495382 153620 495388
rect 153580 492658 153608 495382
rect 153292 492652 153344 492658
rect 153292 492594 153344 492600
rect 153568 492652 153620 492658
rect 153568 492594 153620 492600
rect 153304 483041 153332 492594
rect 153290 483032 153346 483041
rect 153290 482967 153346 482976
rect 153474 483032 153530 483041
rect 153474 482967 153530 482976
rect 153488 476134 153516 482967
rect 153292 476128 153344 476134
rect 153476 476128 153528 476134
rect 153344 476076 153424 476082
rect 153292 476070 153424 476076
rect 153476 476070 153528 476076
rect 153304 476054 153424 476070
rect 153396 466478 153424 476054
rect 153384 466472 153436 466478
rect 153384 466414 153436 466420
rect 153476 466404 153528 466410
rect 153476 466346 153528 466352
rect 153488 463690 153516 466346
rect 153476 463684 153528 463690
rect 153476 463626 153528 463632
rect 153476 456748 153528 456754
rect 153476 456690 153528 456696
rect 153488 454050 153516 456690
rect 153488 454022 153608 454050
rect 153580 447166 153608 454022
rect 153384 447160 153436 447166
rect 153384 447102 153436 447108
rect 153568 447160 153620 447166
rect 153568 447102 153620 447108
rect 153396 444378 153424 447102
rect 153384 444372 153436 444378
rect 153384 444314 153436 444320
rect 153384 437436 153436 437442
rect 153384 437378 153436 437384
rect 153396 434738 153424 437378
rect 153396 434710 153516 434738
rect 153488 425241 153516 434710
rect 153474 425232 153530 425241
rect 153474 425167 153530 425176
rect 153198 425096 153254 425105
rect 153254 425054 153332 425082
rect 153198 425031 153254 425040
rect 153304 418266 153332 425054
rect 153292 418260 153344 418266
rect 153292 418202 153344 418208
rect 153200 418124 153252 418130
rect 153200 418066 153252 418072
rect 153212 408542 153240 418066
rect 153200 408536 153252 408542
rect 153200 408478 153252 408484
rect 153384 408468 153436 408474
rect 153384 408410 153436 408416
rect 153396 398954 153424 408410
rect 153384 398948 153436 398954
rect 153384 398890 153436 398896
rect 153384 396092 153436 396098
rect 153384 396034 153436 396040
rect 153396 395962 153424 396034
rect 153384 395956 153436 395962
rect 153384 395898 153436 395904
rect 153292 389156 153344 389162
rect 153292 389098 153344 389104
rect 153304 379506 153332 389098
rect 153292 379500 153344 379506
rect 153292 379442 153344 379448
rect 153476 379500 153528 379506
rect 153476 379442 153528 379448
rect 153488 371906 153516 379442
rect 153488 371878 153608 371906
rect 153580 367062 153608 371878
rect 153568 367056 153620 367062
rect 153568 366998 153620 367004
rect 153476 357468 153528 357474
rect 153476 357410 153528 357416
rect 153488 350606 153516 357410
rect 153476 350600 153528 350606
rect 153476 350542 153528 350548
rect 153384 350532 153436 350538
rect 153384 350474 153436 350480
rect 153396 341018 153424 350474
rect 153384 341012 153436 341018
rect 153384 340954 153436 340960
rect 153384 340468 153436 340474
rect 153384 340410 153436 340416
rect 153396 331242 153424 340410
rect 153396 331214 153516 331242
rect 153488 318850 153516 331214
rect 153384 318844 153436 318850
rect 153384 318786 153436 318792
rect 153476 318844 153528 318850
rect 153476 318786 153528 318792
rect 153396 311982 153424 318786
rect 153384 311976 153436 311982
rect 153384 311918 153436 311924
rect 153476 311976 153528 311982
rect 153476 311918 153528 311924
rect 153488 302258 153516 311918
rect 153292 302252 153344 302258
rect 153292 302194 153344 302200
rect 153476 302252 153528 302258
rect 153476 302194 153528 302200
rect 153304 302138 153332 302194
rect 153304 302110 153424 302138
rect 153396 292618 153424 302110
rect 153396 292590 153516 292618
rect 153488 282946 153516 292590
rect 153292 282940 153344 282946
rect 153292 282882 153344 282888
rect 153476 282940 153528 282946
rect 153476 282882 153528 282888
rect 153304 282826 153332 282882
rect 153304 282798 153424 282826
rect 153396 280158 153424 282798
rect 153384 280152 153436 280158
rect 153384 280094 153436 280100
rect 153568 273284 153620 273290
rect 153568 273226 153620 273232
rect 153580 270502 153608 273226
rect 153568 270496 153620 270502
rect 153568 270438 153620 270444
rect 153660 260908 153712 260914
rect 153660 260850 153712 260856
rect 153672 254046 153700 260850
rect 153660 254040 153712 254046
rect 153660 253982 153712 253988
rect 153568 253904 153620 253910
rect 153568 253846 153620 253852
rect 153580 244202 153608 253846
rect 153396 244174 153608 244202
rect 153396 241482 153424 244174
rect 153304 241454 153424 241482
rect 153304 234734 153332 241454
rect 153292 234728 153344 234734
rect 153292 234670 153344 234676
rect 153292 234592 153344 234598
rect 153292 234534 153344 234540
rect 153304 231826 153332 234534
rect 153212 231798 153332 231826
rect 153212 225010 153240 231798
rect 153200 225004 153252 225010
rect 153200 224946 153252 224952
rect 153200 222216 153252 222222
rect 153200 222158 153252 222164
rect 153212 215354 153240 222158
rect 153200 215348 153252 215354
rect 153200 215290 153252 215296
rect 153292 215212 153344 215218
rect 153292 215154 153344 215160
rect 153304 212498 153332 215154
rect 153292 212492 153344 212498
rect 153292 212434 153344 212440
rect 153384 202904 153436 202910
rect 153384 202846 153436 202852
rect 151084 202224 151136 202230
rect 151084 202166 151136 202172
rect 146944 202156 146996 202162
rect 146944 202098 146996 202104
rect 145564 201272 145616 201278
rect 145564 201214 145616 201220
rect 153396 201210 153424 202846
rect 153856 202366 153884 518298
rect 157996 202434 158024 553454
rect 160744 532772 160796 532778
rect 160744 532714 160796 532720
rect 159364 518288 159416 518294
rect 159364 518230 159416 518236
rect 159376 202570 159404 518230
rect 159364 202564 159416 202570
rect 159364 202506 159416 202512
rect 160756 202502 160784 532714
rect 162136 202842 162164 553862
rect 175936 398138 175964 583646
rect 270408 583636 270460 583642
rect 270408 583578 270460 583584
rect 195888 562012 195940 562018
rect 195888 561954 195940 561960
rect 192484 506524 192536 506530
rect 192484 506466 192536 506472
rect 175924 398132 175976 398138
rect 175924 398074 175976 398080
rect 168656 395616 168708 395622
rect 168656 395558 168708 395564
rect 162124 202836 162176 202842
rect 162124 202778 162176 202784
rect 160744 202496 160796 202502
rect 160744 202438 160796 202444
rect 157984 202428 158036 202434
rect 157984 202370 158036 202376
rect 153844 202360 153896 202366
rect 153844 202302 153896 202308
rect 168380 202292 168432 202298
rect 168380 202234 168432 202240
rect 153384 201204 153436 201210
rect 153384 201146 153436 201152
rect 168392 200002 168420 202234
rect 168668 200002 168696 395558
rect 179512 395548 179564 395554
rect 179512 395490 179564 395496
rect 169116 202836 169168 202842
rect 169116 202778 169168 202784
rect 169128 200002 169156 202778
rect 176936 202564 176988 202570
rect 176936 202506 176988 202512
rect 176948 200002 176976 202506
rect 178040 202496 178092 202502
rect 178040 202438 178092 202444
rect 178052 200002 178080 202438
rect 178684 202156 178736 202162
rect 178684 202098 178736 202104
rect 178696 200002 178724 202098
rect 179524 200002 179552 395490
rect 192496 342922 192524 506466
rect 195704 409488 195756 409494
rect 195704 409430 195756 409436
rect 195612 409216 195664 409222
rect 195612 409158 195664 409164
rect 195520 409148 195572 409154
rect 195520 409090 195572 409096
rect 192484 342916 192536 342922
rect 192484 342858 192536 342864
rect 195532 205018 195560 409090
rect 195520 205012 195572 205018
rect 195520 204954 195572 204960
rect 195624 204950 195652 409158
rect 195716 205154 195744 409430
rect 195796 409420 195848 409426
rect 195796 409362 195848 409368
rect 195704 205148 195756 205154
rect 195704 205090 195756 205096
rect 195808 205086 195836 409362
rect 195900 205222 195928 561954
rect 197084 561944 197136 561950
rect 197084 561886 197136 561892
rect 208676 561944 208728 561950
rect 208676 561886 208728 561892
rect 217876 561944 217928 561950
rect 217876 561886 217928 561892
rect 196992 561876 197044 561882
rect 196992 561818 197044 561824
rect 196900 410168 196952 410174
rect 196900 410110 196952 410116
rect 196808 409556 196860 409562
rect 196808 409498 196860 409504
rect 196716 409352 196768 409358
rect 196716 409294 196768 409300
rect 196624 409284 196676 409290
rect 196624 409226 196676 409232
rect 196636 205290 196664 409226
rect 196728 205358 196756 409294
rect 196716 205352 196768 205358
rect 196716 205294 196768 205300
rect 196624 205284 196676 205290
rect 196624 205226 196676 205232
rect 195888 205216 195940 205222
rect 195888 205158 195940 205164
rect 195796 205080 195848 205086
rect 195796 205022 195848 205028
rect 195612 204944 195664 204950
rect 195612 204886 195664 204892
rect 182180 202428 182232 202434
rect 182180 202370 182232 202376
rect 181260 202360 181312 202366
rect 181260 202302 181312 202308
rect 180340 202224 180392 202230
rect 180340 202166 180392 202172
rect 180352 200002 180380 202166
rect 181272 200002 181300 202302
rect 182192 200002 182220 202370
rect 196820 201822 196848 409498
rect 196912 202774 196940 410110
rect 196900 202768 196952 202774
rect 197004 202745 197032 561818
rect 197096 202881 197124 561886
rect 205548 561876 205600 561882
rect 205548 561818 205600 561824
rect 197268 561808 197320 561814
rect 197268 561750 197320 561756
rect 197176 560244 197228 560250
rect 197176 560186 197228 560192
rect 197082 202872 197138 202881
rect 197082 202807 197138 202816
rect 196900 202710 196952 202716
rect 196990 202736 197046 202745
rect 196990 202671 197046 202680
rect 197188 202201 197216 560186
rect 197280 202473 197308 561750
rect 202052 560244 202104 560250
rect 202052 560186 202104 560192
rect 202064 559994 202092 560186
rect 202064 559966 202446 559994
rect 205560 559980 205588 561818
rect 208688 559980 208716 561886
rect 214748 561808 214800 561814
rect 211618 561776 211674 561785
rect 214748 561750 214800 561756
rect 211618 561711 211674 561720
rect 211632 559980 211660 561711
rect 214760 559980 214788 561750
rect 217888 559980 217916 561886
rect 222198 556200 222254 556209
rect 222198 556135 222254 556144
rect 198646 534168 198702 534177
rect 198646 534103 198702 534112
rect 198554 524648 198610 524657
rect 198554 524583 198610 524592
rect 198280 521008 198332 521014
rect 198280 520950 198332 520956
rect 198188 520940 198240 520946
rect 198188 520882 198240 520888
rect 198096 518288 198148 518294
rect 198096 518230 198148 518236
rect 198004 407244 198056 407250
rect 198004 407186 198056 407192
rect 197728 406564 197780 406570
rect 197728 406506 197780 406512
rect 197740 365702 197768 406506
rect 198016 397458 198044 407186
rect 198004 397452 198056 397458
rect 198004 397394 198056 397400
rect 198002 378720 198058 378729
rect 198002 378655 198058 378664
rect 197910 374368 197966 374377
rect 197910 374303 197966 374312
rect 197818 370288 197874 370297
rect 197818 370223 197874 370232
rect 197728 365696 197780 365702
rect 197728 365638 197780 365644
rect 197726 361856 197782 361865
rect 197726 361791 197782 361800
rect 197542 357504 197598 357513
rect 197542 357439 197598 357448
rect 197450 353424 197506 353433
rect 197450 353359 197506 353368
rect 197358 349072 197414 349081
rect 197358 349007 197414 349016
rect 197372 202502 197400 349007
rect 197464 203726 197492 353359
rect 197452 203720 197504 203726
rect 197452 203662 197504 203668
rect 197556 202570 197584 357439
rect 197634 344992 197690 345001
rect 197634 344927 197690 344936
rect 197648 202638 197676 344927
rect 197740 203930 197768 361791
rect 197728 203924 197780 203930
rect 197728 203866 197780 203872
rect 197832 203658 197860 370223
rect 197820 203652 197872 203658
rect 197820 203594 197872 203600
rect 197636 202632 197688 202638
rect 197636 202574 197688 202580
rect 197544 202564 197596 202570
rect 197544 202506 197596 202512
rect 197360 202496 197412 202502
rect 197266 202464 197322 202473
rect 197360 202438 197412 202444
rect 197266 202399 197322 202408
rect 197174 202192 197230 202201
rect 197924 202162 197952 374303
rect 198016 203862 198044 378655
rect 198108 339046 198136 518230
rect 198096 339040 198148 339046
rect 198096 338982 198148 338988
rect 198200 338774 198228 520882
rect 198292 338842 198320 520950
rect 198462 399664 198518 399673
rect 198462 399599 198518 399608
rect 198370 387152 198426 387161
rect 198370 387087 198426 387096
rect 198280 338836 198332 338842
rect 198280 338778 198332 338784
rect 198188 338768 198240 338774
rect 198188 338710 198240 338716
rect 198004 203856 198056 203862
rect 198004 203798 198056 203804
rect 198384 203590 198412 387087
rect 198476 203794 198504 399599
rect 198464 203788 198516 203794
rect 198464 203730 198516 203736
rect 198372 203584 198424 203590
rect 198372 203526 198424 203532
rect 197174 202127 197230 202136
rect 197912 202156 197964 202162
rect 197912 202098 197964 202104
rect 196808 201816 196860 201822
rect 196808 201758 196860 201764
rect 198568 201550 198596 524583
rect 198660 201958 198688 534103
rect 198738 529272 198794 529281
rect 198738 529207 198794 529216
rect 198648 201952 198700 201958
rect 198648 201894 198700 201900
rect 198752 201890 198780 529207
rect 199384 521144 199436 521150
rect 199384 521086 199436 521092
rect 198830 403744 198886 403753
rect 198830 403679 198886 403688
rect 198844 202230 198872 403679
rect 198922 395312 198978 395321
rect 198922 395247 198978 395256
rect 198832 202224 198884 202230
rect 198832 202166 198884 202172
rect 198936 202094 198964 395247
rect 199014 391232 199070 391241
rect 199014 391167 199070 391176
rect 199028 203998 199056 391167
rect 199106 382800 199162 382809
rect 199106 382735 199162 382744
rect 199016 203992 199068 203998
rect 199016 203934 199068 203940
rect 199120 202842 199148 382735
rect 199198 365936 199254 365945
rect 199198 365871 199254 365880
rect 199108 202836 199160 202842
rect 199108 202778 199160 202784
rect 199212 202434 199240 365871
rect 199292 342916 199344 342922
rect 199292 342858 199344 342864
rect 199200 202428 199252 202434
rect 199200 202370 199252 202376
rect 198924 202088 198976 202094
rect 198924 202030 198976 202036
rect 198740 201884 198792 201890
rect 198740 201826 198792 201832
rect 199304 201754 199332 342858
rect 199396 338910 199424 521086
rect 199476 521076 199528 521082
rect 199476 521018 199528 521024
rect 199488 338978 199516 521018
rect 200224 520118 200606 520146
rect 202892 520118 203550 520146
rect 199752 410100 199804 410106
rect 199752 410042 199804 410048
rect 199568 409692 199620 409698
rect 199568 409634 199620 409640
rect 199476 338972 199528 338978
rect 199476 338914 199528 338920
rect 199384 338904 199436 338910
rect 199384 338846 199436 338852
rect 199292 201748 199344 201754
rect 199292 201690 199344 201696
rect 199580 201686 199608 409634
rect 199660 409624 199712 409630
rect 199660 409566 199712 409572
rect 199568 201680 199620 201686
rect 199568 201622 199620 201628
rect 199672 201618 199700 409566
rect 199764 202026 199792 410042
rect 199936 410032 199988 410038
rect 199936 409974 199988 409980
rect 199844 409896 199896 409902
rect 199844 409838 199896 409844
rect 199856 202706 199884 409838
rect 199844 202700 199896 202706
rect 199844 202642 199896 202648
rect 199948 202094 199976 409974
rect 200028 409964 200080 409970
rect 200028 409906 200080 409912
rect 200040 202842 200068 409906
rect 200224 342922 200252 520118
rect 200580 410168 200632 410174
rect 200580 410110 200632 410116
rect 200592 408748 200620 410110
rect 202892 409698 202920 520118
rect 206664 517546 206692 520132
rect 205640 517540 205692 517546
rect 205640 517482 205692 517488
rect 206652 517540 206704 517546
rect 206652 517482 206704 517488
rect 203338 410408 203394 410417
rect 203338 410343 203394 410352
rect 202880 409692 202932 409698
rect 202880 409634 202932 409640
rect 203352 408748 203380 410343
rect 205652 409630 205680 517482
rect 206284 410440 206336 410446
rect 206284 410382 206336 410388
rect 205640 409624 205692 409630
rect 205640 409566 205692 409572
rect 206296 408748 206324 410382
rect 209044 409896 209096 409902
rect 209044 409838 209096 409844
rect 209056 408748 209084 409838
rect 209792 409562 209820 520132
rect 212552 520118 212934 520146
rect 215312 520118 216062 520146
rect 211988 410508 212040 410514
rect 211988 410450 212040 410456
rect 209780 409556 209832 409562
rect 209780 409498 209832 409504
rect 212000 408748 212028 410450
rect 212552 409494 212580 520118
rect 214748 409964 214800 409970
rect 214748 409906 214800 409912
rect 212540 409488 212592 409494
rect 212540 409430 212592 409436
rect 214760 408748 214788 409906
rect 215312 409426 215340 520118
rect 218992 518294 219020 520132
rect 218980 518288 219032 518294
rect 218980 518230 219032 518236
rect 217692 410100 217744 410106
rect 217692 410042 217744 410048
rect 215300 409420 215352 409426
rect 215300 409362 215352 409368
rect 217704 408748 217732 410042
rect 220452 410032 220504 410038
rect 220452 409974 220504 409980
rect 220464 408748 220492 409974
rect 222212 409222 222240 556135
rect 222290 552120 222346 552129
rect 222290 552055 222346 552064
rect 222200 409216 222252 409222
rect 222200 409158 222252 409164
rect 222304 409154 222332 552055
rect 222566 546952 222622 546961
rect 222566 546887 222622 546896
rect 222474 542600 222530 542609
rect 222474 542535 222530 542544
rect 222382 538384 222438 538393
rect 222382 538319 222438 538328
rect 222396 521150 222424 538319
rect 222384 521144 222436 521150
rect 222384 521086 222436 521092
rect 222488 520946 222516 542535
rect 222580 521082 222608 546887
rect 222658 533352 222714 533361
rect 222658 533287 222714 533296
rect 222568 521076 222620 521082
rect 222568 521018 222620 521024
rect 222672 521014 222700 533287
rect 222750 529000 222806 529009
rect 222750 528935 222806 528944
rect 222660 521008 222712 521014
rect 222660 520950 222712 520956
rect 222476 520940 222528 520946
rect 222476 520882 222528 520888
rect 222764 409358 222792 528935
rect 222842 524512 222898 524521
rect 222842 524447 222898 524456
rect 222752 409352 222804 409358
rect 222752 409294 222804 409300
rect 222856 409290 222884 524447
rect 267280 451376 267332 451382
rect 267280 451318 267332 451324
rect 248972 410848 249024 410854
rect 248972 410790 249024 410796
rect 266544 410848 266596 410854
rect 266544 410790 266596 410796
rect 246028 410780 246080 410786
rect 246028 410722 246080 410728
rect 234620 410712 234672 410718
rect 234620 410654 234672 410660
rect 228916 410644 228968 410650
rect 228916 410586 228968 410592
rect 223396 410576 223448 410582
rect 223396 410518 223448 410524
rect 222844 409284 222896 409290
rect 222844 409226 222896 409232
rect 222292 409148 222344 409154
rect 222292 409090 222344 409096
rect 223408 408748 223436 410518
rect 226154 410136 226210 410145
rect 226154 410071 226210 410080
rect 226168 408748 226196 410071
rect 228928 408748 228956 410586
rect 231858 410272 231914 410281
rect 231858 410207 231914 410216
rect 231872 408748 231900 410207
rect 234632 408748 234660 410654
rect 243268 410372 243320 410378
rect 243268 410314 243320 410320
rect 240324 410304 240376 410310
rect 240324 410246 240376 410252
rect 237564 410236 237616 410242
rect 237564 410178 237616 410184
rect 237576 408748 237604 410178
rect 240336 408748 240364 410246
rect 243280 408748 243308 410314
rect 246040 408748 246068 410722
rect 248984 408748 249012 410790
rect 266360 410440 266412 410446
rect 266360 410382 266412 410388
rect 257436 410168 257488 410174
rect 257436 410110 257488 410116
rect 254676 410100 254728 410106
rect 254676 410042 254728 410048
rect 251732 410032 251784 410038
rect 251732 409974 251784 409980
rect 251744 408748 251772 409974
rect 254688 408748 254716 410042
rect 257448 408748 257476 410110
rect 263138 410000 263194 410009
rect 260380 409964 260432 409970
rect 263138 409935 263194 409944
rect 260380 409906 260432 409912
rect 260392 408748 260420 409906
rect 263152 408748 263180 409935
rect 265900 409896 265952 409902
rect 265900 409838 265952 409844
rect 265912 408748 265940 409838
rect 200212 342916 200264 342922
rect 200212 342858 200264 342864
rect 200592 337822 200620 340068
rect 203352 337890 203380 340068
rect 203340 337884 203392 337890
rect 203340 337826 203392 337832
rect 200580 337816 200632 337822
rect 200580 337758 200632 337764
rect 206112 337686 206140 340068
rect 209056 337958 209084 340068
rect 211830 340054 212488 340082
rect 209964 339040 210016 339046
rect 209964 338982 210016 338988
rect 209044 337952 209096 337958
rect 209044 337894 209096 337900
rect 206100 337680 206152 337686
rect 206100 337622 206152 337628
rect 209976 328506 210004 338982
rect 209780 328500 209832 328506
rect 209780 328442 209832 328448
rect 209964 328500 210016 328506
rect 209964 328442 210016 328448
rect 209792 318782 209820 328442
rect 209780 318776 209832 318782
rect 209780 318718 209832 318724
rect 209780 309188 209832 309194
rect 209780 309130 209832 309136
rect 209792 299470 209820 309130
rect 209780 299464 209832 299470
rect 209780 299406 209832 299412
rect 209780 289876 209832 289882
rect 209780 289818 209832 289824
rect 209792 280158 209820 289818
rect 209780 280152 209832 280158
rect 209780 280094 209832 280100
rect 209780 270564 209832 270570
rect 209780 270506 209832 270512
rect 209792 260846 209820 270506
rect 209780 260840 209832 260846
rect 209780 260782 209832 260788
rect 209780 251320 209832 251326
rect 209780 251262 209832 251268
rect 209792 241505 209820 251262
rect 209778 241496 209834 241505
rect 209778 241431 209834 241440
rect 209962 241496 210018 241505
rect 209962 241431 210018 241440
rect 209976 231878 210004 241431
rect 209780 231872 209832 231878
rect 209780 231814 209832 231820
rect 209964 231872 210016 231878
rect 209964 231814 210016 231820
rect 209792 222193 209820 231814
rect 209778 222184 209834 222193
rect 209778 222119 209834 222128
rect 209962 222184 210018 222193
rect 209962 222119 210018 222128
rect 209976 212566 210004 222119
rect 209780 212560 209832 212566
rect 209780 212502 209832 212508
rect 209964 212560 210016 212566
rect 209964 212502 210016 212508
rect 209792 202858 209820 212502
rect 200028 202836 200080 202842
rect 209792 202830 209912 202858
rect 200028 202778 200080 202784
rect 199936 202088 199988 202094
rect 199936 202030 199988 202036
rect 199752 202020 199804 202026
rect 199752 201962 199804 201968
rect 199660 201612 199712 201618
rect 199660 201554 199712 201560
rect 198556 201544 198608 201550
rect 198556 201486 198608 201492
rect 202880 201544 202932 201550
rect 202880 201486 202932 201492
rect 202892 200002 202920 201486
rect 209884 200258 209912 202830
rect 211712 201884 211764 201890
rect 211712 201826 211764 201832
rect 211158 201648 211214 201657
rect 211158 201583 211214 201592
rect 209872 200252 209924 200258
rect 209872 200194 209924 200200
rect 210286 200252 210338 200258
rect 210286 200194 210338 200200
rect 134168 199974 134228 200002
rect 134352 199974 134596 200002
rect 134720 199974 135056 200002
rect 142540 199974 142876 200002
rect 168392 199974 168544 200002
rect 168668 199974 169004 200002
rect 169128 199974 169372 200002
rect 176948 199974 177192 200002
rect 178052 199974 178112 200002
rect 178696 199974 178940 200002
rect 179524 199974 179860 200002
rect 180352 199974 180688 200002
rect 181272 199974 181608 200002
rect 182192 199974 182436 200002
rect 202860 199974 202920 200002
rect 210298 199988 210326 200194
rect 211172 200002 211200 201583
rect 211140 199974 211200 200002
rect 211724 200002 211752 201826
rect 212460 201550 212488 340054
rect 214104 338972 214156 338978
rect 214104 338914 214156 338920
rect 214116 338042 214144 338914
rect 214024 338014 214144 338042
rect 214024 331362 214052 338014
rect 214760 337754 214788 340068
rect 215300 338904 215352 338910
rect 215300 338846 215352 338852
rect 214748 337748 214800 337754
rect 214748 337690 214800 337696
rect 214012 331356 214064 331362
rect 214012 331298 214064 331304
rect 213920 328500 213972 328506
rect 213920 328442 213972 328448
rect 212538 201920 212594 201929
rect 212538 201855 212594 201864
rect 212448 201544 212500 201550
rect 212448 201486 212500 201492
rect 212552 200002 212580 201855
rect 213458 201784 213514 201793
rect 213458 201719 213514 201728
rect 213472 200002 213500 201719
rect 213932 200258 213960 328442
rect 213920 200252 213972 200258
rect 213920 200194 213972 200200
rect 214610 200252 214662 200258
rect 214610 200194 214662 200200
rect 211724 199974 211968 200002
rect 212552 199974 212888 200002
rect 213472 199974 213716 200002
rect 214622 199988 214650 200194
rect 215312 200002 215340 338846
rect 217520 337890 217548 340068
rect 220464 338026 220492 340068
rect 220820 338836 220872 338842
rect 220820 338778 220872 338784
rect 220452 338020 220504 338026
rect 220452 337962 220504 337968
rect 220084 337952 220136 337958
rect 220084 337894 220136 337900
rect 215944 337884 215996 337890
rect 215944 337826 215996 337832
rect 217508 337884 217560 337890
rect 217508 337826 217560 337832
rect 215956 201890 215984 337826
rect 218058 202056 218114 202065
rect 218058 201991 218114 202000
rect 216036 201952 216088 201958
rect 216036 201894 216088 201900
rect 215944 201884 215996 201890
rect 215944 201826 215996 201832
rect 216048 200002 216076 201894
rect 216864 201612 216916 201618
rect 216864 201554 216916 201560
rect 216876 200002 216904 201554
rect 218072 200002 218100 201991
rect 219532 201748 219584 201754
rect 219532 201690 219584 201696
rect 218612 201680 218664 201686
rect 218612 201622 218664 201628
rect 218624 200002 218652 201622
rect 219544 200002 219572 201690
rect 220096 201550 220124 337894
rect 220358 202872 220414 202881
rect 220358 202807 220414 202816
rect 220084 201544 220136 201550
rect 220084 201486 220136 201492
rect 220372 200002 220400 202807
rect 220832 201822 220860 338778
rect 222200 338768 222252 338774
rect 222200 338710 222252 338716
rect 220820 201816 220872 201822
rect 220820 201758 220872 201764
rect 221280 201816 221332 201822
rect 221280 201758 221332 201764
rect 221292 200002 221320 201758
rect 222212 200002 222240 338710
rect 223224 336870 223252 340068
rect 226168 337958 226196 340068
rect 226156 337952 226208 337958
rect 226156 337894 226208 337900
rect 228928 337278 228956 340068
rect 231872 337346 231900 340068
rect 234632 337822 234660 340068
rect 237288 338768 237340 338774
rect 237194 338736 237250 338745
rect 237288 338710 237340 338716
rect 237194 338671 237250 338680
rect 234620 337816 234672 337822
rect 234620 337758 234672 337764
rect 231860 337340 231912 337346
rect 231860 337282 231912 337288
rect 228916 337272 228968 337278
rect 228916 337214 228968 337220
rect 232504 337272 232556 337278
rect 232504 337214 232556 337220
rect 223212 336864 223264 336870
rect 223212 336806 223264 336812
rect 229744 336864 229796 336870
rect 229744 336806 229796 336812
rect 226892 205352 226944 205358
rect 226892 205294 226944 205300
rect 223854 202736 223910 202745
rect 223854 202671 223910 202680
rect 223028 201748 223080 201754
rect 223028 201690 223080 201696
rect 223040 200002 223068 201690
rect 223868 200002 223896 202671
rect 225142 202600 225198 202609
rect 225142 202535 225198 202544
rect 225156 200002 225184 202535
rect 226338 202464 226394 202473
rect 226338 202399 226394 202408
rect 226352 200002 226380 202399
rect 215312 199974 215464 200002
rect 216048 199974 216384 200002
rect 216876 199974 217212 200002
rect 218072 199974 218132 200002
rect 218624 199974 218960 200002
rect 219544 199974 219880 200002
rect 220372 199974 220708 200002
rect 221292 199974 221536 200002
rect 222212 199974 222456 200002
rect 223040 199974 223284 200002
rect 223868 199974 224204 200002
rect 225156 199974 225492 200002
rect 226320 199974 226380 200002
rect 226904 200002 226932 205294
rect 227904 205284 227956 205290
rect 227904 205226 227956 205232
rect 227916 200002 227944 205226
rect 228640 205216 228692 205222
rect 228640 205158 228692 205164
rect 228652 200002 228680 205158
rect 229560 205148 229612 205154
rect 229560 205090 229612 205096
rect 229100 202088 229152 202094
rect 229100 202030 229152 202036
rect 229112 201822 229140 202030
rect 229100 201816 229152 201822
rect 229100 201758 229152 201764
rect 229572 200002 229600 205090
rect 229756 201686 229784 336806
rect 230480 205080 230532 205086
rect 230480 205022 230532 205028
rect 229744 201680 229796 201686
rect 229744 201622 229796 201628
rect 230492 200002 230520 205022
rect 231216 205012 231268 205018
rect 231216 204954 231268 204960
rect 231228 200002 231256 204954
rect 232134 202328 232190 202337
rect 232134 202263 232190 202272
rect 232148 200002 232176 202263
rect 232410 201920 232466 201929
rect 232410 201855 232466 201864
rect 232424 201822 232452 201855
rect 232516 201822 232544 337214
rect 233240 204944 233292 204950
rect 233240 204886 233292 204892
rect 232412 201816 232464 201822
rect 232412 201758 232464 201764
rect 232504 201816 232556 201822
rect 232504 201758 232556 201764
rect 233252 200002 233280 204886
rect 233422 202192 233478 202201
rect 233422 202127 233478 202136
rect 233436 200002 233464 202127
rect 236644 202020 236696 202026
rect 236644 201962 236696 201968
rect 236656 200002 236684 201962
rect 236736 201816 236788 201822
rect 236736 201758 236788 201764
rect 226904 199974 227240 200002
rect 227916 199974 228068 200002
rect 228652 199974 228988 200002
rect 229572 199974 229816 200002
rect 230492 199974 230736 200002
rect 231228 199974 231564 200002
rect 232148 199974 232484 200002
rect 233252 199974 233312 200002
rect 233436 199974 233772 200002
rect 236348 199974 236684 200002
rect 236748 200002 236776 201758
rect 237208 200002 237236 338671
rect 237300 202026 237328 338710
rect 237576 337278 237604 340068
rect 240152 340054 240350 340082
rect 238116 338020 238168 338026
rect 238116 337962 238168 337968
rect 237748 337816 237800 337822
rect 237748 337758 237800 337764
rect 237564 337272 237616 337278
rect 237564 337214 237616 337220
rect 237288 202020 237340 202026
rect 237288 201962 237340 201968
rect 237380 201680 237432 201686
rect 237380 201622 237432 201628
rect 237392 200002 237420 201622
rect 237760 200002 237788 337758
rect 238024 337204 238076 337210
rect 238024 337146 238076 337152
rect 238036 201686 238064 337146
rect 238128 201822 238156 337962
rect 240048 337816 240100 337822
rect 240048 337758 240100 337764
rect 238760 203992 238812 203998
rect 238760 203934 238812 203940
rect 238668 202020 238720 202026
rect 238668 201962 238720 201968
rect 238680 201929 238708 201962
rect 238666 201920 238722 201929
rect 238666 201855 238722 201864
rect 238116 201816 238168 201822
rect 238116 201758 238168 201764
rect 238024 201680 238076 201686
rect 238024 201622 238076 201628
rect 238208 201612 238260 201618
rect 238208 201554 238260 201560
rect 238220 200002 238248 201554
rect 236748 199974 236808 200002
rect 237208 199974 237268 200002
rect 237392 199974 237636 200002
rect 237760 199974 238096 200002
rect 238220 199974 238556 200002
rect 238772 199918 238800 203934
rect 239680 202836 239732 202842
rect 239680 202778 239732 202784
rect 239220 201952 239272 201958
rect 239220 201894 239272 201900
rect 239232 200002 239260 201894
rect 239692 200002 239720 202778
rect 240060 201958 240088 337758
rect 240152 202842 240180 340054
rect 241428 337884 241480 337890
rect 241428 337826 241480 337832
rect 241440 202842 241468 337826
rect 243096 337822 243124 340068
rect 244188 338836 244240 338842
rect 244188 338778 244240 338784
rect 243084 337816 243136 337822
rect 243084 337758 243136 337764
rect 243084 337272 243136 337278
rect 243084 337214 243136 337220
rect 240140 202836 240192 202842
rect 240140 202778 240192 202784
rect 240508 202836 240560 202842
rect 240508 202778 240560 202784
rect 241428 202836 241480 202842
rect 241428 202778 241480 202784
rect 242992 202836 243044 202842
rect 242992 202778 243044 202784
rect 240048 201952 240100 201958
rect 240048 201894 240100 201900
rect 240520 200002 240548 202778
rect 241520 202768 241572 202774
rect 241520 202710 241572 202716
rect 240968 202088 241020 202094
rect 240968 202030 241020 202036
rect 240980 200002 241008 202030
rect 241060 202020 241112 202026
rect 241060 201962 241112 201968
rect 238924 199974 239260 200002
rect 239384 199974 239720 200002
rect 240304 199974 240548 200002
rect 240672 199974 241008 200002
rect 241072 200002 241100 201962
rect 241532 200002 241560 202710
rect 242072 201952 242124 201958
rect 242072 201894 242124 201900
rect 242084 200002 242112 201894
rect 242164 201884 242216 201890
rect 242164 201826 242216 201832
rect 241072 199974 241132 200002
rect 241532 199974 241592 200002
rect 242052 199974 242112 200002
rect 242176 200002 242204 201826
rect 243004 200002 243032 202778
rect 242176 199974 242420 200002
rect 242880 199974 243032 200002
rect 243096 199918 243124 337214
rect 244096 336864 244148 336870
rect 244096 336806 244148 336812
rect 244004 209772 244056 209778
rect 244004 209714 244056 209720
rect 243176 201748 243228 201754
rect 243176 201690 243228 201696
rect 243188 200002 243216 201690
rect 244016 200002 244044 209714
rect 244108 202842 244136 336806
rect 244200 209778 244228 338778
rect 244924 338020 244976 338026
rect 244924 337962 244976 337968
rect 244188 209772 244240 209778
rect 244188 209714 244240 209720
rect 244096 202836 244148 202842
rect 244096 202778 244148 202784
rect 244740 202632 244792 202638
rect 244740 202574 244792 202580
rect 244648 202020 244700 202026
rect 244648 201962 244700 201968
rect 244660 200002 244688 201962
rect 243188 199974 243340 200002
rect 243708 199974 244044 200002
rect 244628 199974 244688 200002
rect 244752 200002 244780 202574
rect 244936 202502 244964 337962
rect 246040 337890 246068 340068
rect 248616 340054 248814 340082
rect 246028 337884 246080 337890
rect 246028 337826 246080 337832
rect 247684 337816 247736 337822
rect 247684 337758 247736 337764
rect 247592 203992 247644 203998
rect 247592 203934 247644 203940
rect 245200 202700 245252 202706
rect 245200 202642 245252 202648
rect 247500 202700 247552 202706
rect 247500 202642 247552 202648
rect 244924 202496 244976 202502
rect 244924 202438 244976 202444
rect 245212 200002 245240 202642
rect 245660 202564 245712 202570
rect 245660 202506 245712 202512
rect 245672 200002 245700 202506
rect 246028 202496 246080 202502
rect 246028 202438 246080 202444
rect 246040 200002 246068 202438
rect 246488 201544 246540 201550
rect 246488 201486 246540 201492
rect 246500 200002 246528 201486
rect 247512 200002 247540 202642
rect 244752 199974 245088 200002
rect 245212 199974 245456 200002
rect 245672 199974 245916 200002
rect 246040 199974 246376 200002
rect 246500 199974 246836 200002
rect 247204 199974 247540 200002
rect 247604 200002 247632 203934
rect 247696 201958 247724 337758
rect 248616 336870 248644 340054
rect 248696 337952 248748 337958
rect 248696 337894 248748 337900
rect 250996 337952 251048 337958
rect 250996 337894 251048 337900
rect 248604 336864 248656 336870
rect 248604 336806 248656 336812
rect 247684 201952 247736 201958
rect 247684 201894 247736 201900
rect 247776 201612 247828 201618
rect 247776 201554 247828 201560
rect 247788 200002 247816 201554
rect 248708 200002 248736 337894
rect 248788 337340 248840 337346
rect 248788 337282 248840 337288
rect 248800 202450 248828 337282
rect 250536 204060 250588 204066
rect 250536 204002 250588 204008
rect 250076 202496 250128 202502
rect 248800 202422 249288 202450
rect 250076 202438 250128 202444
rect 248972 202360 249024 202366
rect 248972 202302 249024 202308
rect 248984 200002 249012 202302
rect 247604 199974 247664 200002
rect 247788 199974 248124 200002
rect 248492 199974 248736 200002
rect 248952 199974 249012 200002
rect 249260 200002 249288 202422
rect 250088 200002 250116 202438
rect 250548 200002 250576 204002
rect 250904 202632 250956 202638
rect 250904 202574 250956 202580
rect 250916 200002 250944 202574
rect 251008 202502 251036 337894
rect 251744 337686 251772 340068
rect 253664 338904 253716 338910
rect 253664 338846 253716 338852
rect 251732 337680 251784 337686
rect 251732 337622 251784 337628
rect 252468 337680 252520 337686
rect 252468 337622 252520 337628
rect 251824 202836 251876 202842
rect 251824 202778 251876 202784
rect 250996 202496 251048 202502
rect 250996 202438 251048 202444
rect 251456 201544 251508 201550
rect 251456 201486 251508 201492
rect 251468 200002 251496 201486
rect 251836 200002 251864 202778
rect 252376 202768 252428 202774
rect 252376 202710 252428 202716
rect 251916 201884 251968 201890
rect 251916 201826 251968 201832
rect 249260 199974 249412 200002
rect 249872 199974 250116 200002
rect 250240 199974 250576 200002
rect 250700 199974 250944 200002
rect 251160 199974 251496 200002
rect 251620 199974 251864 200002
rect 251928 200002 251956 201826
rect 252388 200002 252416 202710
rect 252480 201754 252508 337622
rect 253572 204128 253624 204134
rect 253572 204070 253624 204076
rect 253112 201952 253164 201958
rect 253112 201894 253164 201900
rect 252468 201748 252520 201754
rect 252468 201690 252520 201696
rect 253124 200002 253152 201894
rect 253584 200002 253612 204070
rect 251928 199974 251988 200002
rect 252388 199974 252448 200002
rect 252908 199974 253152 200002
rect 253276 199974 253612 200002
rect 253676 200002 253704 338846
rect 253756 337884 253808 337890
rect 253756 337826 253808 337832
rect 253768 201958 253796 337826
rect 254504 336870 254532 340068
rect 257448 337822 257476 340068
rect 257712 338972 257764 338978
rect 257712 338914 257764 338920
rect 257436 337816 257488 337822
rect 257436 337758 257488 337764
rect 255320 337340 255372 337346
rect 255320 337282 255372 337288
rect 254492 336864 254544 336870
rect 254492 336806 254544 336812
rect 255332 212566 255360 337282
rect 257724 336734 257752 338914
rect 260208 337958 260236 340068
rect 262128 339176 262180 339182
rect 262128 339118 262180 339124
rect 260196 337952 260248 337958
rect 260196 337894 260248 337900
rect 258724 337748 258776 337754
rect 258724 337690 258776 337696
rect 258264 336864 258316 336870
rect 258264 336806 258316 336812
rect 257712 336728 257764 336734
rect 257712 336670 257764 336676
rect 257804 336728 257856 336734
rect 257804 336670 257856 336676
rect 257816 335306 257844 336670
rect 257804 335300 257856 335306
rect 257804 335242 257856 335248
rect 257712 317484 257764 317490
rect 257712 317426 257764 317432
rect 257724 317393 257752 317426
rect 257710 317384 257766 317393
rect 257710 317319 257766 317328
rect 257802 311808 257858 311817
rect 257802 311743 257858 311752
rect 257816 307766 257844 311743
rect 257804 307760 257856 307766
rect 257804 307702 257856 307708
rect 257896 298172 257948 298178
rect 257896 298114 257948 298120
rect 257908 288454 257936 298114
rect 257804 288448 257856 288454
rect 257804 288390 257856 288396
rect 257896 288448 257948 288454
rect 257896 288390 257948 288396
rect 257816 288318 257844 288390
rect 257804 288312 257856 288318
rect 257804 288254 257856 288260
rect 257896 278792 257948 278798
rect 257896 278734 257948 278740
rect 257908 273306 257936 278734
rect 257816 273278 257936 273306
rect 257816 270502 257844 273278
rect 257804 270496 257856 270502
rect 257804 270438 257856 270444
rect 257804 263560 257856 263566
rect 257804 263502 257856 263508
rect 257816 260846 257844 263502
rect 257804 260840 257856 260846
rect 257804 260782 257856 260788
rect 257804 253836 257856 253842
rect 257804 253778 257856 253784
rect 257816 251190 257844 253778
rect 257804 251184 257856 251190
rect 257804 251126 257856 251132
rect 257712 241528 257764 241534
rect 257712 241470 257764 241476
rect 257724 234666 257752 241470
rect 257712 234660 257764 234666
rect 257712 234602 257764 234608
rect 257804 234524 257856 234530
rect 257804 234466 257856 234472
rect 257816 225078 257844 234466
rect 257804 225072 257856 225078
rect 257804 225014 257856 225020
rect 257712 224936 257764 224942
rect 257712 224878 257764 224884
rect 257724 222086 257752 224878
rect 257712 222080 257764 222086
rect 257712 222022 257764 222028
rect 257988 222080 258040 222086
rect 257988 222022 258040 222028
rect 258000 220833 258028 222022
rect 257802 220824 257858 220833
rect 257802 220759 257858 220768
rect 257986 220824 258042 220833
rect 257986 220759 258042 220768
rect 255320 212560 255372 212566
rect 255320 212502 255372 212508
rect 256240 212560 256292 212566
rect 256240 212502 256292 212508
rect 255780 204196 255832 204202
rect 255780 204138 255832 204144
rect 254032 202428 254084 202434
rect 254032 202370 254084 202376
rect 253756 201952 253808 201958
rect 253756 201894 253808 201900
rect 254044 200002 254072 202370
rect 254860 201952 254912 201958
rect 254860 201894 254912 201900
rect 254872 200002 254900 201894
rect 255228 201612 255280 201618
rect 255228 201554 255280 201560
rect 255240 200002 255268 201554
rect 255792 200002 255820 204138
rect 256148 201884 256200 201890
rect 256148 201826 256200 201832
rect 256160 200002 256188 201826
rect 253676 199974 253736 200002
rect 254044 199974 254196 200002
rect 254656 199974 254900 200002
rect 255024 199974 255268 200002
rect 255484 199974 255820 200002
rect 255944 199974 256188 200002
rect 256252 200002 256280 212502
rect 257816 212242 257844 220759
rect 257816 212214 258028 212242
rect 257160 203924 257212 203930
rect 257160 203866 257212 203872
rect 257066 202192 257122 202201
rect 257066 202127 257122 202136
rect 257080 200002 257108 202127
rect 256252 199974 256404 200002
rect 256772 199974 257108 200002
rect 257172 200002 257200 203866
rect 258000 202910 258028 212214
rect 257712 202904 257764 202910
rect 257712 202846 257764 202852
rect 257988 202904 258040 202910
rect 257988 202846 258040 202852
rect 257724 200410 257752 202846
rect 258172 202292 258224 202298
rect 258172 202234 258224 202240
rect 258080 201476 258132 201482
rect 258080 201418 258132 201424
rect 257678 200382 257752 200410
rect 257172 199974 257232 200002
rect 257678 199988 257706 200382
rect 258092 200002 258120 201418
rect 258060 199974 258120 200002
rect 258184 200002 258212 202234
rect 258276 200138 258304 336806
rect 258736 201618 258764 337690
rect 260380 203856 260432 203862
rect 260380 203798 260432 203804
rect 260196 202428 260248 202434
rect 260196 202370 260248 202376
rect 259460 201680 259512 201686
rect 259460 201622 259512 201628
rect 260104 201680 260156 201686
rect 260104 201622 260156 201628
rect 258724 201612 258776 201618
rect 258724 201554 258776 201560
rect 258276 200110 258856 200138
rect 258828 200002 258856 200110
rect 259472 200002 259500 201622
rect 260116 200002 260144 201622
rect 258184 199974 258520 200002
rect 258828 199974 258980 200002
rect 259440 199974 259500 200002
rect 259808 199974 260144 200002
rect 260208 200002 260236 202370
rect 260392 200002 260420 203798
rect 262140 202366 262168 339118
rect 263152 337890 263180 340068
rect 265926 340054 266308 340082
rect 263140 337884 263192 337890
rect 263140 337826 263192 337832
rect 262772 203788 262824 203794
rect 262772 203730 262824 203736
rect 261668 202360 261720 202366
rect 261668 202302 261720 202308
rect 262128 202360 262180 202366
rect 262128 202302 262180 202308
rect 260840 201816 260892 201822
rect 260840 201758 260892 201764
rect 260852 200002 260880 201758
rect 261680 200002 261708 202302
rect 261944 202292 261996 202298
rect 261944 202234 261996 202240
rect 260208 199974 260268 200002
rect 260392 199974 260728 200002
rect 260852 199974 261188 200002
rect 261556 199974 261708 200002
rect 261956 200002 261984 202234
rect 262678 201648 262734 201657
rect 262678 201583 262734 201592
rect 262692 200002 262720 201583
rect 261956 199974 262016 200002
rect 262476 199974 262720 200002
rect 262784 200002 262812 203730
rect 262956 203720 263008 203726
rect 262956 203662 263008 203668
rect 262968 200002 262996 203662
rect 265256 203652 265308 203658
rect 265256 203594 265308 203600
rect 263600 201748 263652 201754
rect 263600 201690 263652 201696
rect 265164 201748 265216 201754
rect 265164 201690 265216 201696
rect 263612 200002 263640 201690
rect 263876 201612 263928 201618
rect 263876 201554 263928 201560
rect 263888 200002 263916 201554
rect 264888 201544 264940 201550
rect 264888 201486 264940 201492
rect 264900 200002 264928 201486
rect 265176 200002 265204 201690
rect 262784 199974 262844 200002
rect 262968 199974 263304 200002
rect 263612 199974 263764 200002
rect 263888 199974 264224 200002
rect 264592 199974 264928 200002
rect 265052 199974 265204 200002
rect 265268 200002 265296 203594
rect 266280 201822 266308 340054
rect 266268 201816 266320 201822
rect 266268 201758 266320 201764
rect 266174 201512 266230 201521
rect 266174 201447 266230 201456
rect 266188 200002 266216 201447
rect 266372 200138 266400 410382
rect 266452 410032 266504 410038
rect 266452 409974 266504 409980
rect 266464 201210 266492 409974
rect 266556 201550 266584 410790
rect 266636 410712 266688 410718
rect 266636 410654 266688 410660
rect 266648 202706 266676 410654
rect 267004 410644 267056 410650
rect 267004 410586 267056 410592
rect 266912 410576 266964 410582
rect 266912 410518 266964 410524
rect 266820 410372 266872 410378
rect 266820 410314 266872 410320
rect 266728 410304 266780 410310
rect 266728 410246 266780 410252
rect 266740 202842 266768 410246
rect 266728 202836 266780 202842
rect 266728 202778 266780 202784
rect 266636 202700 266688 202706
rect 266636 202642 266688 202648
rect 266832 202366 266860 410314
rect 266820 202360 266872 202366
rect 266820 202302 266872 202308
rect 266924 201958 266952 410518
rect 266912 201952 266964 201958
rect 266912 201894 266964 201900
rect 267016 201618 267044 410586
rect 267096 410508 267148 410514
rect 267096 410450 267148 410456
rect 267108 201686 267136 410450
rect 267186 399664 267242 399673
rect 267186 399599 267242 399608
rect 267200 201754 267228 399599
rect 267292 385694 267320 451318
rect 267740 410780 267792 410786
rect 267740 410722 267792 410728
rect 267648 410236 267700 410242
rect 267648 410178 267700 410184
rect 267556 409964 267608 409970
rect 267556 409906 267608 409912
rect 267280 385688 267332 385694
rect 267280 385630 267332 385636
rect 267278 357504 267334 357513
rect 267278 357439 267334 357448
rect 267188 201748 267240 201754
rect 267188 201690 267240 201696
rect 267096 201680 267148 201686
rect 267096 201622 267148 201628
rect 267004 201612 267056 201618
rect 267004 201554 267056 201560
rect 267292 201550 267320 357439
rect 267370 353424 267426 353433
rect 267370 353359 267426 353368
rect 267384 202094 267412 353359
rect 267462 349072 267518 349081
rect 267462 349007 267518 349016
rect 267372 202088 267424 202094
rect 267372 202030 267424 202036
rect 267476 201890 267504 349007
rect 267568 338978 267596 409906
rect 267556 338972 267608 338978
rect 267556 338914 267608 338920
rect 267660 338774 267688 410178
rect 267648 338768 267700 338774
rect 267648 338710 267700 338716
rect 267556 203584 267608 203590
rect 267556 203526 267608 203532
rect 267464 201884 267516 201890
rect 267464 201826 267516 201832
rect 266544 201544 266596 201550
rect 266544 201486 266596 201492
rect 266636 201544 266688 201550
rect 266636 201486 266688 201492
rect 267280 201544 267332 201550
rect 267280 201486 267332 201492
rect 266452 201204 266504 201210
rect 266452 201146 266504 201152
rect 266372 200122 266492 200138
rect 266372 200116 266504 200122
rect 266372 200110 266452 200116
rect 266452 200058 266504 200064
rect 266464 200027 266492 200058
rect 265268 199974 265512 200002
rect 265972 199974 266216 200002
rect 238760 199912 238812 199918
rect 238760 199854 238812 199860
rect 239496 199912 239548 199918
rect 243084 199912 243136 199918
rect 239548 199860 239844 199866
rect 239496 199854 239844 199860
rect 243084 199854 243136 199860
rect 243820 199912 243872 199918
rect 266648 199866 266676 201486
rect 267568 200138 267596 203526
rect 267752 202570 267780 410722
rect 268752 410168 268804 410174
rect 268752 410110 268804 410116
rect 267830 403744 267886 403753
rect 267830 403679 267886 403688
rect 267844 202774 267872 403679
rect 267922 395312 267978 395321
rect 267922 395247 267978 395256
rect 267936 204066 267964 395247
rect 268014 391232 268070 391241
rect 268014 391167 268070 391176
rect 267924 204060 267976 204066
rect 267924 204002 267976 204008
rect 267832 202768 267884 202774
rect 267832 202710 267884 202716
rect 267740 202564 267792 202570
rect 267740 202506 267792 202512
rect 268028 202026 268056 391167
rect 268106 386880 268162 386889
rect 268106 386815 268162 386824
rect 268120 203998 268148 386815
rect 268198 382800 268254 382809
rect 268198 382735 268254 382744
rect 268212 204202 268240 382735
rect 268290 378448 268346 378457
rect 268290 378383 268346 378392
rect 268200 204196 268252 204202
rect 268200 204138 268252 204144
rect 268108 203992 268160 203998
rect 268108 203934 268160 203940
rect 268304 202638 268332 378383
rect 268382 374368 268438 374377
rect 268382 374303 268438 374312
rect 268292 202632 268344 202638
rect 268292 202574 268344 202580
rect 268396 202502 268424 374303
rect 268474 370016 268530 370025
rect 268474 369951 268530 369960
rect 268384 202496 268436 202502
rect 268384 202438 268436 202444
rect 268488 202434 268516 369951
rect 268566 365936 268622 365945
rect 268566 365871 268622 365880
rect 268476 202428 268528 202434
rect 268476 202370 268528 202376
rect 268580 202230 268608 365871
rect 268658 361584 268714 361593
rect 268658 361519 268714 361528
rect 268568 202224 268620 202230
rect 268568 202166 268620 202172
rect 268016 202020 268068 202026
rect 268016 201962 268068 201968
rect 268200 201680 268252 201686
rect 268200 201622 268252 201628
rect 267740 201612 267792 201618
rect 267740 201554 267792 201560
rect 267648 201204 267700 201210
rect 267648 201146 267700 201152
rect 266728 200116 266780 200122
rect 266728 200058 266780 200064
rect 267476 200110 267596 200138
rect 266740 200002 266768 200058
rect 267476 200002 267504 200110
rect 267660 200002 267688 201146
rect 266740 199974 266800 200002
rect 267260 199974 267504 200002
rect 267628 199974 267688 200002
rect 267752 200002 267780 201554
rect 268212 200002 268240 201622
rect 268672 200002 268700 361519
rect 268764 338842 268792 410110
rect 268844 410100 268896 410106
rect 268844 410042 268896 410048
rect 268856 338910 268884 410042
rect 268936 409896 268988 409902
rect 268936 409838 268988 409844
rect 268948 339182 268976 409838
rect 269026 344992 269082 345001
rect 269026 344927 269082 344936
rect 268936 339176 268988 339182
rect 268936 339118 268988 339124
rect 268844 338904 268896 338910
rect 268844 338846 268896 338852
rect 268752 338836 268804 338842
rect 268752 338778 268804 338784
rect 269040 204134 269068 344927
rect 269028 204128 269080 204134
rect 269028 204070 269080 204076
rect 269488 202156 269540 202162
rect 269488 202098 269540 202104
rect 269120 201816 269172 201822
rect 269120 201758 269172 201764
rect 269132 200002 269160 201758
rect 269500 200002 269528 202098
rect 270420 200002 270448 583578
rect 286324 583568 286376 583574
rect 286324 583510 286376 583516
rect 281356 583024 281408 583030
rect 281356 582966 281408 582972
rect 274546 582584 274602 582593
rect 274546 582519 274602 582528
rect 272524 569968 272576 569974
rect 272524 569910 272576 569916
rect 271788 203652 271840 203658
rect 271788 203594 271840 203600
rect 271420 202564 271472 202570
rect 271420 202506 271472 202512
rect 270960 202224 271012 202230
rect 270960 202166 271012 202172
rect 270972 200002 271000 202166
rect 271432 200002 271460 202506
rect 271800 200002 271828 203594
rect 272248 202836 272300 202842
rect 272248 202778 272300 202784
rect 272260 200002 272288 202778
rect 272536 202570 272564 569910
rect 273168 556232 273220 556238
rect 273168 556174 273220 556180
rect 273180 202842 273208 556174
rect 273168 202836 273220 202842
rect 273168 202778 273220 202784
rect 272524 202564 272576 202570
rect 272524 202506 272576 202512
rect 274560 202502 274588 582519
rect 280068 521688 280120 521694
rect 280068 521630 280120 521636
rect 279424 518968 279476 518974
rect 279424 518910 279476 518916
rect 277308 497276 277360 497282
rect 277308 497218 277360 497224
rect 276664 497208 276716 497214
rect 276664 497150 276716 497156
rect 273996 202496 274048 202502
rect 273996 202438 274048 202444
rect 274548 202496 274600 202502
rect 274548 202438 274600 202444
rect 273628 201680 273680 201686
rect 273628 201622 273680 201628
rect 273640 200002 273668 201622
rect 274008 200002 274036 202438
rect 275284 202428 275336 202434
rect 275284 202370 275336 202376
rect 275296 200002 275324 202370
rect 275744 202360 275796 202366
rect 275744 202302 275796 202308
rect 275756 200002 275784 202302
rect 276676 201686 276704 497150
rect 277320 202502 277348 497218
rect 279436 202502 279464 518910
rect 276940 202496 276992 202502
rect 276940 202438 276992 202444
rect 277308 202496 277360 202502
rect 277308 202438 277360 202444
rect 278688 202496 278740 202502
rect 278688 202438 278740 202444
rect 279424 202496 279476 202502
rect 279424 202438 279476 202444
rect 276664 201680 276716 201686
rect 276664 201622 276716 201628
rect 276952 200002 276980 202438
rect 277308 202292 277360 202298
rect 277308 202234 277360 202240
rect 277320 200002 277348 202234
rect 278700 200002 278728 202438
rect 280080 201618 280108 521630
rect 280528 203584 280580 203590
rect 280528 203526 280580 203532
rect 279240 201612 279292 201618
rect 279240 201554 279292 201560
rect 280068 201612 280120 201618
rect 280068 201554 280120 201560
rect 279252 200002 279280 201554
rect 280540 200002 280568 203526
rect 281368 202502 281396 582966
rect 284944 516180 284996 516186
rect 284944 516122 284996 516128
rect 284116 497820 284168 497826
rect 284116 497762 284168 497768
rect 280988 202496 281040 202502
rect 280988 202438 281040 202444
rect 281356 202496 281408 202502
rect 281356 202438 281408 202444
rect 281000 200002 281028 202438
rect 283564 202156 283616 202162
rect 283564 202098 283616 202104
rect 282644 201612 282696 201618
rect 282644 201554 282696 201560
rect 282276 201544 282328 201550
rect 282276 201486 282328 201492
rect 282288 200002 282316 201486
rect 282656 200002 282684 201554
rect 283576 200002 283604 202098
rect 284128 200138 284156 497762
rect 284208 497684 284260 497690
rect 284208 497626 284260 497632
rect 284036 200110 284156 200138
rect 284036 200002 284064 200110
rect 284220 200002 284248 497626
rect 284956 201550 284984 516122
rect 285588 497412 285640 497418
rect 285588 497354 285640 497360
rect 284944 201544 284996 201550
rect 284944 201486 284996 201492
rect 285600 200002 285628 497354
rect 286336 202366 286364 583510
rect 291844 583228 291896 583234
rect 291844 583170 291896 583176
rect 291108 582820 291160 582826
rect 291108 582762 291160 582768
rect 287704 582480 287756 582486
rect 287704 582422 287756 582428
rect 286876 538280 286928 538286
rect 286876 538222 286928 538228
rect 286416 497004 286468 497010
rect 286416 496946 286468 496952
rect 286428 202434 286456 496946
rect 286416 202428 286468 202434
rect 286416 202370 286468 202376
rect 286324 202360 286376 202366
rect 286324 202302 286376 202308
rect 286232 201544 286284 201550
rect 286232 201486 286284 201492
rect 286244 200002 286272 201486
rect 286888 200002 286916 538222
rect 286968 203788 287020 203794
rect 286968 203730 287020 203736
rect 286980 201550 287008 203730
rect 287520 203720 287572 203726
rect 287520 203662 287572 203668
rect 286968 201544 287020 201550
rect 286968 201486 287020 201492
rect 287532 200002 287560 203662
rect 287716 201618 287744 582422
rect 291016 497752 291068 497758
rect 291016 497694 291068 497700
rect 288348 492720 288400 492726
rect 288348 492662 288400 492668
rect 288360 485926 288388 492662
rect 288348 485920 288400 485926
rect 288348 485862 288400 485868
rect 288256 485716 288308 485722
rect 288256 485658 288308 485664
rect 288268 483002 288296 485658
rect 288256 482996 288308 483002
rect 288256 482938 288308 482944
rect 288256 476060 288308 476066
rect 288256 476002 288308 476008
rect 288268 473362 288296 476002
rect 288268 473334 288388 473362
rect 288360 466546 288388 473334
rect 288348 466540 288400 466546
rect 288348 466482 288400 466488
rect 288256 463820 288308 463826
rect 288256 463762 288308 463768
rect 288268 463690 288296 463762
rect 288256 463684 288308 463690
rect 288256 463626 288308 463632
rect 288256 456748 288308 456754
rect 288256 456690 288308 456696
rect 288268 454050 288296 456690
rect 288268 454022 288388 454050
rect 288360 447234 288388 454022
rect 288348 447228 288400 447234
rect 288348 447170 288400 447176
rect 288348 444440 288400 444446
rect 288268 444388 288348 444394
rect 288268 444382 288400 444388
rect 288268 444378 288388 444382
rect 288256 444372 288388 444378
rect 288308 444366 288388 444372
rect 288256 444314 288308 444320
rect 288268 444283 288296 444314
rect 288256 437436 288308 437442
rect 288256 437378 288308 437384
rect 288268 434738 288296 437378
rect 288268 434710 288388 434738
rect 288360 427922 288388 434710
rect 288348 427916 288400 427922
rect 288348 427858 288400 427864
rect 288348 425128 288400 425134
rect 288268 425076 288348 425082
rect 288268 425070 288400 425076
rect 288268 425066 288388 425070
rect 288072 425060 288124 425066
rect 288072 425002 288124 425008
rect 288256 425060 288388 425066
rect 288308 425054 288388 425060
rect 288256 425002 288308 425008
rect 288084 415426 288112 425002
rect 288268 424971 288296 425002
rect 287992 415398 288112 415426
rect 287992 408406 288020 415398
rect 287980 408400 288032 408406
rect 287980 408342 288032 408348
rect 288348 408400 288400 408406
rect 288348 408342 288400 408348
rect 288360 392193 288388 408342
rect 288346 392184 288402 392193
rect 288346 392119 288402 392128
rect 288162 392048 288218 392057
rect 288162 391983 288218 391992
rect 288176 391950 288204 391983
rect 288164 391944 288216 391950
rect 288164 391886 288216 391892
rect 288348 391944 288400 391950
rect 288348 391886 288400 391892
rect 288360 382265 288388 391886
rect 288346 382256 288402 382265
rect 288346 382191 288402 382200
rect 288530 382256 288586 382265
rect 288530 382191 288586 382200
rect 288544 372638 288572 382191
rect 288348 372632 288400 372638
rect 288348 372574 288400 372580
rect 288532 372632 288584 372638
rect 288532 372574 288584 372580
rect 288360 369918 288388 372574
rect 288348 369912 288400 369918
rect 288348 369854 288400 369860
rect 288348 362976 288400 362982
rect 288348 362918 288400 362924
rect 288360 360262 288388 362918
rect 288348 360256 288400 360262
rect 288348 360198 288400 360204
rect 288348 353320 288400 353326
rect 288348 353262 288400 353268
rect 288360 344622 288388 353262
rect 288348 344616 288400 344622
rect 288348 344558 288400 344564
rect 288348 338156 288400 338162
rect 288348 338098 288400 338104
rect 288360 332042 288388 338098
rect 288348 332036 288400 332042
rect 288348 331978 288400 331984
rect 288164 328500 288216 328506
rect 288164 328442 288216 328448
rect 288176 328370 288204 328442
rect 288164 328364 288216 328370
rect 288164 328306 288216 328312
rect 288348 318844 288400 318850
rect 288348 318786 288400 318792
rect 288360 313410 288388 318786
rect 288348 313404 288400 313410
rect 288348 313346 288400 313352
rect 288348 309188 288400 309194
rect 288348 309130 288400 309136
rect 288360 302258 288388 309130
rect 288348 302252 288400 302258
rect 288348 302194 288400 302200
rect 288348 299532 288400 299538
rect 288348 299474 288400 299480
rect 288360 294098 288388 299474
rect 288348 294092 288400 294098
rect 288348 294034 288400 294040
rect 288164 289876 288216 289882
rect 288164 289818 288216 289824
rect 288176 289746 288204 289818
rect 288164 289740 288216 289746
rect 288164 289682 288216 289688
rect 288348 280220 288400 280226
rect 288348 280162 288400 280168
rect 288360 274786 288388 280162
rect 288348 274780 288400 274786
rect 288348 274722 288400 274728
rect 288164 270564 288216 270570
rect 288164 270506 288216 270512
rect 288176 270434 288204 270506
rect 288164 270428 288216 270434
rect 288164 270370 288216 270376
rect 288348 260908 288400 260914
rect 288348 260850 288400 260856
rect 288360 256034 288388 260850
rect 288176 256006 288388 256034
rect 288176 251274 288204 256006
rect 288176 251246 288296 251274
rect 288268 251190 288296 251246
rect 288256 251184 288308 251190
rect 288256 251126 288308 251132
rect 288348 241528 288400 241534
rect 288348 241470 288400 241476
rect 288360 236026 288388 241470
rect 288348 236020 288400 236026
rect 288348 235962 288400 235968
rect 288164 231872 288216 231878
rect 288254 231840 288310 231849
rect 288216 231820 288254 231826
rect 288164 231814 288254 231820
rect 288176 231798 288254 231814
rect 288254 231775 288310 231784
rect 288530 231840 288586 231849
rect 288530 231775 288586 231784
rect 288544 222222 288572 231775
rect 288348 222216 288400 222222
rect 288348 222158 288400 222164
rect 288532 222216 288584 222222
rect 288532 222158 288584 222164
rect 288360 215370 288388 222158
rect 288176 215342 288388 215370
rect 288176 212566 288204 215342
rect 288072 212560 288124 212566
rect 288072 212502 288124 212508
rect 288164 212560 288216 212566
rect 288164 212502 288216 212508
rect 288084 205714 288112 212502
rect 290924 210452 290976 210458
rect 290924 210394 290976 210400
rect 287992 205686 288112 205714
rect 287704 201612 287756 201618
rect 287704 201554 287756 201560
rect 287992 200002 288020 205686
rect 290556 202836 290608 202842
rect 290556 202778 290608 202784
rect 289268 202768 289320 202774
rect 289268 202710 289320 202716
rect 288808 202632 288860 202638
rect 288808 202574 288860 202580
rect 288820 200002 288848 202574
rect 289280 200002 289308 202710
rect 289544 202088 289596 202094
rect 289544 202030 289596 202036
rect 289556 200002 289584 202030
rect 290568 200002 290596 202778
rect 290936 200138 290964 210394
rect 291028 202842 291056 497694
rect 291120 210458 291148 582762
rect 291108 210452 291160 210458
rect 291108 210394 291160 210400
rect 291016 202836 291068 202842
rect 291016 202778 291068 202784
rect 291384 202836 291436 202842
rect 291384 202778 291436 202784
rect 290936 200110 291056 200138
rect 291028 200002 291056 200110
rect 291396 200002 291424 202778
rect 291856 202774 291884 583170
rect 298928 583160 298980 583166
rect 298928 583102 298980 583108
rect 294604 583092 294656 583098
rect 294604 583034 294656 583040
rect 293868 509312 293920 509318
rect 293868 509254 293920 509260
rect 292304 497344 292356 497350
rect 292304 497286 292356 497292
rect 292212 203924 292264 203930
rect 292212 203866 292264 203872
rect 291844 202768 291896 202774
rect 291844 202710 291896 202716
rect 292224 200138 292252 203866
rect 292316 202842 292344 497286
rect 292488 203856 292540 203862
rect 292488 203798 292540 203804
rect 292304 202836 292356 202842
rect 292304 202778 292356 202784
rect 292224 200110 292344 200138
rect 292316 200002 292344 200110
rect 292500 200002 292528 203798
rect 293132 202836 293184 202842
rect 293132 202778 293184 202784
rect 293144 200002 293172 202778
rect 293880 200002 293908 509254
rect 294420 204264 294472 204270
rect 294420 204206 294472 204212
rect 294432 200002 294460 204206
rect 294616 202842 294644 583034
rect 298652 582888 298704 582894
rect 298652 582830 298704 582836
rect 298468 582548 298520 582554
rect 298468 582490 298520 582496
rect 296718 575784 296774 575793
rect 296718 575719 296774 575728
rect 296732 575550 296760 575719
rect 296720 575544 296772 575550
rect 296720 575486 296772 575492
rect 297454 572928 297510 572937
rect 297454 572863 297510 572872
rect 296442 565856 296498 565865
rect 296442 565791 296498 565800
rect 295984 532908 296036 532914
rect 295984 532850 296036 532856
rect 295996 521626 296024 532850
rect 295340 521620 295392 521626
rect 295340 521562 295392 521568
rect 295984 521620 296036 521626
rect 295984 521562 296036 521568
rect 295352 521286 295380 521562
rect 295340 521280 295392 521286
rect 295340 521222 295392 521228
rect 295352 406774 295380 521222
rect 295340 406768 295392 406774
rect 295340 406710 295392 406716
rect 295352 405890 295380 406710
rect 295340 405884 295392 405890
rect 295340 405826 295392 405832
rect 295984 405884 296036 405890
rect 295984 405826 296036 405832
rect 295996 385762 296024 405826
rect 295984 385756 296036 385762
rect 295984 385698 296036 385704
rect 294880 203992 294932 203998
rect 294880 203934 294932 203940
rect 294604 202836 294656 202842
rect 294604 202778 294656 202784
rect 294892 200002 294920 203934
rect 296168 203448 296220 203454
rect 296168 203390 296220 203396
rect 295800 202836 295852 202842
rect 295800 202778 295852 202784
rect 295812 200002 295840 202778
rect 296180 200002 296208 203390
rect 296456 202842 296484 565791
rect 296902 563408 296958 563417
rect 296902 563343 296958 563352
rect 296916 563106 296944 563343
rect 296904 563100 296956 563106
rect 296904 563042 296956 563048
rect 297086 556880 297142 556889
rect 297086 556815 297142 556824
rect 297100 556238 297128 556815
rect 297088 556232 297140 556238
rect 297088 556174 297140 556180
rect 297362 541104 297418 541113
rect 297362 541039 297418 541048
rect 296534 531448 296590 531457
rect 296534 531383 296590 531392
rect 296444 202836 296496 202842
rect 296444 202778 296496 202784
rect 296548 200002 296576 531383
rect 297086 522200 297142 522209
rect 297086 522135 297142 522144
rect 297100 521694 297128 522135
rect 297088 521688 297140 521694
rect 297088 521630 297140 521636
rect 297376 337550 297404 541039
rect 297468 532914 297496 572863
rect 298006 570072 298062 570081
rect 298006 570007 298062 570016
rect 298020 569974 298048 570007
rect 298008 569968 298060 569974
rect 298008 569910 298060 569916
rect 298006 560416 298062 560425
rect 298006 560351 298062 560360
rect 297914 553616 297970 553625
rect 297914 553551 297970 553560
rect 297822 544096 297878 544105
rect 297822 544031 297878 544040
rect 297730 538384 297786 538393
rect 297730 538319 297786 538328
rect 297744 538286 297772 538319
rect 297732 538280 297784 538286
rect 297732 538222 297784 538228
rect 297456 532908 297508 532914
rect 297456 532850 297508 532856
rect 297454 528864 297510 528873
rect 297454 528799 297510 528808
rect 297468 518226 297496 528799
rect 297730 519208 297786 519217
rect 297730 519143 297786 519152
rect 297744 518974 297772 519143
rect 297732 518968 297784 518974
rect 297732 518910 297784 518916
rect 297456 518220 297508 518226
rect 297456 518162 297508 518168
rect 297730 516216 297786 516225
rect 297730 516151 297732 516160
rect 297784 516151 297786 516160
rect 297732 516122 297784 516128
rect 297730 513496 297786 513505
rect 297730 513431 297786 513440
rect 297638 509688 297694 509697
rect 297638 509623 297694 509632
rect 297652 509318 297680 509623
rect 297640 509312 297692 509318
rect 297640 509254 297692 509260
rect 297638 506696 297694 506705
rect 297638 506631 297694 506640
rect 297652 506530 297680 506631
rect 297640 506524 297692 506530
rect 297640 506466 297692 506472
rect 297364 337544 297416 337550
rect 297364 337486 297416 337492
rect 297744 202502 297772 513431
rect 297732 202496 297784 202502
rect 297732 202438 297784 202444
rect 297836 201958 297864 544031
rect 297928 204202 297956 553551
rect 297916 204196 297968 204202
rect 297916 204138 297968 204144
rect 298020 203250 298048 560351
rect 298480 498846 298508 582490
rect 298560 582412 298612 582418
rect 298560 582354 298612 582360
rect 298468 498840 298520 498846
rect 298468 498782 298520 498788
rect 298572 498302 298600 582354
rect 298664 498982 298692 582830
rect 298744 582752 298796 582758
rect 298744 582694 298796 582700
rect 298652 498976 298704 498982
rect 298652 498918 298704 498924
rect 298560 498296 298612 498302
rect 298560 498238 298612 498244
rect 298008 203244 298060 203250
rect 298008 203186 298060 203192
rect 298756 202842 298784 582694
rect 298836 582616 298888 582622
rect 298836 582558 298888 582564
rect 298848 498914 298876 582558
rect 298940 499118 298968 583102
rect 299020 582956 299072 582962
rect 299020 582898 299072 582904
rect 298928 499112 298980 499118
rect 298928 499054 298980 499060
rect 299032 499050 299060 582898
rect 300492 582684 300544 582690
rect 300492 582626 300544 582632
rect 299388 579692 299440 579698
rect 299388 579634 299440 579640
rect 299294 550760 299350 550769
rect 299294 550695 299350 550704
rect 299202 547904 299258 547913
rect 299202 547839 299258 547848
rect 299110 525872 299166 525881
rect 299110 525807 299166 525816
rect 299020 499044 299072 499050
rect 299020 498986 299072 498992
rect 298836 498908 298888 498914
rect 298836 498850 298888 498856
rect 299020 204060 299072 204066
rect 299020 204002 299072 204008
rect 297916 202836 297968 202842
rect 297916 202778 297968 202784
rect 298744 202836 298796 202842
rect 298744 202778 298796 202784
rect 298928 202836 298980 202842
rect 298928 202778 298980 202784
rect 297824 201952 297876 201958
rect 297824 201894 297876 201900
rect 297548 201884 297600 201890
rect 297548 201826 297600 201832
rect 297560 200002 297588 201826
rect 297928 200002 297956 202778
rect 298376 201748 298428 201754
rect 298376 201690 298428 201696
rect 298388 200002 298416 201690
rect 267752 199974 268088 200002
rect 268212 199974 268548 200002
rect 268672 199974 269008 200002
rect 269132 199974 269376 200002
rect 269500 199974 269836 200002
rect 270296 199974 270448 200002
rect 270664 199974 271000 200002
rect 271124 199974 271460 200002
rect 271584 199974 271828 200002
rect 272044 199974 272288 200002
rect 273332 199974 273668 200002
rect 273792 199974 274036 200002
rect 275080 199974 275324 200002
rect 275448 199974 275784 200002
rect 276828 199974 276980 200002
rect 277196 199974 277348 200002
rect 278576 199974 278728 200002
rect 278944 199974 279280 200002
rect 280232 199974 280568 200002
rect 280692 199974 281028 200002
rect 281980 199974 282316 200002
rect 282440 199974 282684 200002
rect 283360 199974 283604 200002
rect 283728 199974 284064 200002
rect 284188 199974 284248 200002
rect 285476 199974 285628 200002
rect 285936 199974 286272 200002
rect 286764 199974 286916 200002
rect 287224 199974 287560 200002
rect 287684 199974 288020 200002
rect 288512 199974 288848 200002
rect 288972 199974 289308 200002
rect 289432 199974 289584 200002
rect 290260 199974 290596 200002
rect 290720 199974 291056 200002
rect 291180 199974 291424 200002
rect 292008 199974 292344 200002
rect 292468 199974 292528 200002
rect 292928 199974 293172 200002
rect 293756 199974 293908 200002
rect 294216 199974 294460 200002
rect 294584 199974 294920 200002
rect 295504 199974 295840 200002
rect 295964 199974 296208 200002
rect 296332 199974 296576 200002
rect 297252 199974 297588 200002
rect 297712 199974 297956 200002
rect 298080 199974 298416 200002
rect 298940 200002 298968 202778
rect 299032 202042 299060 204002
rect 299124 202774 299152 525807
rect 299112 202768 299164 202774
rect 299112 202710 299164 202716
rect 299216 202706 299244 547839
rect 299204 202700 299256 202706
rect 299204 202642 299256 202648
rect 299032 202014 299152 202042
rect 299124 200002 299152 202014
rect 299308 201618 299336 550695
rect 299400 202570 299428 579634
rect 299480 579352 299532 579358
rect 299480 579294 299532 579300
rect 299388 202564 299440 202570
rect 299388 202506 299440 202512
rect 299492 201686 299520 579294
rect 299570 535460 299626 535469
rect 299570 535395 299626 535404
rect 299584 201822 299612 535395
rect 299662 503908 299718 503917
rect 299662 503843 299718 503852
rect 299676 202638 299704 503843
rect 300504 499186 300532 582626
rect 302804 579972 302832 583646
rect 307024 583636 307076 583642
rect 307024 583578 307076 583584
rect 307036 579972 307064 583578
rect 319720 583568 319772 583574
rect 319720 583510 319772 583516
rect 313464 582480 313516 582486
rect 313464 582422 313516 582428
rect 309232 582412 309284 582418
rect 309232 582354 309284 582360
rect 309244 579972 309272 582354
rect 313476 579972 313504 582422
rect 319732 579972 319760 583510
rect 347504 583500 347556 583506
rect 347504 583442 347556 583448
rect 324136 583432 324188 583438
rect 324136 583374 324188 583380
rect 321928 582548 321980 582554
rect 321928 582490 321980 582496
rect 321940 579972 321968 582490
rect 324148 579972 324176 583374
rect 334624 583364 334676 583370
rect 334624 583306 334676 583312
rect 328368 583228 328420 583234
rect 328368 583170 328420 583176
rect 326160 583024 326212 583030
rect 326160 582966 326212 582972
rect 326172 579972 326200 582966
rect 328380 579972 328408 583170
rect 332600 582616 332652 582622
rect 332600 582558 332652 582564
rect 332612 579972 332640 582558
rect 334636 579972 334664 583306
rect 345296 583296 345348 583302
rect 345296 583238 345348 583244
rect 341064 583160 341116 583166
rect 341064 583102 341116 583108
rect 338856 583092 338908 583098
rect 338856 583034 338908 583040
rect 338868 579972 338896 583034
rect 341076 579972 341104 583102
rect 345308 579972 345336 583238
rect 347516 579972 347544 583442
rect 353760 582956 353812 582962
rect 353760 582898 353812 582904
rect 351736 582820 351788 582826
rect 351736 582762 351788 582768
rect 349526 582448 349582 582457
rect 349526 582383 349582 582392
rect 349540 579972 349568 582383
rect 351748 579972 351776 582762
rect 353772 579972 353800 582898
rect 355968 582888 356020 582894
rect 355968 582830 356020 582836
rect 355980 579972 356008 582830
rect 360200 582752 360252 582758
rect 360200 582694 360252 582700
rect 357992 582616 358044 582622
rect 357992 582558 358044 582564
rect 358004 579972 358032 582558
rect 360212 579972 360240 582694
rect 362408 582684 362460 582690
rect 362408 582626 362460 582632
rect 366640 582684 366692 582690
rect 366640 582626 366692 582632
rect 378876 582684 378928 582690
rect 378876 582626 378928 582632
rect 362420 579972 362448 582626
rect 366652 579972 366680 582626
rect 378416 582616 378468 582622
rect 368662 582584 368718 582593
rect 378416 582558 378468 582564
rect 368662 582519 368718 582528
rect 370872 582548 370924 582554
rect 368676 579972 368704 582519
rect 370872 582490 370924 582496
rect 370884 579972 370912 582490
rect 372896 582412 372948 582418
rect 372896 582354 372948 582360
rect 372908 579972 372936 582354
rect 304828 579698 305026 579714
rect 304816 579692 305026 579698
rect 304868 579686 305026 579692
rect 304816 579634 304868 579640
rect 300676 579352 300728 579358
rect 300610 579300 300676 579306
rect 300610 579294 300728 579300
rect 310980 579352 311032 579358
rect 315212 579352 315264 579358
rect 311032 579300 311282 579306
rect 310980 579294 311282 579300
rect 317420 579352 317472 579358
rect 315264 579300 315514 579306
rect 315212 579294 315514 579300
rect 330208 579352 330260 579358
rect 317472 579300 317722 579306
rect 317420 579294 317722 579300
rect 336648 579352 336700 579358
rect 330260 579300 330418 579306
rect 330208 579294 330418 579300
rect 342996 579352 343048 579358
rect 336700 579300 336858 579306
rect 336648 579294 336858 579300
rect 364248 579352 364300 579358
rect 343048 579300 343298 579306
rect 342996 579294 343298 579300
rect 375380 579352 375432 579358
rect 364300 579300 364458 579306
rect 364248 579294 364458 579300
rect 300610 579278 300716 579294
rect 310992 579278 311282 579294
rect 315224 579278 315514 579294
rect 317432 579278 317722 579294
rect 330220 579278 330418 579294
rect 336660 579278 336858 579294
rect 343008 579278 343298 579294
rect 364260 579278 364458 579294
rect 375130 579300 375380 579306
rect 375130 579294 375432 579300
rect 375130 579278 375420 579294
rect 377154 579278 377260 579306
rect 300610 500126 300716 500154
rect 304842 500126 304948 500154
rect 300492 499180 300544 499186
rect 300492 499122 300544 499128
rect 300688 495394 300716 500126
rect 302424 498296 302476 498302
rect 302424 498238 302476 498244
rect 301504 497072 301556 497078
rect 301504 497014 301556 497020
rect 300596 495366 300716 495394
rect 300596 485858 300624 495366
rect 299940 485852 299992 485858
rect 299940 485794 299992 485800
rect 300584 485852 300636 485858
rect 300584 485794 300636 485800
rect 299952 476134 299980 485794
rect 299756 476128 299808 476134
rect 299940 476128 299992 476134
rect 299808 476076 299888 476082
rect 299756 476070 299888 476076
rect 299940 476070 299992 476076
rect 299768 476054 299888 476070
rect 299860 473346 299888 476054
rect 299848 473340 299900 473346
rect 299848 473282 299900 473288
rect 299848 466404 299900 466410
rect 299848 466346 299900 466352
rect 299860 463706 299888 466346
rect 299860 463678 299980 463706
rect 299952 456822 299980 463678
rect 299756 456816 299808 456822
rect 299940 456816 299992 456822
rect 299808 456764 299888 456770
rect 299756 456758 299888 456764
rect 299940 456758 299992 456764
rect 299768 456742 299888 456758
rect 299860 454034 299888 456742
rect 299848 454028 299900 454034
rect 299848 453970 299900 453976
rect 299848 447092 299900 447098
rect 299848 447034 299900 447040
rect 299860 444394 299888 447034
rect 299860 444366 299980 444394
rect 299952 437510 299980 444366
rect 299756 437504 299808 437510
rect 299940 437504 299992 437510
rect 299808 437452 299888 437458
rect 299756 437446 299888 437452
rect 299940 437446 299992 437452
rect 299768 437430 299888 437446
rect 299860 434722 299888 437430
rect 299848 434716 299900 434722
rect 299848 434658 299900 434664
rect 299848 427780 299900 427786
rect 299848 427722 299900 427728
rect 299860 425082 299888 427722
rect 299860 425054 299980 425082
rect 299952 418198 299980 425054
rect 299756 418192 299808 418198
rect 299940 418192 299992 418198
rect 299808 418140 299888 418146
rect 299756 418134 299888 418140
rect 299940 418134 299992 418140
rect 299768 418118 299888 418134
rect 299860 415410 299888 418118
rect 299848 415404 299900 415410
rect 299848 415346 299900 415352
rect 299940 405748 299992 405754
rect 299940 405690 299992 405696
rect 299952 396098 299980 405690
rect 299848 396092 299900 396098
rect 299848 396034 299900 396040
rect 299940 396092 299992 396098
rect 299940 396034 299992 396040
rect 299860 389178 299888 396034
rect 299860 389150 299980 389178
rect 299952 376786 299980 389150
rect 299848 376780 299900 376786
rect 299848 376722 299900 376728
rect 299940 376780 299992 376786
rect 299940 376722 299992 376728
rect 299860 369866 299888 376722
rect 299860 369838 299980 369866
rect 299952 360210 299980 369838
rect 299768 360182 299980 360210
rect 299768 360074 299796 360182
rect 299768 360046 299888 360074
rect 299860 350538 299888 360046
rect 299848 350532 299900 350538
rect 299848 350474 299900 350480
rect 299940 350464 299992 350470
rect 299940 350406 299992 350412
rect 299952 337618 299980 350406
rect 299940 337612 299992 337618
rect 299940 337554 299992 337560
rect 301412 204128 301464 204134
rect 301412 204070 301464 204076
rect 299664 202632 299716 202638
rect 299664 202574 299716 202580
rect 300124 202360 300176 202366
rect 300124 202302 300176 202308
rect 299572 201816 299624 201822
rect 299572 201758 299624 201764
rect 299480 201680 299532 201686
rect 299480 201622 299532 201628
rect 299296 201612 299348 201618
rect 299296 201554 299348 201560
rect 300136 200002 300164 202302
rect 300768 202020 300820 202026
rect 300768 201962 300820 201968
rect 300780 200002 300808 201962
rect 301424 200002 301452 204070
rect 301516 202842 301544 497014
rect 302148 496868 302200 496874
rect 302148 496810 302200 496816
rect 302160 381546 302188 496810
rect 301596 381540 301648 381546
rect 301596 381482 301648 381488
rect 302148 381540 302200 381546
rect 302148 381482 302200 381488
rect 301608 338094 301636 381482
rect 301596 338088 301648 338094
rect 301596 338030 301648 338036
rect 301504 202836 301556 202842
rect 301504 202778 301556 202784
rect 301872 202428 301924 202434
rect 301872 202370 301924 202376
rect 301884 200002 301912 202370
rect 302436 200002 302464 498238
rect 302620 497622 302648 500004
rect 302608 497616 302660 497622
rect 302608 497558 302660 497564
rect 304540 497616 304592 497622
rect 304540 497558 304592 497564
rect 302620 496874 302648 497558
rect 302608 496868 302660 496874
rect 302608 496810 302660 496816
rect 304552 492697 304580 497558
rect 304170 492688 304226 492697
rect 304170 492623 304226 492632
rect 304538 492688 304594 492697
rect 304538 492623 304594 492632
rect 304184 485858 304212 492623
rect 304172 485852 304224 485858
rect 304172 485794 304224 485800
rect 304264 485716 304316 485722
rect 304264 485658 304316 485664
rect 304276 483002 304304 485658
rect 304264 482996 304316 483002
rect 304264 482938 304316 482944
rect 304448 482996 304500 483002
rect 304448 482938 304500 482944
rect 304460 473385 304488 482938
rect 304262 473376 304318 473385
rect 304446 473376 304502 473385
rect 304262 473311 304264 473320
rect 304316 473311 304318 473320
rect 304356 473340 304408 473346
rect 304264 473282 304316 473288
rect 304446 473311 304502 473320
rect 304356 473282 304408 473288
rect 304368 466290 304396 473282
rect 304276 466262 304396 466290
rect 304276 456890 304304 466262
rect 304264 456884 304316 456890
rect 304264 456826 304316 456832
rect 304264 456748 304316 456754
rect 304264 456690 304316 456696
rect 304276 454034 304304 456690
rect 304264 454028 304316 454034
rect 304264 453970 304316 453976
rect 304356 454028 304408 454034
rect 304356 453970 304408 453976
rect 304368 452606 304396 453970
rect 304356 452600 304408 452606
rect 304356 452542 304408 452548
rect 304172 434784 304224 434790
rect 304172 434726 304224 434732
rect 304184 425082 304212 434726
rect 304184 425054 304304 425082
rect 304276 418266 304304 425054
rect 304264 418260 304316 418266
rect 304264 418202 304316 418208
rect 304172 418124 304224 418130
rect 304172 418066 304224 418072
rect 304184 405770 304212 418066
rect 304184 405742 304304 405770
rect 304276 398954 304304 405742
rect 304264 398948 304316 398954
rect 304264 398890 304316 398896
rect 304264 398812 304316 398818
rect 304264 398754 304316 398760
rect 304276 389230 304304 398754
rect 304264 389224 304316 389230
rect 304264 389166 304316 389172
rect 304172 389156 304224 389162
rect 304172 389098 304224 389104
rect 304184 386458 304212 389098
rect 304184 386430 304304 386458
rect 304276 386374 304304 386430
rect 304264 386368 304316 386374
rect 304264 386310 304316 386316
rect 304264 379364 304316 379370
rect 304264 379306 304316 379312
rect 304276 369918 304304 379306
rect 304264 369912 304316 369918
rect 304264 369854 304316 369860
rect 304172 369844 304224 369850
rect 304172 369786 304224 369792
rect 304184 360262 304212 369786
rect 304172 360256 304224 360262
rect 304172 360198 304224 360204
rect 304264 360188 304316 360194
rect 304264 360130 304316 360136
rect 304276 357270 304304 360130
rect 304264 357264 304316 357270
rect 304264 357206 304316 357212
rect 304264 347880 304316 347886
rect 304264 347822 304316 347828
rect 304276 342938 304304 347822
rect 304184 342910 304304 342938
rect 304184 338099 304212 342910
rect 304170 338090 304226 338099
rect 304170 338025 304226 338034
rect 304446 337920 304502 337929
rect 304446 337855 304502 337864
rect 304460 321450 304488 337855
rect 304276 321422 304488 321450
rect 304276 318782 304304 321422
rect 304264 318776 304316 318782
rect 304264 318718 304316 318724
rect 304264 309256 304316 309262
rect 304264 309198 304316 309204
rect 304276 309126 304304 309198
rect 304264 309120 304316 309126
rect 304264 309062 304316 309068
rect 304264 301708 304316 301714
rect 304264 301650 304316 301656
rect 304276 299470 304304 301650
rect 304264 299464 304316 299470
rect 304264 299406 304316 299412
rect 304264 289944 304316 289950
rect 304264 289886 304316 289892
rect 304276 289814 304304 289886
rect 304264 289808 304316 289814
rect 304264 289750 304316 289756
rect 304264 282804 304316 282810
rect 304264 282746 304316 282752
rect 304276 280158 304304 282746
rect 304264 280152 304316 280158
rect 304264 280094 304316 280100
rect 304264 270632 304316 270638
rect 304264 270574 304316 270580
rect 304276 270502 304304 270574
rect 304264 270496 304316 270502
rect 304264 270438 304316 270444
rect 304448 270496 304500 270502
rect 304448 270438 304500 270444
rect 304460 260953 304488 270438
rect 304078 260944 304134 260953
rect 304078 260879 304134 260888
rect 304446 260944 304502 260953
rect 304446 260879 304502 260888
rect 304092 260846 304120 260879
rect 304080 260840 304132 260846
rect 304080 260782 304132 260788
rect 304264 251252 304316 251258
rect 304264 251194 304316 251200
rect 304276 251138 304304 251194
rect 304184 251110 304304 251138
rect 304184 244322 304212 251110
rect 304172 244316 304224 244322
rect 304172 244258 304224 244264
rect 304172 241528 304224 241534
rect 304172 241470 304224 241476
rect 304184 241398 304212 241470
rect 304172 241392 304224 241398
rect 304172 241334 304224 241340
rect 304172 231872 304224 231878
rect 304262 231840 304318 231849
rect 304224 231820 304262 231826
rect 304172 231814 304262 231820
rect 304184 231798 304262 231814
rect 304262 231775 304318 231784
rect 304538 231840 304594 231849
rect 304538 231775 304594 231784
rect 304552 222222 304580 231775
rect 304356 222216 304408 222222
rect 304356 222158 304408 222164
rect 304540 222216 304592 222222
rect 304540 222158 304592 222164
rect 304368 213450 304396 222158
rect 304172 213444 304224 213450
rect 304172 213386 304224 213392
rect 304356 213444 304408 213450
rect 304356 213386 304408 213392
rect 304184 212514 304212 213386
rect 304092 212486 304212 212514
rect 304092 205698 304120 212486
rect 304080 205692 304132 205698
rect 304080 205634 304132 205640
rect 304264 204196 304316 204202
rect 304264 204138 304316 204144
rect 302884 203312 302936 203318
rect 302884 203254 302936 203260
rect 302896 200002 302924 203254
rect 304080 202904 304132 202910
rect 304080 202846 304132 202852
rect 302976 202700 303028 202706
rect 302976 202642 303028 202648
rect 298940 199974 299000 200002
rect 299124 199974 299368 200002
rect 299828 199974 300164 200002
rect 300748 199974 300808 200002
rect 301116 199974 301452 200002
rect 301576 199974 301912 200002
rect 302404 199974 302464 200002
rect 302864 199974 302924 200002
rect 302988 200002 303016 202642
rect 303896 202496 303948 202502
rect 303896 202438 303948 202444
rect 303908 200002 303936 202438
rect 304092 202434 304120 202846
rect 304080 202428 304132 202434
rect 304080 202370 304132 202376
rect 304276 200002 304304 204138
rect 304920 202502 304948 500126
rect 306472 498840 306524 498846
rect 306472 498782 306524 498788
rect 305644 496936 305696 496942
rect 305644 496878 305696 496884
rect 305656 202842 305684 496878
rect 305644 202836 305696 202842
rect 305644 202778 305696 202784
rect 304908 202496 304960 202502
rect 304908 202438 304960 202444
rect 305644 202020 305696 202026
rect 305644 201962 305696 201968
rect 305000 201544 305052 201550
rect 305000 201486 305052 201492
rect 305012 200002 305040 201486
rect 305656 200002 305684 201962
rect 306484 201754 306512 498782
rect 306852 497010 306880 500004
rect 308968 499990 309074 500018
rect 308968 497010 308996 499990
rect 310612 499112 310664 499118
rect 310612 499054 310664 499060
rect 309140 498908 309192 498914
rect 309140 498850 309192 498856
rect 310428 498908 310480 498914
rect 310428 498850 310480 498856
rect 309048 498840 309100 498846
rect 309048 498782 309100 498788
rect 306840 497004 306892 497010
rect 306840 496946 306892 496952
rect 308956 497004 309008 497010
rect 308956 496946 309008 496952
rect 308404 496868 308456 496874
rect 308404 496810 308456 496816
rect 306656 204196 306708 204202
rect 306656 204138 306708 204144
rect 306472 201748 306524 201754
rect 306472 201690 306524 201696
rect 306668 200002 306696 204138
rect 308416 202434 308444 496810
rect 309060 215234 309088 498782
rect 308876 215206 309088 215234
rect 308876 205714 308904 215206
rect 308784 205686 308904 205714
rect 307024 202428 307076 202434
rect 307024 202370 307076 202376
rect 308404 202428 308456 202434
rect 308404 202370 308456 202376
rect 307036 200002 307064 202370
rect 307300 201748 307352 201754
rect 307300 201690 307352 201696
rect 308404 201748 308456 201754
rect 308404 201690 308456 201696
rect 302988 199974 303324 200002
rect 303908 199974 304152 200002
rect 304276 199974 304612 200002
rect 305012 199974 305072 200002
rect 305656 199974 305900 200002
rect 306360 199974 306696 200002
rect 306820 199974 307064 200002
rect 307312 200002 307340 201690
rect 308416 200002 308444 201690
rect 308784 200002 308812 205686
rect 309152 202842 309180 498850
rect 309140 202836 309192 202842
rect 309140 202778 309192 202784
rect 309600 202836 309652 202842
rect 309600 202778 309652 202784
rect 309140 202496 309192 202502
rect 309140 202438 309192 202444
rect 307312 199974 307648 200002
rect 308108 199974 308444 200002
rect 308568 199974 308812 200002
rect 309152 200002 309180 202438
rect 309612 200002 309640 202778
rect 310440 200002 310468 498850
rect 310624 202502 310652 499054
rect 311084 497214 311112 500004
rect 311900 499180 311952 499186
rect 311900 499122 311952 499128
rect 311072 497208 311124 497214
rect 311072 497150 311124 497156
rect 311912 202842 311940 499122
rect 313292 497962 313320 500004
rect 314844 499044 314896 499050
rect 314844 498986 314896 498992
rect 313280 497956 313332 497962
rect 313280 497898 313332 497904
rect 313556 203516 313608 203522
rect 313556 203458 313608 203464
rect 311900 202836 311952 202842
rect 311900 202778 311952 202784
rect 312544 202836 312596 202842
rect 312544 202778 312596 202784
rect 310612 202496 310664 202502
rect 310612 202438 310664 202444
rect 311256 202496 311308 202502
rect 311256 202438 311308 202444
rect 311164 201952 311216 201958
rect 311164 201894 311216 201900
rect 311176 200002 311204 201894
rect 309152 199974 309396 200002
rect 309612 199974 309856 200002
rect 310316 199974 310468 200002
rect 311144 199974 311204 200002
rect 311268 200002 311296 202438
rect 311992 201816 312044 201822
rect 311992 201758 312044 201764
rect 312004 200002 312032 201758
rect 311268 199974 311604 200002
rect 311972 199974 312032 200002
rect 312556 200002 312584 202778
rect 313568 200002 313596 203458
rect 314856 202842 314884 498986
rect 315316 496874 315344 500004
rect 316040 498976 316092 498982
rect 316040 498918 316092 498924
rect 317328 498976 317380 498982
rect 317328 498918 317380 498924
rect 315948 497208 316000 497214
rect 315948 497150 316000 497156
rect 315304 496868 315356 496874
rect 315304 496810 315356 496816
rect 314844 202836 314896 202842
rect 314844 202778 314896 202784
rect 315580 202836 315632 202842
rect 315580 202778 315632 202784
rect 315304 202088 315356 202094
rect 315304 202030 315356 202036
rect 313648 201884 313700 201890
rect 313648 201826 313700 201832
rect 312556 199974 312892 200002
rect 313352 199974 313596 200002
rect 313660 200002 313688 201826
rect 314936 201612 314988 201618
rect 314936 201554 314988 201560
rect 314948 200002 314976 201554
rect 315316 200002 315344 202030
rect 315396 202020 315448 202026
rect 315396 201962 315448 201968
rect 313660 199974 313720 200002
rect 314640 199974 314976 200002
rect 315100 199974 315344 200002
rect 315408 200002 315436 201962
rect 315592 200002 315620 202778
rect 315960 202094 315988 497150
rect 316052 202094 316080 498918
rect 317340 204762 317368 498918
rect 317524 497282 317552 500004
rect 319732 498137 319760 500004
rect 321468 499044 321520 499050
rect 321468 498986 321520 498992
rect 319718 498128 319774 498137
rect 319718 498063 319774 498072
rect 320088 497956 320140 497962
rect 320088 497898 320140 497904
rect 317512 497276 317564 497282
rect 317512 497218 317564 497224
rect 317064 204734 317368 204762
rect 315948 202088 316000 202094
rect 315948 202030 316000 202036
rect 316040 202088 316092 202094
rect 316040 202030 316092 202036
rect 317064 200002 317092 204734
rect 320100 202774 320128 497898
rect 321480 202774 321508 498986
rect 321756 497146 321784 500004
rect 321744 497140 321796 497146
rect 321744 497082 321796 497088
rect 321744 497004 321796 497010
rect 321744 496946 321796 496952
rect 319260 202768 319312 202774
rect 319260 202710 319312 202716
rect 320088 202768 320140 202774
rect 320088 202710 320140 202716
rect 320548 202768 320600 202774
rect 320548 202710 320600 202716
rect 321468 202768 321520 202774
rect 321468 202710 321520 202716
rect 317144 202088 317196 202094
rect 317144 202030 317196 202036
rect 318616 202088 318668 202094
rect 318616 202030 318668 202036
rect 315408 199974 315468 200002
rect 315592 199974 315928 200002
rect 316756 199974 317092 200002
rect 317156 200002 317184 202030
rect 318628 200002 318656 202030
rect 319272 200002 319300 202710
rect 320560 200002 320588 202710
rect 320640 202020 320692 202026
rect 320640 201962 320692 201968
rect 317156 199974 317216 200002
rect 318504 199974 318656 200002
rect 318964 199974 319300 200002
rect 320252 199974 320588 200002
rect 320652 200002 320680 201962
rect 321756 200002 321784 496946
rect 323964 496942 323992 500004
rect 324228 499112 324280 499118
rect 324228 499054 324280 499060
rect 323952 496936 324004 496942
rect 323952 496878 324004 496884
rect 322940 203380 322992 203386
rect 322940 203322 322992 203328
rect 322952 202434 322980 203322
rect 322940 202428 322992 202434
rect 322940 202370 322992 202376
rect 322756 201884 322808 201890
rect 322756 201826 322808 201832
rect 322768 200002 322796 201826
rect 324044 201544 324096 201550
rect 324044 201486 324096 201492
rect 324056 200002 324084 201486
rect 324240 200002 324268 499054
rect 325988 497078 326016 500004
rect 327092 499990 328210 500018
rect 329852 499990 330234 500018
rect 331232 499990 332442 500018
rect 325976 497072 326028 497078
rect 325976 497014 326028 497020
rect 325148 203244 325200 203250
rect 325148 203186 325200 203192
rect 320652 199974 320712 200002
rect 321756 199974 322000 200002
rect 322460 199974 322796 200002
rect 323748 199974 324084 200002
rect 324208 199974 324268 200002
rect 325160 200002 325188 203186
rect 325700 202700 325752 202706
rect 325700 202642 325752 202648
rect 325712 200002 325740 202642
rect 327092 201550 327120 499990
rect 329852 337482 329880 499990
rect 330484 496868 330536 496874
rect 330484 496810 330536 496816
rect 329840 337476 329892 337482
rect 329840 337418 329892 337424
rect 330496 201958 330524 496810
rect 331232 203318 331260 499990
rect 334452 497894 334480 500004
rect 334440 497888 334492 497894
rect 334440 497830 334492 497836
rect 336660 496874 336688 500004
rect 338868 498030 338896 500004
rect 338856 498024 338908 498030
rect 338856 497966 338908 497972
rect 338764 497888 338816 497894
rect 338764 497830 338816 497836
rect 337384 497276 337436 497282
rect 337384 497218 337436 497224
rect 336648 496868 336700 496874
rect 336648 496810 336700 496816
rect 333888 362976 333940 362982
rect 333888 362918 333940 362924
rect 333796 347064 333848 347070
rect 333796 347006 333848 347012
rect 331220 203312 331272 203318
rect 331220 203254 331272 203260
rect 333152 202768 333204 202774
rect 333152 202710 333204 202716
rect 332508 202428 332560 202434
rect 332508 202370 332560 202376
rect 330484 201952 330536 201958
rect 330484 201894 330536 201900
rect 327080 201544 327132 201550
rect 327080 201486 327132 201492
rect 332520 200002 332548 202370
rect 333164 200002 333192 202710
rect 333808 200274 333836 347006
rect 333900 202774 333928 362918
rect 333888 202768 333940 202774
rect 333888 202710 333940 202716
rect 337396 202094 337424 497218
rect 338776 202638 338804 497830
rect 340144 496868 340196 496874
rect 340144 496810 340196 496816
rect 338764 202632 338816 202638
rect 338764 202574 338816 202580
rect 340156 202162 340184 496810
rect 340892 204270 340920 500004
rect 343100 496874 343128 500004
rect 345124 497418 345152 500004
rect 347332 498098 347360 500004
rect 347320 498092 347372 498098
rect 347320 498034 347372 498040
rect 345112 497412 345164 497418
rect 345112 497354 345164 497360
rect 349356 497214 349384 500004
rect 351564 497350 351592 500004
rect 353312 499990 353602 500018
rect 351552 497344 351604 497350
rect 351552 497286 351604 497292
rect 349344 497208 349396 497214
rect 349344 497150 349396 497156
rect 343088 496868 343140 496874
rect 343088 496810 343140 496816
rect 344928 385824 344980 385830
rect 344928 385766 344980 385772
rect 343548 385212 343600 385218
rect 343548 385154 343600 385160
rect 342168 347336 342220 347342
rect 342168 347278 342220 347284
rect 340880 204264 340932 204270
rect 340880 204206 340932 204212
rect 342076 202768 342128 202774
rect 342076 202710 342128 202716
rect 341432 202632 341484 202638
rect 341432 202574 341484 202580
rect 340144 202156 340196 202162
rect 340144 202098 340196 202104
rect 337384 202088 337436 202094
rect 337384 202030 337436 202036
rect 333716 200246 333836 200274
rect 333716 200138 333744 200246
rect 333624 200110 333744 200138
rect 333624 200002 333652 200110
rect 341444 200002 341472 202574
rect 342088 200002 342116 202710
rect 342180 202638 342208 347278
rect 343560 202638 343588 385154
rect 344008 202700 344060 202706
rect 344008 202642 344060 202648
rect 342168 202632 342220 202638
rect 342168 202574 342220 202580
rect 343088 202632 343140 202638
rect 343088 202574 343140 202580
rect 343548 202632 343600 202638
rect 343548 202574 343600 202580
rect 343100 200002 343128 202574
rect 344020 200002 344048 202642
rect 344940 200002 344968 385766
rect 349068 385552 349120 385558
rect 349068 385494 349120 385500
rect 347688 385280 347740 385286
rect 347688 385222 347740 385228
rect 347596 369912 347648 369918
rect 347596 369854 347648 369860
rect 345756 204264 345808 204270
rect 345756 204206 345808 204212
rect 345768 200002 345796 204206
rect 347608 202638 347636 369854
rect 346676 202632 346728 202638
rect 346676 202574 346728 202580
rect 347596 202632 347648 202638
rect 347596 202574 347648 202580
rect 346688 200002 346716 202574
rect 347700 200138 347728 385222
rect 348332 202156 348384 202162
rect 348332 202098 348384 202104
rect 347516 200110 347728 200138
rect 347516 200002 347544 200110
rect 348344 200002 348372 202098
rect 349080 200002 349108 385494
rect 353208 385348 353260 385354
rect 353208 385290 353260 385296
rect 351828 376780 351880 376786
rect 351828 376722 351880 376728
rect 350448 347404 350500 347410
rect 350448 347346 350500 347352
rect 350460 202774 350488 347346
rect 351840 202774 351868 376722
rect 349988 202768 350040 202774
rect 349988 202710 350040 202716
rect 350448 202768 350500 202774
rect 350448 202710 350500 202716
rect 351000 202768 351052 202774
rect 351000 202710 351052 202716
rect 351828 202768 351880 202774
rect 351828 202710 351880 202716
rect 350000 200002 350028 202710
rect 351012 200002 351040 202710
rect 353220 202094 353248 385290
rect 353312 203454 353340 499990
rect 355796 497282 355824 500004
rect 358004 497962 358032 500004
rect 357992 497956 358044 497962
rect 357992 497898 358044 497904
rect 360028 497554 360056 500004
rect 362236 497894 362264 500004
rect 364260 498166 364288 500004
rect 364248 498160 364300 498166
rect 364248 498102 364300 498108
rect 362224 497888 362276 497894
rect 362224 497830 362276 497836
rect 366468 497622 366496 500004
rect 368492 497826 368520 500004
rect 369872 499990 370714 500018
rect 368480 497820 368532 497826
rect 368480 497762 368532 497768
rect 366456 497616 366508 497622
rect 366456 497558 366508 497564
rect 360016 497548 360068 497554
rect 360016 497490 360068 497496
rect 355784 497276 355836 497282
rect 355784 497218 355836 497224
rect 369124 385620 369176 385626
rect 369124 385562 369176 385568
rect 355876 385484 355928 385490
rect 355876 385426 355928 385432
rect 354588 353320 354640 353326
rect 354588 353262 354640 353268
rect 354496 347200 354548 347206
rect 354496 347142 354548 347148
rect 353300 203448 353352 203454
rect 353300 203390 353352 203396
rect 353576 202156 353628 202162
rect 353576 202098 353628 202104
rect 352748 202088 352800 202094
rect 352748 202030 352800 202036
rect 353208 202088 353260 202094
rect 353208 202030 353260 202036
rect 351736 202020 351788 202026
rect 351736 201962 351788 201968
rect 351748 200002 351776 201962
rect 352760 200002 352788 202030
rect 353588 200002 353616 202098
rect 354508 200002 354536 347142
rect 354600 202162 354628 353262
rect 354588 202156 354640 202162
rect 354588 202098 354640 202104
rect 355324 201544 355376 201550
rect 355324 201486 355376 201492
rect 355336 200002 355364 201486
rect 325160 199974 325496 200002
rect 325712 199974 325956 200002
rect 332488 199974 332548 200002
rect 332856 199974 333192 200002
rect 333316 199974 333652 200002
rect 341136 199974 341472 200002
rect 342056 199974 342116 200002
rect 342884 199974 343128 200002
rect 343712 199974 344048 200002
rect 344632 199974 344968 200002
rect 345460 199974 345796 200002
rect 346380 199974 346716 200002
rect 347208 199974 347544 200002
rect 348128 199974 348372 200002
rect 348956 199974 349108 200002
rect 349876 199974 350028 200002
rect 350704 199974 351040 200002
rect 351624 199974 351776 200002
rect 352452 199974 352788 200002
rect 353280 199974 353616 200002
rect 354200 199974 354536 200002
rect 355028 199974 355364 200002
rect 355888 200002 355916 385426
rect 357348 385416 357400 385422
rect 357348 385358 357400 385364
rect 355968 385144 356020 385150
rect 355968 385086 356020 385092
rect 355980 201550 356008 385086
rect 355968 201544 356020 201550
rect 355968 201486 356020 201492
rect 357360 200138 357388 385358
rect 367008 385076 367060 385082
rect 367008 385018 367060 385024
rect 364248 374060 364300 374066
rect 364248 374002 364300 374008
rect 360108 347676 360160 347682
rect 360108 347618 360160 347624
rect 358728 347540 358780 347546
rect 358728 347482 358780 347488
rect 357900 201952 357952 201958
rect 357900 201894 357952 201900
rect 357084 200110 357388 200138
rect 357084 200002 357112 200110
rect 357912 200002 357940 201894
rect 358740 200002 358768 347482
rect 360120 201550 360148 347618
rect 362868 347608 362920 347614
rect 362868 347550 362920 347556
rect 362776 347472 362828 347478
rect 362776 347414 362828 347420
rect 361488 347268 361540 347274
rect 361488 347210 361540 347216
rect 361396 347132 361448 347138
rect 361396 347074 361448 347080
rect 361408 201550 361436 347074
rect 359648 201544 359700 201550
rect 359648 201486 359700 201492
rect 360108 201544 360160 201550
rect 360108 201486 360160 201492
rect 360568 201544 360620 201550
rect 360568 201486 360620 201492
rect 361396 201544 361448 201550
rect 361396 201486 361448 201492
rect 359660 200002 359688 201486
rect 360580 200002 360608 201486
rect 361500 200138 361528 347210
rect 362788 201550 362816 347414
rect 362316 201544 362368 201550
rect 362316 201486 362368 201492
rect 362776 201544 362828 201550
rect 362776 201486 362828 201492
rect 361408 200110 361528 200138
rect 361408 200002 361436 200110
rect 362328 200002 362356 201486
rect 362880 200002 362908 347550
rect 364260 200138 364288 374002
rect 367020 202162 367048 385018
rect 366180 202156 366232 202162
rect 366180 202098 366232 202104
rect 367008 202156 367060 202162
rect 367008 202098 367060 202104
rect 365352 202020 365404 202026
rect 365352 201962 365404 201968
rect 364892 201748 364944 201754
rect 364892 201690 364944 201696
rect 364076 200110 364288 200138
rect 364076 200002 364104 200110
rect 364904 200002 364932 201690
rect 365364 200002 365392 201962
rect 366192 200002 366220 202098
rect 369136 202026 369164 385562
rect 369872 203658 369900 499990
rect 372724 497486 372752 500004
rect 374932 497690 374960 500004
rect 377140 497758 377168 500004
rect 377128 497752 377180 497758
rect 377128 497694 377180 497700
rect 374920 497684 374972 497690
rect 374920 497626 374972 497632
rect 372712 497480 372764 497486
rect 372712 497422 372764 497428
rect 375288 387116 375340 387122
rect 375288 387058 375340 387064
rect 369860 203652 369912 203658
rect 369860 203594 369912 203600
rect 375300 202366 375328 387058
rect 375748 202836 375800 202842
rect 375748 202778 375800 202784
rect 374460 202360 374512 202366
rect 374460 202302 374512 202308
rect 375288 202360 375340 202366
rect 375288 202302 375340 202308
rect 369124 202020 369176 202026
rect 369124 201962 369176 201968
rect 366916 201816 366968 201822
rect 366916 201758 366968 201764
rect 366928 200002 366956 201758
rect 374472 200002 374500 202302
rect 375760 200002 375788 202778
rect 377232 202570 377260 579278
rect 377310 565856 377366 565865
rect 377310 565791 377366 565800
rect 377324 203794 377352 565791
rect 377402 563136 377458 563145
rect 377402 563071 377458 563080
rect 377416 203998 377444 563071
rect 378138 560212 378194 560221
rect 378138 560147 378194 560156
rect 377494 556608 377550 556617
rect 377494 556543 377550 556552
rect 377404 203992 377456 203998
rect 377404 203934 377456 203940
rect 377312 203788 377364 203794
rect 377312 203730 377364 203736
rect 377220 202564 377272 202570
rect 377220 202506 377272 202512
rect 377508 202502 377536 556543
rect 377496 202496 377548 202502
rect 377496 202438 377548 202444
rect 378152 202298 378180 560147
rect 378230 550692 378286 550701
rect 378230 550627 378286 550636
rect 378140 202292 378192 202298
rect 378140 202234 378192 202240
rect 376484 202156 376536 202162
rect 376484 202098 376536 202104
rect 376496 200002 376524 202098
rect 378244 201890 378272 550627
rect 378322 547700 378378 547709
rect 378322 547635 378378 547644
rect 378336 202230 378364 547635
rect 378428 499118 378456 582558
rect 378692 582548 378744 582554
rect 378692 582490 378744 582496
rect 378600 582412 378652 582418
rect 378600 582354 378652 582360
rect 378508 579352 378560 579358
rect 378508 579294 378560 579300
rect 378416 499112 378468 499118
rect 378416 499054 378468 499060
rect 378520 499050 378548 579294
rect 378508 499044 378560 499050
rect 378508 498986 378560 498992
rect 378612 498846 378640 582354
rect 378704 498914 378732 582490
rect 378784 556232 378836 556238
rect 378784 556174 378836 556180
rect 378692 498908 378744 498914
rect 378692 498850 378744 498856
rect 378600 498840 378652 498846
rect 378600 498782 378652 498788
rect 378796 202842 378824 556174
rect 378888 498982 378916 582626
rect 380622 575512 380678 575521
rect 380622 575447 380678 575456
rect 379518 569120 379574 569129
rect 379518 569055 379574 569064
rect 378966 515536 379022 515545
rect 378966 515471 379022 515480
rect 378876 498976 378928 498982
rect 378876 498918 378928 498924
rect 378784 202836 378836 202842
rect 378784 202778 378836 202784
rect 378980 202366 379008 515471
rect 379532 203522 379560 569055
rect 379610 553480 379666 553489
rect 379610 553415 379666 553424
rect 379624 204134 379652 553415
rect 379702 543824 379758 543833
rect 379702 543759 379758 543768
rect 379612 204128 379664 204134
rect 379612 204070 379664 204076
rect 379716 203726 379744 543759
rect 379794 537568 379850 537577
rect 379794 537503 379850 537512
rect 379808 203930 379836 537503
rect 379886 534576 379942 534585
rect 379886 534511 379942 534520
rect 379796 203924 379848 203930
rect 379796 203866 379848 203872
rect 379900 203862 379928 534511
rect 379978 531448 380034 531457
rect 379978 531383 380034 531392
rect 379888 203856 379940 203862
rect 379888 203798 379940 203804
rect 379704 203720 379756 203726
rect 379704 203662 379756 203668
rect 379992 203590 380020 531383
rect 380530 528728 380586 528737
rect 380530 528663 380586 528672
rect 380070 525056 380126 525065
rect 380070 524991 380126 525000
rect 379980 203584 380032 203590
rect 379980 203526 380032 203532
rect 379520 203516 379572 203522
rect 379520 203458 379572 203464
rect 378968 202360 379020 202366
rect 378968 202302 379020 202308
rect 378324 202224 378376 202230
rect 378324 202166 378376 202172
rect 378232 201884 378284 201890
rect 378232 201826 378284 201832
rect 380084 201686 380112 524991
rect 380162 521792 380218 521801
rect 380162 521727 380218 521736
rect 380176 203386 380204 521727
rect 380254 512544 380310 512553
rect 380254 512479 380310 512488
rect 380164 203380 380216 203386
rect 380164 203322 380216 203328
rect 380072 201680 380124 201686
rect 380072 201622 380124 201628
rect 380268 201618 380296 512479
rect 380346 509416 380402 509425
rect 380346 509351 380402 509360
rect 380360 204066 380388 509351
rect 380438 506560 380494 506569
rect 380438 506495 380494 506504
rect 380452 500954 380480 506495
rect 380440 500948 380492 500954
rect 380440 500890 380492 500896
rect 380440 500812 380492 500818
rect 380440 500754 380492 500760
rect 380452 204202 380480 500754
rect 380544 337414 380572 528663
rect 380636 407930 380664 575447
rect 420184 556300 420236 556306
rect 420184 556242 420236 556248
rect 380714 519208 380770 519217
rect 380714 519143 380770 519152
rect 380728 503130 380756 519143
rect 380716 503124 380768 503130
rect 380716 503066 380768 503072
rect 380714 503024 380770 503033
rect 380714 502959 380770 502968
rect 380728 500818 380756 502959
rect 380716 500812 380768 500818
rect 380716 500754 380768 500760
rect 380624 407924 380676 407930
rect 380624 407866 380676 407872
rect 416964 407856 417016 407862
rect 416964 407798 417016 407804
rect 402980 407788 403032 407794
rect 402980 407730 403032 407736
rect 402992 393310 403020 407730
rect 411260 407244 411312 407250
rect 411260 407186 411312 407192
rect 402980 393304 403032 393310
rect 402980 393246 403032 393252
rect 403900 393304 403952 393310
rect 403900 393246 403952 393252
rect 388260 385756 388312 385762
rect 388260 385698 388312 385704
rect 385868 385552 385920 385558
rect 385868 385494 385920 385500
rect 385880 383316 385908 385494
rect 388272 383316 388300 385698
rect 392860 385620 392912 385626
rect 392860 385562 392912 385568
rect 390468 385076 390520 385082
rect 390468 385018 390520 385024
rect 390480 383316 390508 385018
rect 392872 383316 392900 385562
rect 399668 385484 399720 385490
rect 399668 385426 399720 385432
rect 397460 385280 397512 385286
rect 397460 385222 397512 385228
rect 395068 385212 395120 385218
rect 395068 385154 395120 385160
rect 395080 383316 395108 385154
rect 397472 383316 397500 385222
rect 399680 383316 399708 385426
rect 402060 385348 402112 385354
rect 402060 385290 402112 385296
rect 402072 383316 402100 385290
rect 403912 383330 403940 393246
rect 408868 385824 408920 385830
rect 408868 385766 408920 385772
rect 406660 385416 406712 385422
rect 406660 385358 406712 385364
rect 403912 383302 404294 383330
rect 406672 383316 406700 385358
rect 408880 383316 408908 385766
rect 411272 383316 411300 407186
rect 416872 407176 416924 407182
rect 416872 407118 416924 407124
rect 416596 389428 416648 389434
rect 416596 389370 416648 389376
rect 414664 389360 414716 389366
rect 414664 389302 414716 389308
rect 413468 385144 413520 385150
rect 413468 385086 413520 385092
rect 413480 383316 413508 385086
rect 380900 381540 380952 381546
rect 380900 381482 380952 381488
rect 380912 381449 380940 381482
rect 380898 381440 380954 381449
rect 380898 381375 380954 381384
rect 380898 377224 380954 377233
rect 380898 377159 380954 377168
rect 380912 376786 380940 377159
rect 380900 376780 380952 376786
rect 380900 376722 380952 376728
rect 380898 374096 380954 374105
rect 380898 374031 380900 374040
rect 380952 374031 380954 374040
rect 380900 374002 380952 374008
rect 380898 370424 380954 370433
rect 380898 370359 380954 370368
rect 380912 369918 380940 370359
rect 380900 369912 380952 369918
rect 380900 369854 380952 369860
rect 381634 367432 381690 367441
rect 381634 367367 381690 367376
rect 380898 363624 380954 363633
rect 380898 363559 380954 363568
rect 380912 362982 380940 363559
rect 380900 362976 380952 362982
rect 380900 362918 380952 362924
rect 380898 353560 380954 353569
rect 380898 353495 380954 353504
rect 380912 353326 380940 353495
rect 380900 353320 380952 353326
rect 380900 353262 380952 353268
rect 381544 347744 381596 347750
rect 381544 347686 381596 347692
rect 380532 337408 380584 337414
rect 380532 337350 380584 337356
rect 380440 204196 380492 204202
rect 380440 204138 380492 204144
rect 380348 204060 380400 204066
rect 380348 204002 380400 204008
rect 381556 201754 381584 347686
rect 381648 340678 381676 367367
rect 381726 360360 381782 360369
rect 381726 360295 381782 360304
rect 381740 340746 381768 360295
rect 381818 356824 381874 356833
rect 381818 356759 381874 356768
rect 381728 340740 381780 340746
rect 381728 340682 381780 340688
rect 381636 340672 381688 340678
rect 381636 340614 381688 340620
rect 381832 340542 381860 356759
rect 383672 350118 384606 350146
rect 383672 340610 383700 350118
rect 386800 347750 386828 350132
rect 386788 347744 386840 347750
rect 386788 347686 386840 347692
rect 389008 347342 389036 350132
rect 391400 347682 391428 350132
rect 391388 347676 391440 347682
rect 391388 347618 391440 347624
rect 393608 347546 393636 350132
rect 393596 347540 393648 347546
rect 393596 347482 393648 347488
rect 396000 347410 396028 350132
rect 398208 347614 398236 350132
rect 398196 347608 398248 347614
rect 398196 347550 398248 347556
rect 395988 347404 396040 347410
rect 395988 347346 396040 347352
rect 388996 347336 389048 347342
rect 388996 347278 389048 347284
rect 400600 347206 400628 350132
rect 402808 347478 402836 350132
rect 404372 350118 405214 350146
rect 402796 347472 402848 347478
rect 402796 347414 402848 347420
rect 400588 347200 400640 347206
rect 400588 347142 400640 347148
rect 404372 340814 404400 350118
rect 407408 347274 407436 350132
rect 408512 350118 409814 350146
rect 407396 347268 407448 347274
rect 407396 347210 407448 347216
rect 408512 340882 408540 350118
rect 412008 347070 412036 350132
rect 414400 347138 414428 350132
rect 414388 347132 414440 347138
rect 414388 347074 414440 347080
rect 411996 347064 412048 347070
rect 411996 347006 412048 347012
rect 408500 340876 408552 340882
rect 408500 340818 408552 340824
rect 404360 340808 404412 340814
rect 404360 340750 404412 340756
rect 383660 340604 383712 340610
rect 383660 340546 383712 340552
rect 381820 340536 381872 340542
rect 381820 340478 381872 340484
rect 401508 337612 401560 337618
rect 401508 337554 401560 337560
rect 401520 202842 401548 337554
rect 411168 337544 411220 337550
rect 411168 337486 411220 337492
rect 408408 337476 408460 337482
rect 408408 337418 408460 337424
rect 400588 202836 400640 202842
rect 400588 202778 400640 202784
rect 401508 202836 401560 202842
rect 401508 202778 401560 202784
rect 381544 201748 381596 201754
rect 381544 201690 381596 201696
rect 380256 201612 380308 201618
rect 380256 201554 380308 201560
rect 400600 200002 400628 202778
rect 400956 202564 401008 202570
rect 400956 202506 401008 202512
rect 400968 200002 400996 202506
rect 408420 200002 408448 337418
rect 411076 202224 411128 202230
rect 411076 202166 411128 202172
rect 410156 201748 410208 201754
rect 410156 201690 410208 201696
rect 409236 201680 409288 201686
rect 409236 201622 409288 201628
rect 409248 200002 409276 201622
rect 410168 200002 410196 201690
rect 355888 199974 355948 200002
rect 356776 199974 357112 200002
rect 357696 199974 357940 200002
rect 358524 199974 358768 200002
rect 359444 199974 359688 200002
rect 360272 199974 360608 200002
rect 361192 199974 361436 200002
rect 362020 199974 362356 200002
rect 362848 199974 362908 200002
rect 363768 199974 364104 200002
rect 364596 199974 364932 200002
rect 365056 199974 365392 200002
rect 365976 199974 366220 200002
rect 366804 199974 366956 200002
rect 374164 199974 374500 200002
rect 375452 199974 375788 200002
rect 376372 199974 376524 200002
rect 400292 199974 400628 200002
rect 400752 199974 400996 200002
rect 408112 199974 408448 200002
rect 408940 199974 409276 200002
rect 409860 199974 410196 200002
rect 411088 200002 411116 202166
rect 411180 201754 411208 337486
rect 413928 337408 413980 337414
rect 413928 337350 413980 337356
rect 413192 202496 413244 202502
rect 413192 202438 413244 202444
rect 412272 201884 412324 201890
rect 412272 201826 412324 201832
rect 411168 201748 411220 201754
rect 411168 201690 411220 201696
rect 412284 200002 412312 201826
rect 413204 200002 413232 202438
rect 413940 200002 413968 337350
rect 414676 202570 414704 389302
rect 416044 374060 416096 374066
rect 416044 374002 416096 374008
rect 415398 363964 415454 363973
rect 415398 363899 415454 363908
rect 415412 202638 415440 363899
rect 415400 202632 415452 202638
rect 415400 202574 415452 202580
rect 414664 202564 414716 202570
rect 414664 202506 414716 202512
rect 416056 202502 416084 374002
rect 416412 212560 416464 212566
rect 416412 212502 416464 212508
rect 416044 202496 416096 202502
rect 416044 202438 416096 202444
rect 415768 202428 415820 202434
rect 415768 202370 415820 202376
rect 414940 202292 414992 202298
rect 414940 202234 414992 202240
rect 414952 200002 414980 202234
rect 415780 200002 415808 202370
rect 416424 200002 416452 212502
rect 416608 202434 416636 389370
rect 416688 389224 416740 389230
rect 416688 389166 416740 389172
rect 416700 212566 416728 389166
rect 416884 380905 416912 407118
rect 416870 380896 416926 380905
rect 416870 380831 416926 380840
rect 416778 376952 416834 376961
rect 416778 376887 416834 376896
rect 416688 212560 416740 212566
rect 416688 212502 416740 212508
rect 416596 202428 416648 202434
rect 416596 202370 416648 202376
rect 416792 202366 416820 376887
rect 416976 374649 417004 407798
rect 418068 389292 418120 389298
rect 418068 389234 418120 389240
rect 416962 374640 417018 374649
rect 416962 374575 417018 374584
rect 416870 370152 416926 370161
rect 416870 370087 416926 370096
rect 416884 202706 416912 370087
rect 416962 367160 417018 367169
rect 416962 367095 417018 367104
rect 416872 202700 416924 202706
rect 416872 202642 416924 202648
rect 416780 202360 416832 202366
rect 416780 202302 416832 202308
rect 416976 201958 417004 367095
rect 417054 360224 417110 360233
rect 417054 360159 417110 360168
rect 417068 204270 417096 360159
rect 417146 356552 417202 356561
rect 417146 356487 417202 356496
rect 417056 204264 417108 204270
rect 417056 204206 417108 204212
rect 417160 202774 417188 356487
rect 417238 353424 417294 353433
rect 417238 353359 417294 353368
rect 417148 202768 417200 202774
rect 417148 202710 417200 202716
rect 417252 202094 417280 353359
rect 418080 202434 418108 389234
rect 417516 202428 417568 202434
rect 417516 202370 417568 202376
rect 418068 202428 418120 202434
rect 418068 202370 418120 202376
rect 417240 202088 417292 202094
rect 417240 202030 417292 202036
rect 416964 201952 417016 201958
rect 416964 201894 417016 201900
rect 417528 200002 417556 202370
rect 420196 201822 420224 556242
rect 420184 201816 420236 201822
rect 420184 201758 420236 201764
rect 411088 199974 411148 200002
rect 411976 199974 412312 200002
rect 412896 199974 413232 200002
rect 413724 199974 413968 200002
rect 414644 199974 414980 200002
rect 415472 199974 415808 200002
rect 416392 199974 416452 200002
rect 417220 199974 417556 200002
rect 243872 199860 244168 199866
rect 243820 199854 244168 199860
rect 239508 199838 239844 199854
rect 243832 199838 244168 199854
rect 266340 199838 266676 199866
rect 433904 157321 433932 699654
rect 433996 159361 434024 700674
rect 434088 161265 434116 700878
rect 434168 700800 434220 700806
rect 434168 700742 434220 700748
rect 434180 163577 434208 700742
rect 434352 700664 434404 700670
rect 434352 700606 434404 700612
rect 434260 700324 434312 700330
rect 434260 700266 434312 700272
rect 434272 169697 434300 700266
rect 434258 169688 434314 169697
rect 434258 169623 434314 169632
rect 434364 165617 434392 700606
rect 434444 700460 434496 700466
rect 434444 700402 434496 700408
rect 438124 700460 438176 700466
rect 438124 700402 438176 700408
rect 434456 167793 434484 700402
rect 434720 681760 434772 681766
rect 434720 681702 434772 681708
rect 434536 294024 434588 294030
rect 434536 293966 434588 293972
rect 434548 186289 434576 293966
rect 434534 186280 434590 186289
rect 434534 186215 434590 186224
rect 434732 172009 434760 681702
rect 434812 623824 434864 623830
rect 434812 623766 434864 623772
rect 434824 173913 434852 623766
rect 436744 438932 436796 438938
rect 436744 438874 436796 438880
rect 436100 385688 436152 385694
rect 436100 385630 436152 385636
rect 434904 336796 434956 336802
rect 434904 336738 434956 336744
rect 434916 184657 434944 336738
rect 435088 251252 435140 251258
rect 435088 251194 435140 251200
rect 434994 196208 435050 196217
rect 434994 196143 435050 196152
rect 434902 184648 434958 184657
rect 434902 184583 434958 184592
rect 434810 173904 434866 173913
rect 434810 173839 434866 173848
rect 434718 172000 434774 172009
rect 434718 171935 434774 171944
rect 434442 167784 434498 167793
rect 434442 167719 434498 167728
rect 434350 165608 434406 165617
rect 434350 165543 434406 165552
rect 434166 163568 434222 163577
rect 434166 163503 434222 163512
rect 434074 161256 434130 161265
rect 434074 161191 434130 161200
rect 433982 159352 434038 159361
rect 433982 159287 434038 159296
rect 433890 157312 433946 157321
rect 433890 157247 433946 157256
rect 134064 122392 134116 122398
rect 134064 122334 134116 122340
rect 134062 121952 134118 121961
rect 134062 121887 134118 121896
rect 134076 120834 134104 121887
rect 134064 120828 134116 120834
rect 134064 120770 134116 120776
rect 133972 120692 134024 120698
rect 133972 120634 134024 120640
rect 135168 120352 135220 120358
rect 135168 120294 135220 120300
rect 133892 120006 134320 120034
rect 134536 120006 134872 120034
rect 133786 117872 133842 117881
rect 133786 117807 133842 117816
rect 133800 117298 133828 117807
rect 133788 117292 133840 117298
rect 133788 117234 133840 117240
rect 133788 115932 133840 115938
rect 133788 115874 133840 115880
rect 133800 106321 133828 115874
rect 133786 106312 133842 106321
rect 133786 106247 133842 106256
rect 133604 41404 133656 41410
rect 133604 41346 133656 41352
rect 133512 37324 133564 37330
rect 133512 37266 133564 37272
rect 132408 30320 132460 30326
rect 132408 30262 132460 30268
rect 133524 29034 133552 37266
rect 133328 29028 133380 29034
rect 133328 28970 133380 28976
rect 133512 29028 133564 29034
rect 133512 28970 133564 28976
rect 133340 27606 133368 28970
rect 133328 27600 133380 27606
rect 133328 27542 133380 27548
rect 132224 22092 132276 22098
rect 132224 22034 132276 22040
rect 133328 19304 133380 19310
rect 133328 19246 133380 19252
rect 133340 9722 133368 19246
rect 133144 9716 133196 9722
rect 133144 9658 133196 9664
rect 133328 9716 133380 9722
rect 133328 9658 133380 9664
rect 133156 8634 133184 9658
rect 133144 8628 133196 8634
rect 133144 8570 133196 8576
rect 131764 8288 131816 8294
rect 131764 8230 131816 8236
rect 133788 8288 133840 8294
rect 133788 8230 133840 8236
rect 131396 7200 131448 7206
rect 131396 7142 131448 7148
rect 130384 4480 130436 4486
rect 130384 4422 130436 4428
rect 131408 480 131436 7142
rect 132592 7064 132644 7070
rect 132592 7006 132644 7012
rect 132604 480 132632 7006
rect 133800 480 133828 8230
rect 133892 7614 133920 120006
rect 133970 117736 134026 117745
rect 134154 117736 134210 117745
rect 134026 117694 134154 117722
rect 133970 117671 134026 117680
rect 134154 117671 134210 117680
rect 134536 115938 134564 120006
rect 135180 119406 135208 120294
rect 186608 120290 186944 120306
rect 186596 120284 186944 120290
rect 186648 120278 186944 120284
rect 393852 120278 394188 120306
rect 425684 120278 426112 120306
rect 186596 120226 186648 120232
rect 145024 120154 145268 120170
rect 145012 120148 145268 120154
rect 145064 120142 145268 120148
rect 159468 120142 159988 120170
rect 164988 120142 165508 120170
rect 145012 120090 145064 120096
rect 135364 120006 135516 120034
rect 135732 120006 136068 120034
rect 136712 120006 136864 120034
rect 135168 119400 135220 119406
rect 135168 119342 135220 119348
rect 135260 117700 135312 117706
rect 135260 117642 135312 117648
rect 135272 117570 135300 117642
rect 135260 117564 135312 117570
rect 135260 117506 135312 117512
rect 134524 115932 134576 115938
rect 134524 115874 134576 115880
rect 135260 113892 135312 113898
rect 135260 113834 135312 113840
rect 133970 106312 134026 106321
rect 133970 106247 133972 106256
rect 134024 106247 134026 106256
rect 133972 106218 134024 106224
rect 133972 106140 134024 106146
rect 133972 106082 134024 106088
rect 133984 91746 134012 106082
rect 133984 91718 134104 91746
rect 134076 60738 134104 91718
rect 133984 60710 134104 60738
rect 133984 60602 134012 60710
rect 133984 60574 134104 60602
rect 134076 41426 134104 60574
rect 133984 41398 134104 41426
rect 133984 41290 134012 41398
rect 133984 41262 134104 41290
rect 134076 22114 134104 41262
rect 133984 22086 134104 22114
rect 133984 21978 134012 22086
rect 133984 21950 134104 21978
rect 134076 7750 134104 21950
rect 135272 7818 135300 113834
rect 135260 7812 135312 7818
rect 135260 7754 135312 7760
rect 134064 7744 134116 7750
rect 134064 7686 134116 7692
rect 135364 7682 135392 120006
rect 135444 117564 135496 117570
rect 135444 117506 135496 117512
rect 135456 9178 135484 117506
rect 135732 113898 135760 120006
rect 135720 113892 135772 113898
rect 135720 113834 135772 113840
rect 136732 112532 136784 112538
rect 136732 112474 136784 112480
rect 135444 9172 135496 9178
rect 135444 9114 135496 9120
rect 136744 7886 136772 112474
rect 136836 8974 136864 120006
rect 136928 120006 137356 120034
rect 137572 120006 137908 120034
rect 136824 8968 136876 8974
rect 136824 8910 136876 8916
rect 136732 7880 136784 7886
rect 136732 7822 136784 7828
rect 136088 7744 136140 7750
rect 136088 7686 136140 7692
rect 135352 7676 135404 7682
rect 135352 7618 135404 7624
rect 133880 7608 133932 7614
rect 133880 7550 133932 7556
rect 134892 7608 134944 7614
rect 134892 7550 134944 7556
rect 134904 480 134932 7550
rect 136100 480 136128 7686
rect 136928 3466 136956 120006
rect 137572 112538 137600 120006
rect 138538 119785 138566 120020
rect 138860 120006 139196 120034
rect 139504 120006 139748 120034
rect 140056 120006 140392 120034
rect 140792 120006 141036 120034
rect 141252 120006 141588 120034
rect 142232 120006 142384 120034
rect 138524 119776 138580 119785
rect 138524 119711 138580 119720
rect 138860 119338 138888 120006
rect 138296 119332 138348 119338
rect 138296 119274 138348 119280
rect 138848 119332 138900 119338
rect 138848 119274 138900 119280
rect 138308 113914 138336 119274
rect 138124 113886 138336 113914
rect 139400 113892 139452 113898
rect 137560 112532 137612 112538
rect 137560 112474 137612 112480
rect 138124 99498 138152 113886
rect 139400 113834 139452 113840
rect 138032 99470 138152 99498
rect 138032 96626 138060 99470
rect 138020 96620 138072 96626
rect 138020 96562 138072 96568
rect 138112 89684 138164 89690
rect 138112 89626 138164 89632
rect 138124 86986 138152 89626
rect 138124 86958 138244 86986
rect 138216 12458 138244 86958
rect 138032 12430 138244 12458
rect 137284 7676 137336 7682
rect 137284 7618 137336 7624
rect 136916 3460 136968 3466
rect 136916 3402 136968 3408
rect 137296 480 137324 7618
rect 138032 3534 138060 12430
rect 139412 4894 139440 113834
rect 139504 9042 139532 120006
rect 140056 113898 140084 120006
rect 140792 118998 140820 120006
rect 140780 118992 140832 118998
rect 140780 118934 140832 118940
rect 140792 113914 140820 118934
rect 140044 113892 140096 113898
rect 140792 113886 141004 113914
rect 140044 113834 140096 113840
rect 140780 111920 140832 111926
rect 140780 111862 140832 111868
rect 139492 9036 139544 9042
rect 139492 8978 139544 8984
rect 139676 7812 139728 7818
rect 139676 7754 139728 7760
rect 139400 4888 139452 4894
rect 139400 4830 139452 4836
rect 138480 4480 138532 4486
rect 138480 4422 138532 4428
rect 138020 3528 138072 3534
rect 138020 3470 138072 3476
rect 138492 480 138520 4422
rect 139688 480 139716 7754
rect 140792 3670 140820 111862
rect 140976 99482 141004 113886
rect 141252 111926 141280 120006
rect 142252 118924 142304 118930
rect 142252 118866 142304 118872
rect 141240 111920 141292 111926
rect 141240 111862 141292 111868
rect 140964 99476 141016 99482
rect 140964 99418 141016 99424
rect 140872 99408 140924 99414
rect 140872 99350 140924 99356
rect 140884 95198 140912 99350
rect 140872 95192 140924 95198
rect 140872 95134 140924 95140
rect 140964 86896 141016 86902
rect 140964 86838 141016 86844
rect 140976 84182 141004 86838
rect 140964 84176 141016 84182
rect 140964 84118 141016 84124
rect 141056 74588 141108 74594
rect 141056 74530 141108 74536
rect 141068 58002 141096 74530
rect 140872 57996 140924 58002
rect 140872 57938 140924 57944
rect 141056 57996 141108 58002
rect 141056 57938 141108 57944
rect 140884 57866 140912 57938
rect 140872 57860 140924 57866
rect 140872 57802 140924 57808
rect 140964 48340 141016 48346
rect 140964 48282 141016 48288
rect 140976 48226 141004 48282
rect 140976 48198 141096 48226
rect 141068 38690 141096 48198
rect 140872 38684 140924 38690
rect 140872 38626 140924 38632
rect 141056 38684 141108 38690
rect 141056 38626 141108 38632
rect 140884 38593 140912 38626
rect 140870 38584 140926 38593
rect 140870 38519 140926 38528
rect 140962 29064 141018 29073
rect 140962 28999 141018 29008
rect 140976 28966 141004 28999
rect 140964 28960 141016 28966
rect 140964 28902 141016 28908
rect 140872 19440 140924 19446
rect 140872 19382 140924 19388
rect 140884 19310 140912 19382
rect 140872 19304 140924 19310
rect 140872 19246 140924 19252
rect 141056 9716 141108 9722
rect 141056 9658 141108 9664
rect 141068 7954 141096 9658
rect 141056 7948 141108 7954
rect 141056 7890 141108 7896
rect 140872 7880 140924 7886
rect 140872 7822 140924 7828
rect 140780 3664 140832 3670
rect 140780 3606 140832 3612
rect 140884 480 140912 7822
rect 142068 4888 142120 4894
rect 142068 4830 142120 4836
rect 142080 480 142108 4830
rect 142264 4826 142292 118866
rect 142252 4820 142304 4826
rect 142252 4762 142304 4768
rect 142356 3602 142384 120006
rect 142540 120006 142876 120034
rect 143092 120006 143428 120034
rect 143552 120006 144072 120034
rect 144196 120006 144716 120034
rect 145576 120006 145912 120034
rect 146312 120006 146556 120034
rect 146772 120006 147108 120034
rect 142540 118930 142568 120006
rect 142528 118924 142580 118930
rect 142528 118866 142580 118872
rect 143092 117586 143120 120006
rect 143000 117570 143120 117586
rect 142988 117564 143120 117570
rect 143040 117558 143120 117564
rect 142988 117506 143040 117512
rect 143264 8968 143316 8974
rect 143264 8910 143316 8916
rect 142344 3596 142396 3602
rect 142344 3538 142396 3544
rect 143276 480 143304 8910
rect 143552 3738 143580 120006
rect 143724 117564 143776 117570
rect 143724 117506 143776 117512
rect 143632 109064 143684 109070
rect 143632 109006 143684 109012
rect 143644 9110 143672 109006
rect 143632 9104 143684 9110
rect 143632 9046 143684 9052
rect 143540 3732 143592 3738
rect 143540 3674 143592 3680
rect 143736 3330 143764 117506
rect 144196 109070 144224 120006
rect 145576 118425 145604 120006
rect 145562 118416 145618 118425
rect 145562 118351 145618 118360
rect 144184 109064 144236 109070
rect 144184 109006 144236 109012
rect 145012 96688 145064 96694
rect 145012 96630 145064 96636
rect 145024 89706 145052 96630
rect 145024 89678 145144 89706
rect 145116 67658 145144 89678
rect 145012 67652 145064 67658
rect 145012 67594 145064 67600
rect 145104 67652 145156 67658
rect 145104 67594 145156 67600
rect 145024 64870 145052 67594
rect 145012 64864 145064 64870
rect 145012 64806 145064 64812
rect 144920 55276 144972 55282
rect 144920 55218 144972 55224
rect 144932 47002 144960 55218
rect 144932 46974 145052 47002
rect 145024 46918 145052 46974
rect 145012 46912 145064 46918
rect 145012 46854 145064 46860
rect 144920 46844 144972 46850
rect 144920 46786 144972 46792
rect 144932 22098 144960 46786
rect 144920 22092 144972 22098
rect 144920 22034 144972 22040
rect 145104 22092 145156 22098
rect 145104 22034 145156 22040
rect 145116 4962 145144 22034
rect 145104 4956 145156 4962
rect 145104 4898 145156 4904
rect 145656 4820 145708 4826
rect 145656 4762 145708 4768
rect 144460 3460 144512 3466
rect 144460 3402 144512 3408
rect 143724 3324 143776 3330
rect 143724 3266 143776 3272
rect 144472 480 144500 3402
rect 145668 480 145696 4762
rect 146312 3806 146340 120006
rect 146772 119354 146800 120006
rect 147738 119762 147766 120020
rect 148060 120006 148396 120034
rect 148520 120006 148948 120034
rect 149072 120006 149592 120034
rect 149900 120006 150236 120034
rect 150452 120006 150788 120034
rect 147738 119734 147812 119762
rect 146404 119326 146800 119354
rect 146404 3874 146432 119326
rect 147784 118726 147812 119734
rect 147772 118720 147824 118726
rect 147772 118662 147824 118668
rect 147784 5030 147812 118662
rect 148060 117366 148088 120006
rect 148048 117360 148100 117366
rect 148048 117302 148100 117308
rect 148520 113914 148548 120006
rect 149072 118794 149100 120006
rect 149060 118788 149112 118794
rect 149060 118730 149112 118736
rect 147968 113886 148548 113914
rect 147968 89706 147996 113886
rect 147968 89678 148180 89706
rect 148152 85542 148180 89678
rect 148140 85536 148192 85542
rect 148140 85478 148192 85484
rect 147956 75948 148008 75954
rect 147956 75890 148008 75896
rect 147968 67658 147996 75890
rect 147956 67652 148008 67658
rect 147956 67594 148008 67600
rect 148048 67652 148100 67658
rect 148048 67594 148100 67600
rect 148060 51134 148088 67594
rect 148048 51128 148100 51134
rect 148048 51070 148100 51076
rect 147956 51060 148008 51066
rect 147956 51002 148008 51008
rect 147968 46918 147996 51002
rect 147956 46912 148008 46918
rect 147956 46854 148008 46860
rect 147864 46844 147916 46850
rect 147864 46786 147916 46792
rect 147876 24206 147904 46786
rect 147864 24200 147916 24206
rect 147864 24142 147916 24148
rect 148048 24200 148100 24206
rect 148048 24142 148100 24148
rect 148060 5098 148088 24142
rect 148048 5092 148100 5098
rect 148048 5034 148100 5040
rect 147772 5024 147824 5030
rect 147772 4966 147824 4972
rect 149072 4865 149100 118730
rect 149900 117910 149928 120006
rect 149888 117904 149940 117910
rect 149888 117846 149940 117852
rect 150452 5658 150480 120006
rect 151418 119762 151446 120020
rect 151970 119762 151998 120020
rect 151372 119734 151446 119762
rect 151924 119734 151998 119762
rect 152292 120006 152628 120034
rect 151372 115938 151400 119734
rect 151924 117745 151952 119734
rect 151910 117736 151966 117745
rect 151910 117671 151966 117680
rect 150808 115932 150860 115938
rect 150808 115874 150860 115880
rect 151360 115932 151412 115938
rect 151360 115874 151412 115880
rect 150820 95402 150848 115874
rect 151820 113892 151872 113898
rect 151820 113834 151872 113840
rect 150624 95396 150676 95402
rect 150624 95338 150676 95344
rect 150808 95396 150860 95402
rect 150808 95338 150860 95344
rect 150636 95198 150664 95338
rect 150624 95192 150676 95198
rect 150624 95134 150676 95140
rect 150716 85604 150768 85610
rect 150716 85546 150768 85552
rect 150544 80102 150572 80133
rect 150728 80102 150756 85546
rect 150532 80096 150584 80102
rect 150716 80096 150768 80102
rect 150584 80044 150716 80050
rect 150532 80038 150768 80044
rect 150544 80022 150756 80038
rect 150728 70514 150756 80022
rect 150716 70508 150768 70514
rect 150716 70450 150768 70456
rect 150624 70372 150676 70378
rect 150624 70314 150676 70320
rect 150636 60738 150664 70314
rect 150544 60722 150664 60738
rect 150532 60716 150664 60722
rect 150584 60710 150664 60716
rect 150716 60716 150768 60722
rect 150532 60658 150584 60664
rect 150716 60658 150768 60664
rect 150728 51762 150756 60658
rect 150728 51734 150940 51762
rect 150912 50946 150940 51734
rect 150820 50918 150940 50946
rect 150820 46918 150848 50918
rect 150808 46912 150860 46918
rect 150808 46854 150860 46860
rect 150624 37324 150676 37330
rect 150624 37266 150676 37272
rect 150636 33862 150664 37266
rect 150624 33856 150676 33862
rect 150624 33798 150676 33804
rect 150808 33856 150860 33862
rect 150808 33798 150860 33804
rect 150820 24290 150848 33798
rect 150728 24262 150848 24290
rect 150728 19378 150756 24262
rect 150624 19372 150676 19378
rect 150624 19314 150676 19320
rect 150716 19372 150768 19378
rect 150716 19314 150768 19320
rect 150636 12458 150664 19314
rect 150636 12430 150756 12458
rect 150452 5630 150664 5658
rect 150440 5568 150492 5574
rect 150440 5510 150492 5516
rect 149244 4956 149296 4962
rect 149244 4898 149296 4904
rect 149058 4856 149114 4865
rect 149058 4791 149114 4800
rect 146392 3868 146444 3874
rect 146392 3810 146444 3816
rect 146300 3800 146352 3806
rect 146300 3742 146352 3748
rect 146852 3732 146904 3738
rect 146852 3674 146904 3680
rect 146864 480 146892 3674
rect 148048 2848 148100 2854
rect 148048 2790 148100 2796
rect 148060 480 148088 2790
rect 149256 480 149284 4898
rect 150452 480 150480 5510
rect 150636 3942 150664 5630
rect 150728 5166 150756 12430
rect 151832 9246 151860 113834
rect 151820 9240 151872 9246
rect 151820 9182 151872 9188
rect 150716 5160 150768 5166
rect 150716 5102 150768 5108
rect 151924 4010 151952 117671
rect 152292 113898 152320 120006
rect 153258 119762 153286 120020
rect 153488 120006 153824 120034
rect 154132 120006 154468 120034
rect 154684 120006 155112 120034
rect 155328 120006 155664 120034
rect 156064 120006 156308 120034
rect 156616 120006 156952 120034
rect 157352 120006 157504 120034
rect 157904 120006 158148 120034
rect 153258 119734 153332 119762
rect 152280 113892 152332 113898
rect 152280 113834 152332 113840
rect 153200 113892 153252 113898
rect 153200 113834 153252 113840
rect 152740 5024 152792 5030
rect 152740 4966 152792 4972
rect 151912 4004 151964 4010
rect 151912 3946 151964 3952
rect 150624 3936 150676 3942
rect 150624 3878 150676 3884
rect 151544 3800 151596 3806
rect 151544 3742 151596 3748
rect 151556 480 151584 3742
rect 152752 480 152780 4966
rect 153212 4146 153240 113834
rect 153304 5234 153332 119734
rect 153488 118561 153516 120006
rect 153474 118552 153530 118561
rect 153474 118487 153530 118496
rect 154132 113898 154160 120006
rect 154120 113892 154172 113898
rect 154120 113834 154172 113840
rect 154684 9314 154712 120006
rect 155328 118658 155356 120006
rect 155316 118652 155368 118658
rect 155316 118594 155368 118600
rect 155960 113892 156012 113898
rect 155960 113834 156012 113840
rect 154672 9308 154724 9314
rect 154672 9250 154724 9256
rect 155972 6186 156000 113834
rect 156064 9382 156092 120006
rect 156616 113898 156644 120006
rect 157352 117570 157380 120006
rect 157340 117564 157392 117570
rect 157340 117506 157392 117512
rect 157904 115977 157932 120006
rect 158778 119762 158806 120020
rect 159008 120006 159344 120034
rect 158778 119734 158852 119762
rect 157522 115968 157578 115977
rect 157522 115903 157578 115912
rect 157890 115968 157946 115977
rect 157890 115903 157946 115912
rect 156604 113892 156656 113898
rect 156604 113834 156656 113840
rect 157536 106282 157564 115903
rect 157524 106276 157576 106282
rect 157524 106218 157576 106224
rect 157616 99340 157668 99346
rect 157616 99282 157668 99288
rect 157628 96642 157656 99282
rect 157628 96614 157748 96642
rect 157720 75954 157748 96614
rect 157340 75948 157392 75954
rect 157340 75890 157392 75896
rect 157708 75948 157760 75954
rect 157708 75890 157760 75896
rect 157352 70417 157380 75890
rect 157338 70408 157394 70417
rect 157338 70343 157394 70352
rect 157338 66328 157394 66337
rect 157338 66263 157394 66272
rect 157352 64870 157380 66263
rect 157340 64864 157392 64870
rect 157340 64806 157392 64812
rect 157432 55276 157484 55282
rect 157432 55218 157484 55224
rect 157444 51814 157472 55218
rect 157432 51808 157484 51814
rect 157432 51750 157484 51756
rect 157616 38684 157668 38690
rect 157616 38626 157668 38632
rect 157628 22114 157656 38626
rect 157536 22086 157656 22114
rect 157536 12458 157564 22086
rect 157352 12430 157564 12458
rect 156052 9376 156104 9382
rect 156052 9318 156104 9324
rect 155960 6180 156012 6186
rect 155960 6122 156012 6128
rect 153292 5228 153344 5234
rect 153292 5170 153344 5176
rect 155132 5092 155184 5098
rect 155132 5034 155184 5040
rect 153200 4140 153252 4146
rect 153200 4082 153252 4088
rect 153936 3868 153988 3874
rect 153936 3810 153988 3816
rect 153948 480 153976 3810
rect 155144 480 155172 5034
rect 156328 4140 156380 4146
rect 156328 4082 156380 4088
rect 156340 480 156368 4082
rect 157352 4078 157380 12430
rect 158824 8022 158852 119734
rect 159008 117638 159036 120006
rect 159468 119354 159496 120142
rect 159100 119326 159496 119354
rect 160204 120006 160632 120034
rect 160848 120006 161184 120034
rect 161492 120006 161828 120034
rect 162136 120006 162472 120034
rect 162872 120006 163024 120034
rect 163332 120006 163668 120034
rect 158996 117632 159048 117638
rect 158996 117574 159048 117580
rect 159100 113880 159128 119326
rect 158916 113852 159128 113880
rect 158812 8016 158864 8022
rect 158812 7958 158864 7964
rect 157524 6180 157576 6186
rect 157524 6122 157576 6128
rect 157340 4072 157392 4078
rect 157340 4014 157392 4020
rect 157536 480 157564 6122
rect 158720 5160 158772 5166
rect 158720 5102 158772 5108
rect 158732 480 158760 5102
rect 158916 3398 158944 113852
rect 160204 9450 160232 120006
rect 160848 117842 160876 120006
rect 160836 117836 160888 117842
rect 160836 117778 160888 117784
rect 161388 101448 161440 101454
rect 161388 101390 161440 101396
rect 161400 93022 161428 101390
rect 161388 93016 161440 93022
rect 161388 92958 161440 92964
rect 160192 9444 160244 9450
rect 160192 9386 160244 9392
rect 161492 6254 161520 120006
rect 162136 115977 162164 120006
rect 162872 117774 162900 120006
rect 163332 119354 163360 120006
rect 164298 119762 164326 120020
rect 164528 120006 164864 120034
rect 164298 119734 164372 119762
rect 162964 119326 163360 119354
rect 162860 117768 162912 117774
rect 162860 117710 162912 117716
rect 161754 115968 161810 115977
rect 161754 115903 161810 115912
rect 162122 115968 162178 115977
rect 162122 115903 162178 115912
rect 161768 101454 161796 115903
rect 161756 101448 161808 101454
rect 161756 101390 161808 101396
rect 162964 96694 162992 119326
rect 162952 96688 163004 96694
rect 162952 96630 163004 96636
rect 162860 96620 162912 96626
rect 162860 96562 162912 96568
rect 162872 95198 162900 96562
rect 162860 95192 162912 95198
rect 162860 95134 162912 95140
rect 161664 93016 161716 93022
rect 161664 92958 161716 92964
rect 161676 85542 161704 92958
rect 162952 86896 163004 86902
rect 162952 86838 163004 86844
rect 161664 85536 161716 85542
rect 161664 85478 161716 85484
rect 161756 85536 161808 85542
rect 161756 85478 161808 85484
rect 161768 70310 161796 85478
rect 161756 70304 161808 70310
rect 161756 70246 161808 70252
rect 161756 70168 161808 70174
rect 161756 70110 161808 70116
rect 161768 60874 161796 70110
rect 162964 67794 162992 86838
rect 162952 67788 163004 67794
rect 162952 67730 163004 67736
rect 162952 67652 163004 67658
rect 162952 67594 163004 67600
rect 162964 66230 162992 67594
rect 162952 66224 163004 66230
rect 162952 66166 163004 66172
rect 161676 60846 161796 60874
rect 161676 60738 161704 60846
rect 161584 60722 161704 60738
rect 161572 60716 161704 60722
rect 161624 60710 161704 60716
rect 161756 60716 161808 60722
rect 161572 60658 161624 60664
rect 161756 60658 161808 60664
rect 161768 51134 161796 60658
rect 162952 56636 163004 56642
rect 162952 56578 163004 56584
rect 161756 51128 161808 51134
rect 161756 51070 161808 51076
rect 161756 50924 161808 50930
rect 161756 50866 161808 50872
rect 161768 38570 161796 50866
rect 162964 48634 162992 56578
rect 162872 48606 162992 48634
rect 162872 48346 162900 48606
rect 162860 48340 162912 48346
rect 162860 48282 162912 48288
rect 162952 48340 163004 48346
rect 162952 48282 163004 48288
rect 162964 46918 162992 48282
rect 162952 46912 163004 46918
rect 162952 46854 163004 46860
rect 161768 38542 161888 38570
rect 161860 29034 161888 38542
rect 162952 37324 163004 37330
rect 162952 37266 163004 37272
rect 161756 29028 161808 29034
rect 161756 28970 161808 28976
rect 161848 29028 161900 29034
rect 161848 28970 161900 28976
rect 161768 22778 161796 28970
rect 162964 27606 162992 37266
rect 162952 27600 163004 27606
rect 162952 27542 163004 27548
rect 161756 22772 161808 22778
rect 161756 22714 161808 22720
rect 162952 18012 163004 18018
rect 162952 17954 163004 17960
rect 162964 12510 162992 17954
rect 162952 12504 163004 12510
rect 162952 12446 163004 12452
rect 162860 12436 162912 12442
rect 162860 12378 162912 12384
rect 161756 11892 161808 11898
rect 161756 11834 161808 11840
rect 161768 9518 161796 11834
rect 162872 9654 162900 12378
rect 162860 9648 162912 9654
rect 162860 9590 162912 9596
rect 164344 9586 164372 119734
rect 164528 118522 164556 120006
rect 164988 119354 165016 120142
rect 164620 119326 165016 119354
rect 165724 120006 166152 120034
rect 166368 120006 166704 120034
rect 167104 120006 167348 120034
rect 167656 120006 167992 120034
rect 168392 120006 168544 120034
rect 168852 120006 169188 120034
rect 169740 120006 169984 120034
rect 164516 118516 164568 118522
rect 164516 118458 164568 118464
rect 164620 113880 164648 119326
rect 164436 113852 164648 113880
rect 164332 9580 164384 9586
rect 164332 9522 164384 9528
rect 161756 9512 161808 9518
rect 161756 9454 161808 9460
rect 164436 6322 164464 113852
rect 164424 6316 164476 6322
rect 164424 6258 164476 6264
rect 161480 6248 161532 6254
rect 161480 6190 161532 6196
rect 165724 5302 165752 120006
rect 166368 117706 166396 120006
rect 166356 117700 166408 117706
rect 166356 117642 166408 117648
rect 167000 113892 167052 113898
rect 167000 113834 167052 113840
rect 167012 5370 167040 113834
rect 167104 8906 167132 120006
rect 167656 113898 167684 120006
rect 168392 117434 168420 120006
rect 168852 119354 168880 120006
rect 168484 119326 168880 119354
rect 168380 117428 168432 117434
rect 168380 117370 168432 117376
rect 167644 113892 167696 113898
rect 167644 113834 167696 113840
rect 168484 12510 168512 119326
rect 169852 113892 169904 113898
rect 169852 113834 169904 113840
rect 168472 12504 168524 12510
rect 168472 12446 168524 12452
rect 168380 9716 168432 9722
rect 168380 9658 168432 9664
rect 167092 8900 167144 8906
rect 167092 8842 167144 8848
rect 168392 6390 168420 9658
rect 169864 8838 169892 113834
rect 169852 8832 169904 8838
rect 169852 8774 169904 8780
rect 168380 6384 168432 6390
rect 168380 6326 168432 6332
rect 169956 5438 169984 120006
rect 170048 120006 170384 120034
rect 170692 120006 171028 120034
rect 171244 120006 171580 120034
rect 171888 120006 172224 120034
rect 172624 120006 172868 120034
rect 173084 120006 173420 120034
rect 173912 120006 174064 120034
rect 174372 120006 174708 120034
rect 175260 120006 175596 120034
rect 170048 118114 170076 120006
rect 170036 118108 170088 118114
rect 170036 118050 170088 118056
rect 170404 118108 170456 118114
rect 170404 118050 170456 118056
rect 169944 5432 169996 5438
rect 169944 5374 169996 5380
rect 167000 5364 167052 5370
rect 167000 5306 167052 5312
rect 165712 5296 165764 5302
rect 165712 5238 165764 5244
rect 167092 5296 167144 5302
rect 167092 5238 167144 5244
rect 163504 5228 163556 5234
rect 163504 5170 163556 5176
rect 161112 4004 161164 4010
rect 161112 3946 161164 3952
rect 159916 3528 159968 3534
rect 159916 3470 159968 3476
rect 158904 3392 158956 3398
rect 158904 3334 158956 3340
rect 159928 480 159956 3470
rect 161124 480 161152 3946
rect 162308 3596 162360 3602
rect 162308 3538 162360 3544
rect 162320 480 162348 3538
rect 163516 480 163544 5170
rect 165620 4344 165672 4350
rect 165620 4286 165672 4292
rect 164700 3936 164752 3942
rect 164700 3878 164752 3884
rect 164712 480 164740 3878
rect 165632 3534 165660 4286
rect 165896 3664 165948 3670
rect 165896 3606 165948 3612
rect 165620 3528 165672 3534
rect 165620 3470 165672 3476
rect 165908 480 165936 3606
rect 167104 480 167132 5238
rect 168288 4276 168340 4282
rect 168288 4218 168340 4224
rect 168196 4004 168248 4010
rect 168196 3946 168248 3952
rect 168208 480 168236 3946
rect 168300 3738 168328 4218
rect 170416 4078 170444 118050
rect 170692 113898 170720 120006
rect 170680 113892 170732 113898
rect 170680 113834 170732 113840
rect 171244 5506 171272 120006
rect 171888 117978 171916 120006
rect 171876 117972 171928 117978
rect 171876 117914 171928 117920
rect 171784 117360 171836 117366
rect 171784 117302 171836 117308
rect 171796 5658 171824 117302
rect 172520 113892 172572 113898
rect 172520 113834 172572 113840
rect 171520 5630 171824 5658
rect 171232 5500 171284 5506
rect 171232 5442 171284 5448
rect 170588 5364 170640 5370
rect 170588 5306 170640 5312
rect 170404 4072 170456 4078
rect 170404 4014 170456 4020
rect 168288 3732 168340 3738
rect 168288 3674 168340 3680
rect 169392 3732 169444 3738
rect 169392 3674 169444 3680
rect 169404 480 169432 3674
rect 170600 480 170628 5306
rect 171520 3874 171548 5630
rect 171692 5500 171744 5506
rect 171692 5442 171744 5448
rect 171508 3868 171560 3874
rect 171508 3810 171560 3816
rect 171704 3806 171732 5442
rect 172532 4758 172560 113834
rect 172624 6458 172652 120006
rect 173084 113898 173112 120006
rect 173912 118182 173940 120006
rect 174372 119354 174400 120006
rect 174004 119326 174400 119354
rect 173900 118176 173952 118182
rect 173900 118118 173952 118124
rect 174004 115938 174032 119326
rect 175278 118008 175334 118017
rect 174544 117972 174596 117978
rect 175278 117943 175334 117952
rect 174544 117914 174596 117920
rect 173992 115932 174044 115938
rect 173992 115874 174044 115880
rect 174360 115932 174412 115938
rect 174360 115874 174412 115880
rect 174372 114510 174400 115874
rect 174360 114504 174412 114510
rect 174360 114446 174412 114452
rect 173072 113892 173124 113898
rect 173072 113834 173124 113840
rect 174176 104916 174228 104922
rect 174176 104858 174228 104864
rect 174188 97238 174216 104858
rect 174176 97232 174228 97238
rect 174176 97174 174228 97180
rect 173900 95260 173952 95266
rect 173900 95202 173952 95208
rect 173912 86986 173940 95202
rect 173912 86958 174032 86986
rect 174004 80186 174032 86958
rect 173912 80158 174032 80186
rect 173912 77330 173940 80158
rect 173912 77302 174032 77330
rect 174004 67658 174032 77302
rect 173992 67652 174044 67658
rect 173992 67594 174044 67600
rect 174084 67516 174136 67522
rect 174084 67458 174136 67464
rect 174096 64870 174124 67458
rect 174084 64864 174136 64870
rect 174084 64806 174136 64812
rect 174268 64864 174320 64870
rect 174268 64806 174320 64812
rect 174280 45626 174308 64806
rect 173992 45620 174044 45626
rect 173992 45562 174044 45568
rect 174268 45620 174320 45626
rect 174268 45562 174320 45568
rect 174004 40730 174032 45562
rect 173992 40724 174044 40730
rect 173992 40666 174044 40672
rect 174084 26308 174136 26314
rect 174084 26250 174136 26256
rect 174096 22166 174124 26250
rect 174084 22160 174136 22166
rect 174084 22102 174136 22108
rect 174084 22024 174136 22030
rect 174084 21966 174136 21972
rect 174096 12458 174124 21966
rect 174004 12430 174124 12458
rect 174004 8770 174032 12430
rect 173992 8764 174044 8770
rect 173992 8706 174044 8712
rect 172612 6452 172664 6458
rect 172612 6394 172664 6400
rect 172520 4752 172572 4758
rect 172520 4694 172572 4700
rect 174556 4146 174584 117914
rect 175292 117706 175320 117943
rect 175280 117700 175332 117706
rect 175280 117642 175332 117648
rect 175464 117700 175516 117706
rect 175464 117642 175516 117648
rect 175372 113892 175424 113898
rect 175372 113834 175424 113840
rect 175384 6594 175412 113834
rect 175476 8702 175504 117642
rect 175464 8696 175516 8702
rect 175464 8638 175516 8644
rect 175372 6588 175424 6594
rect 175372 6530 175424 6536
rect 175568 4690 175596 120006
rect 175660 120006 175904 120034
rect 176212 120006 176548 120034
rect 176764 120006 177100 120034
rect 177408 120006 177744 120034
rect 178144 120006 178388 120034
rect 178604 120006 178940 120034
rect 179432 120006 179584 120034
rect 179892 120006 180228 120034
rect 180780 120006 180932 120034
rect 175660 118318 175688 120006
rect 175924 118516 175976 118522
rect 175924 118458 175976 118464
rect 175648 118312 175700 118318
rect 175648 118254 175700 118260
rect 175556 4684 175608 4690
rect 175556 4626 175608 4632
rect 171784 4140 171836 4146
rect 171784 4082 171836 4088
rect 174544 4140 174596 4146
rect 174544 4082 174596 4088
rect 171692 3800 171744 3806
rect 171692 3742 171744 3748
rect 171796 480 171824 4082
rect 174176 4072 174228 4078
rect 174176 4014 174228 4020
rect 172980 3800 173032 3806
rect 172980 3742 173032 3748
rect 172992 480 173020 3742
rect 174188 480 174216 4014
rect 175936 3942 175964 118458
rect 176016 118312 176068 118318
rect 176016 118254 176068 118260
rect 176028 4010 176056 118254
rect 176212 113898 176240 120006
rect 176200 113892 176252 113898
rect 176200 113834 176252 113840
rect 176764 4622 176792 120006
rect 177408 118250 177436 120006
rect 177396 118244 177448 118250
rect 177396 118186 177448 118192
rect 177304 118176 177356 118182
rect 177304 118118 177356 118124
rect 176752 4616 176804 4622
rect 176752 4558 176804 4564
rect 176016 4004 176068 4010
rect 176016 3946 176068 3952
rect 175924 3936 175976 3942
rect 175924 3878 175976 3884
rect 176568 3868 176620 3874
rect 176568 3810 176620 3816
rect 175372 3528 175424 3534
rect 175372 3470 175424 3476
rect 175384 480 175412 3470
rect 176580 480 176608 3810
rect 177316 3534 177344 118118
rect 178040 113892 178092 113898
rect 178040 113834 178092 113840
rect 178052 4554 178080 113834
rect 178144 6662 178172 120006
rect 178604 113898 178632 120006
rect 179328 118244 179380 118250
rect 179328 118186 179380 118192
rect 178592 113892 178644 113898
rect 178592 113834 178644 113840
rect 178132 6656 178184 6662
rect 178132 6598 178184 6604
rect 178040 4548 178092 4554
rect 178040 4490 178092 4496
rect 177764 4140 177816 4146
rect 177764 4082 177816 4088
rect 177304 3528 177356 3534
rect 177304 3470 177356 3476
rect 177776 480 177804 4082
rect 179340 610 179368 118186
rect 179432 118046 179460 120006
rect 179892 119354 179920 120006
rect 179524 119326 179920 119354
rect 179420 118040 179472 118046
rect 179420 117982 179472 117988
rect 179524 113880 179552 119326
rect 179432 113852 179552 113880
rect 179432 109018 179460 113852
rect 179432 108990 179552 109018
rect 179524 106282 179552 108990
rect 179512 106276 179564 106282
rect 179512 106218 179564 106224
rect 179512 99340 179564 99346
rect 179512 99282 179564 99288
rect 179524 96642 179552 99282
rect 179524 96614 179644 96642
rect 179616 89758 179644 96614
rect 179420 89752 179472 89758
rect 179604 89752 179656 89758
rect 179472 89700 179552 89706
rect 179420 89694 179552 89700
rect 179604 89694 179656 89700
rect 179432 89678 179552 89694
rect 179524 89570 179552 89678
rect 179524 89542 179736 89570
rect 179708 77466 179736 89542
rect 179616 77438 179736 77466
rect 179616 77330 179644 77438
rect 179616 77302 179736 77330
rect 179708 70514 179736 77302
rect 179696 70508 179748 70514
rect 179696 70450 179748 70456
rect 179604 70372 179656 70378
rect 179604 70314 179656 70320
rect 179616 60738 179644 70314
rect 179432 60710 179644 60738
rect 179432 56574 179460 60710
rect 179420 56568 179472 56574
rect 179420 56510 179472 56516
rect 179512 46980 179564 46986
rect 179512 46922 179564 46928
rect 179524 46866 179552 46922
rect 179524 46838 179736 46866
rect 179708 37505 179736 46838
rect 179694 37496 179750 37505
rect 179694 37431 179750 37440
rect 179418 37360 179474 37369
rect 179418 37295 179474 37304
rect 179432 37262 179460 37295
rect 179420 37256 179472 37262
rect 179420 37198 179472 37204
rect 179512 27668 179564 27674
rect 179512 27610 179564 27616
rect 179524 22114 179552 27610
rect 179524 22086 179736 22114
rect 179708 19310 179736 22086
rect 179696 19304 179748 19310
rect 179696 19246 179748 19252
rect 179788 9716 179840 9722
rect 179788 9658 179840 9664
rect 179800 9602 179828 9658
rect 179800 9574 179920 9602
rect 179892 3262 179920 9574
rect 180904 6730 180932 120006
rect 181088 120006 181424 120034
rect 181548 120006 182068 120034
rect 182284 120006 182620 120034
rect 182928 120006 183264 120034
rect 183572 120006 183908 120034
rect 184124 120006 184460 120034
rect 184952 120006 185104 120034
rect 185412 120006 185748 120034
rect 186300 120006 186544 120034
rect 181088 118590 181116 120006
rect 181548 119354 181576 120006
rect 181180 119326 181576 119354
rect 181076 118584 181128 118590
rect 181076 118526 181128 118532
rect 181180 113880 181208 119326
rect 180996 113852 181208 113880
rect 180996 6798 181024 113852
rect 182284 6866 182312 120006
rect 182928 118386 182956 120006
rect 182916 118380 182968 118386
rect 182916 118322 182968 118328
rect 183468 118040 183520 118046
rect 183468 117982 183520 117988
rect 182272 6860 182324 6866
rect 182272 6802 182324 6808
rect 180984 6792 181036 6798
rect 180984 6734 181036 6740
rect 180892 6724 180944 6730
rect 180892 6666 180944 6672
rect 180156 3936 180208 3942
rect 180156 3878 180208 3884
rect 179880 3256 179932 3262
rect 179880 3198 179932 3204
rect 178960 604 179012 610
rect 178960 546 179012 552
rect 179328 604 179380 610
rect 179328 546 179380 552
rect 178972 480 179000 546
rect 180168 480 180196 3878
rect 183480 3330 183508 117982
rect 182548 3324 182600 3330
rect 182548 3266 182600 3272
rect 183468 3324 183520 3330
rect 183468 3266 183520 3272
rect 181352 3256 181404 3262
rect 181352 3198 181404 3204
rect 181364 480 181392 3198
rect 182560 480 182588 3266
rect 183572 3194 183600 120006
rect 184124 115977 184152 120006
rect 184952 118697 184980 120006
rect 185412 119354 185440 120006
rect 185044 119326 185440 119354
rect 184938 118688 184994 118697
rect 184938 118623 184994 118632
rect 183834 115968 183890 115977
rect 183834 115903 183890 115912
rect 184110 115968 184166 115977
rect 184110 115903 184166 115912
rect 183848 109018 183876 115903
rect 185044 113880 185072 119326
rect 186044 118380 186096 118386
rect 186044 118322 186096 118328
rect 185676 117904 185728 117910
rect 185676 117846 185728 117852
rect 185584 117768 185636 117774
rect 185584 117710 185636 117716
rect 183756 108990 183876 109018
rect 184952 113852 185072 113880
rect 183756 101266 183784 108990
rect 183664 101238 183784 101266
rect 183664 89758 183692 101238
rect 183652 89752 183704 89758
rect 183652 89694 183704 89700
rect 183744 89616 183796 89622
rect 183744 89558 183796 89564
rect 183756 75954 183784 89558
rect 183744 75948 183796 75954
rect 183744 75890 183796 75896
rect 183836 75948 183888 75954
rect 183836 75890 183888 75896
rect 183848 70802 183876 75890
rect 183756 70774 183876 70802
rect 183756 60738 183784 70774
rect 183664 60722 183784 60738
rect 183652 60716 183784 60722
rect 183704 60710 183784 60716
rect 183836 60716 183888 60722
rect 183652 60658 183704 60664
rect 183836 60658 183888 60664
rect 183848 48346 183876 60658
rect 183836 48340 183888 48346
rect 183836 48282 183888 48288
rect 183928 48340 183980 48346
rect 183928 48282 183980 48288
rect 183940 45558 183968 48282
rect 183928 45552 183980 45558
rect 183928 45494 183980 45500
rect 183744 27668 183796 27674
rect 183744 27610 183796 27616
rect 183756 26246 183784 27610
rect 183744 26240 183796 26246
rect 183744 26182 183796 26188
rect 183836 16652 183888 16658
rect 183836 16594 183888 16600
rect 183848 6050 183876 16594
rect 184952 8090 184980 113852
rect 184940 8084 184992 8090
rect 184940 8026 184992 8032
rect 183836 6044 183888 6050
rect 183836 5986 183888 5992
rect 185596 4078 185624 117710
rect 185688 4146 185716 117846
rect 186056 114594 186084 118322
rect 186056 114566 186176 114594
rect 186148 106350 186176 114566
rect 186412 113892 186464 113898
rect 186412 113834 186464 113840
rect 186136 106344 186188 106350
rect 186136 106286 186188 106292
rect 186228 106208 186280 106214
rect 186228 106150 186280 106156
rect 186240 103494 186268 106150
rect 186228 103488 186280 103494
rect 186228 103430 186280 103436
rect 186320 93900 186372 93906
rect 186320 93842 186372 93848
rect 186332 75954 186360 93842
rect 186228 75948 186280 75954
rect 186228 75890 186280 75896
rect 186320 75948 186372 75954
rect 186320 75890 186372 75896
rect 186240 58002 186268 75890
rect 186228 57996 186280 58002
rect 186228 57938 186280 57944
rect 186320 57928 186372 57934
rect 186320 57870 186372 57876
rect 186332 55214 186360 57870
rect 186320 55208 186372 55214
rect 186320 55150 186372 55156
rect 186228 45620 186280 45626
rect 186228 45562 186280 45568
rect 186240 45506 186268 45562
rect 186240 45478 186360 45506
rect 186332 40730 186360 45478
rect 186320 40724 186372 40730
rect 186320 40666 186372 40672
rect 186228 27124 186280 27130
rect 186228 27066 186280 27072
rect 186240 12510 186268 27066
rect 186228 12504 186280 12510
rect 186228 12446 186280 12452
rect 186044 12436 186096 12442
rect 186044 12378 186096 12384
rect 185676 4140 185728 4146
rect 185676 4082 185728 4088
rect 185584 4072 185636 4078
rect 185584 4014 185636 4020
rect 183744 4004 183796 4010
rect 183744 3946 183796 3952
rect 183560 3188 183612 3194
rect 183560 3130 183612 3136
rect 183756 480 183784 3946
rect 184848 3188 184900 3194
rect 184848 3130 184900 3136
rect 184860 480 184888 3130
rect 186056 480 186084 12378
rect 186424 6225 186452 113834
rect 186410 6216 186466 6225
rect 186410 6151 186466 6160
rect 186516 6118 186544 120006
rect 186608 113898 186636 120226
rect 192128 120142 192464 120170
rect 196268 120142 196696 120170
rect 198108 120142 198536 120170
rect 248892 120142 249412 120170
rect 187068 120006 187496 120034
rect 187712 120006 188140 120034
rect 188448 120006 188784 120034
rect 189184 120006 189336 120034
rect 189644 120006 189980 120034
rect 190472 120006 190624 120034
rect 191024 120006 191176 120034
rect 187068 119354 187096 120006
rect 186700 119326 187096 119354
rect 186596 113892 186648 113898
rect 186596 113834 186648 113840
rect 186700 113778 186728 119326
rect 186608 113750 186728 113778
rect 186504 6112 186556 6118
rect 186504 6054 186556 6060
rect 186608 3126 186636 113750
rect 187712 6526 187740 120006
rect 188448 118153 188476 120006
rect 188434 118144 188490 118153
rect 188434 118079 188490 118088
rect 189080 111580 189132 111586
rect 189080 111522 189132 111528
rect 187700 6520 187752 6526
rect 187700 6462 187752 6468
rect 189092 5982 189120 111522
rect 189184 8158 189212 120006
rect 189644 111586 189672 120006
rect 190368 118584 190420 118590
rect 190368 118526 190420 118532
rect 189632 111580 189684 111586
rect 189632 111522 189684 111528
rect 189172 8152 189224 8158
rect 189172 8094 189224 8100
rect 189080 5976 189132 5982
rect 189080 5918 189132 5924
rect 187240 5432 187292 5438
rect 187240 5374 187292 5380
rect 186596 3120 186648 3126
rect 186596 3062 186648 3068
rect 187252 480 187280 5374
rect 190380 4146 190408 118526
rect 190472 118454 190500 120006
rect 190460 118448 190512 118454
rect 190460 118390 190512 118396
rect 191024 116006 191052 120006
rect 191806 119762 191834 120020
rect 191806 119734 191880 119762
rect 190736 116000 190788 116006
rect 190736 115942 190788 115948
rect 191012 116000 191064 116006
rect 191012 115942 191064 115948
rect 190748 111058 190776 115942
rect 190748 111030 190960 111058
rect 190932 96801 190960 111030
rect 190918 96792 190974 96801
rect 190918 96727 190974 96736
rect 190642 96656 190698 96665
rect 190642 96591 190698 96600
rect 190656 89758 190684 96591
rect 190644 89752 190696 89758
rect 190644 89694 190696 89700
rect 190736 89616 190788 89622
rect 190736 89558 190788 89564
rect 190748 80866 190776 89558
rect 190656 80838 190776 80866
rect 190656 75954 190684 80838
rect 190552 75948 190604 75954
rect 190552 75890 190604 75896
rect 190644 75948 190696 75954
rect 190644 75890 190696 75896
rect 190564 75834 190592 75890
rect 190564 75806 190684 75834
rect 190656 60722 190684 75806
rect 190644 60716 190696 60722
rect 190644 60658 190696 60664
rect 190828 60716 190880 60722
rect 190828 60658 190880 60664
rect 190840 51082 190868 60658
rect 190748 51054 190868 51082
rect 190748 45558 190776 51054
rect 190736 45552 190788 45558
rect 190736 45494 190788 45500
rect 190644 40724 190696 40730
rect 190644 40666 190696 40672
rect 190656 27606 190684 40666
rect 190644 27600 190696 27606
rect 190644 27542 190696 27548
rect 190460 18012 190512 18018
rect 190460 17954 190512 17960
rect 190472 15994 190500 17954
rect 190472 15966 190776 15994
rect 189632 4140 189684 4146
rect 189632 4082 189684 4088
rect 190368 4140 190420 4146
rect 190368 4082 190420 4088
rect 188436 4072 188488 4078
rect 188436 4014 188488 4020
rect 188448 480 188476 4014
rect 189644 480 189672 4082
rect 190748 3058 190776 15966
rect 191852 5914 191880 119734
rect 192128 119406 192156 120142
rect 192680 120006 193016 120034
rect 193232 120006 193660 120034
rect 193968 120006 194304 120034
rect 192116 119400 192168 119406
rect 192036 119360 192116 119388
rect 191932 113892 191984 113898
rect 191932 113834 191984 113840
rect 191944 8226 191972 113834
rect 192036 109070 192064 119360
rect 192116 119342 192168 119348
rect 192680 113898 192708 120006
rect 192668 113892 192720 113898
rect 192668 113834 192720 113840
rect 192024 109064 192076 109070
rect 192024 109006 192076 109012
rect 192208 108996 192260 109002
rect 192208 108938 192260 108944
rect 192220 100042 192248 108938
rect 192220 100014 192340 100042
rect 192312 89758 192340 100014
rect 192300 89752 192352 89758
rect 192300 89694 192352 89700
rect 192392 89616 192444 89622
rect 192392 89558 192444 89564
rect 192404 84182 192432 89558
rect 192392 84176 192444 84182
rect 192392 84118 192444 84124
rect 192208 74588 192260 74594
rect 192208 74530 192260 74536
rect 192220 70514 192248 74530
rect 192208 70508 192260 70514
rect 192208 70450 192260 70456
rect 192116 70372 192168 70378
rect 192116 70314 192168 70320
rect 192128 60858 192156 70314
rect 192116 60852 192168 60858
rect 192116 60794 192168 60800
rect 192116 60716 192168 60722
rect 192116 60658 192168 60664
rect 192128 56574 192156 60658
rect 192116 56568 192168 56574
rect 192116 56510 192168 56516
rect 192116 46980 192168 46986
rect 192116 46922 192168 46928
rect 192128 45898 192156 46922
rect 192116 45892 192168 45898
rect 192116 45834 192168 45840
rect 192208 41336 192260 41342
rect 192208 41278 192260 41284
rect 192220 31754 192248 41278
rect 192208 31748 192260 31754
rect 192208 31690 192260 31696
rect 192208 27600 192260 27606
rect 192208 27542 192260 27548
rect 192220 26246 192248 27542
rect 192208 26240 192260 26246
rect 192208 26182 192260 26188
rect 192208 16652 192260 16658
rect 192208 16594 192260 16600
rect 191932 8220 191984 8226
rect 191932 8162 191984 8168
rect 191840 5908 191892 5914
rect 191840 5850 191892 5856
rect 192220 5846 192248 16594
rect 192208 5840 192260 5846
rect 192208 5782 192260 5788
rect 193232 5778 193260 120006
rect 193968 118289 193996 120006
rect 194842 119762 194870 120020
rect 194796 119734 194870 119762
rect 195164 120006 195500 120034
rect 195992 120006 196144 120034
rect 194508 118448 194560 118454
rect 194508 118390 194560 118396
rect 193954 118280 194010 118289
rect 193954 118215 194010 118224
rect 193864 117564 193916 117570
rect 193864 117506 193916 117512
rect 193220 5772 193272 5778
rect 193220 5714 193272 5720
rect 190828 4140 190880 4146
rect 190828 4082 190880 4088
rect 190736 3052 190788 3058
rect 190736 2994 190788 3000
rect 190840 480 190868 4082
rect 193220 3324 193272 3330
rect 193220 3266 193272 3272
rect 192024 3188 192076 3194
rect 192024 3130 192076 3136
rect 192036 480 192064 3130
rect 193232 480 193260 3266
rect 193876 3126 193904 117506
rect 194416 3392 194468 3398
rect 194416 3334 194468 3340
rect 193864 3120 193916 3126
rect 193864 3062 193916 3068
rect 194428 480 194456 3334
rect 194520 3330 194548 118390
rect 194692 113892 194744 113898
rect 194692 113834 194744 113840
rect 194704 5710 194732 113834
rect 194692 5704 194744 5710
rect 194692 5646 194744 5652
rect 194508 3324 194560 3330
rect 194508 3266 194560 3272
rect 194796 2990 194824 119734
rect 195164 113898 195192 120006
rect 195992 117706 196020 120006
rect 195980 117700 196032 117706
rect 195980 117642 196032 117648
rect 195888 117632 195940 117638
rect 195888 117574 195940 117580
rect 195152 113892 195204 113898
rect 195152 113834 195204 113840
rect 194784 2984 194836 2990
rect 194784 2926 194836 2932
rect 195900 626 195928 117574
rect 196268 116634 196296 120142
rect 197326 119762 197354 120020
rect 197648 120006 197984 120034
rect 197326 119734 197400 119762
rect 197268 117700 197320 117706
rect 197268 117642 197320 117648
rect 196084 116606 196296 116634
rect 196084 7546 196112 116606
rect 196072 7540 196124 7546
rect 196072 7482 196124 7488
rect 197280 3534 197308 117642
rect 197372 5642 197400 119734
rect 197648 117609 197676 120006
rect 197634 117600 197690 117609
rect 197634 117535 197690 117544
rect 198108 116634 198136 120142
rect 197464 116606 198136 116634
rect 198844 120006 199180 120034
rect 199488 120006 199824 120034
rect 200224 120006 200376 120034
rect 200684 120006 201020 120034
rect 198740 116612 198792 116618
rect 197464 7410 197492 116606
rect 198740 116554 198792 116560
rect 197452 7404 197504 7410
rect 197452 7346 197504 7352
rect 198752 7274 198780 116554
rect 198844 7478 198872 120006
rect 199488 116618 199516 120006
rect 199476 116612 199528 116618
rect 199476 116554 199528 116560
rect 200120 116612 200172 116618
rect 200120 116554 200172 116560
rect 198832 7472 198884 7478
rect 198832 7414 198884 7420
rect 198740 7268 198792 7274
rect 198740 7210 198792 7216
rect 200132 7138 200160 116554
rect 200224 7342 200252 120006
rect 200684 116618 200712 120006
rect 201650 119762 201678 120020
rect 201604 119734 201678 119762
rect 201880 120006 202216 120034
rect 202860 120006 203104 120034
rect 201408 117564 201460 117570
rect 201408 117506 201460 117512
rect 200672 116612 200724 116618
rect 200672 116554 200724 116560
rect 200212 7336 200264 7342
rect 200212 7278 200264 7284
rect 200120 7132 200172 7138
rect 200120 7074 200172 7080
rect 197360 5636 197412 5642
rect 197360 5578 197412 5584
rect 201420 3534 201448 117506
rect 201500 116612 201552 116618
rect 201500 116554 201552 116560
rect 201512 7070 201540 116554
rect 201604 7206 201632 119734
rect 201880 116618 201908 120006
rect 201868 116612 201920 116618
rect 201868 116554 201920 116560
rect 202972 116612 203024 116618
rect 202972 116554 203024 116560
rect 202880 114572 202932 114578
rect 202880 114514 202932 114520
rect 202892 7614 202920 114514
rect 202984 7750 203012 116554
rect 203076 8294 203104 120006
rect 203168 120006 203504 120034
rect 203720 120006 204056 120034
rect 204364 120006 204700 120034
rect 204916 120006 205252 120034
rect 205744 120006 205896 120034
rect 206204 120006 206540 120034
rect 203168 114578 203196 120006
rect 203720 116618 203748 120006
rect 203708 116612 203760 116618
rect 203708 116554 203760 116560
rect 204260 116612 204312 116618
rect 204260 116554 204312 116560
rect 203156 114572 203208 114578
rect 203156 114514 203208 114520
rect 203064 8288 203116 8294
rect 203064 8230 203116 8236
rect 202972 7744 203024 7750
rect 202972 7686 203024 7692
rect 202880 7608 202932 7614
rect 202880 7550 202932 7556
rect 201592 7200 201644 7206
rect 201592 7142 201644 7148
rect 201500 7064 201552 7070
rect 201500 7006 201552 7012
rect 203800 4752 203852 4758
rect 203800 4694 203852 4700
rect 196808 3528 196860 3534
rect 196808 3470 196860 3476
rect 197268 3528 197320 3534
rect 197268 3470 197320 3476
rect 200396 3528 200448 3534
rect 200396 3470 200448 3476
rect 201408 3528 201460 3534
rect 201408 3470 201460 3476
rect 195624 598 195928 626
rect 195624 480 195652 598
rect 196820 480 196848 3470
rect 199200 3052 199252 3058
rect 199200 2994 199252 3000
rect 198004 2984 198056 2990
rect 198004 2926 198056 2932
rect 198016 480 198044 2926
rect 199212 480 199240 2994
rect 200408 480 200436 3470
rect 202696 3120 202748 3126
rect 202696 3062 202748 3068
rect 201500 2916 201552 2922
rect 201500 2858 201552 2864
rect 201512 480 201540 2858
rect 202708 480 202736 3062
rect 203812 2922 203840 4694
rect 204168 4616 204220 4622
rect 204168 4558 204220 4564
rect 203892 3188 203944 3194
rect 203892 3130 203944 3136
rect 203800 2916 203852 2922
rect 203800 2858 203852 2864
rect 203904 480 203932 3130
rect 204180 2990 204208 4558
rect 204272 4486 204300 116554
rect 204364 7682 204392 120006
rect 204916 116618 204944 120006
rect 204904 116612 204956 116618
rect 204904 116554 204956 116560
rect 205640 113892 205692 113898
rect 205640 113834 205692 113840
rect 205652 7886 205680 113834
rect 205640 7880 205692 7886
rect 205640 7822 205692 7828
rect 205744 7818 205772 120006
rect 206204 113898 206232 120006
rect 207078 119762 207106 120020
rect 207032 119734 207106 119762
rect 207216 120006 207736 120034
rect 208380 120006 208716 120034
rect 206192 113892 206244 113898
rect 206192 113834 206244 113840
rect 205732 7812 205784 7818
rect 205732 7754 205784 7760
rect 204352 7676 204404 7682
rect 204352 7618 204404 7624
rect 207032 4894 207060 119734
rect 207216 89826 207244 120006
rect 208308 117496 208360 117502
rect 208308 117438 208360 117444
rect 207204 89820 207256 89826
rect 207204 89762 207256 89768
rect 207204 89684 207256 89690
rect 207204 89626 207256 89632
rect 207216 86986 207244 89626
rect 207216 86958 207336 86986
rect 207308 80850 207336 86958
rect 207296 80844 207348 80850
rect 207296 80786 207348 80792
rect 207296 77308 207348 77314
rect 207296 77250 207348 77256
rect 207308 77194 207336 77250
rect 207216 77166 207336 77194
rect 207216 56794 207244 77166
rect 207216 56766 207336 56794
rect 207308 56658 207336 56766
rect 207216 56630 207336 56658
rect 207216 56574 207244 56630
rect 207204 56568 207256 56574
rect 207204 56510 207256 56516
rect 207480 38684 207532 38690
rect 207480 38626 207532 38632
rect 207492 28966 207520 38626
rect 207480 28960 207532 28966
rect 207480 28902 207532 28908
rect 207204 19440 207256 19446
rect 207256 19388 207336 19394
rect 207204 19382 207336 19388
rect 207216 19366 207336 19382
rect 207308 19310 207336 19366
rect 207296 19304 207348 19310
rect 207296 19246 207348 19252
rect 207204 9716 207256 9722
rect 207204 9658 207256 9664
rect 207216 8974 207244 9658
rect 207204 8968 207256 8974
rect 207204 8910 207256 8916
rect 207020 4888 207072 4894
rect 207020 4830 207072 4836
rect 205088 4684 205140 4690
rect 205088 4626 205140 4632
rect 204260 4480 204312 4486
rect 204260 4422 204312 4428
rect 204168 2984 204220 2990
rect 204168 2926 204220 2932
rect 205100 480 205128 4626
rect 208320 3534 208348 117438
rect 208492 113892 208544 113898
rect 208492 113834 208544 113840
rect 208400 12504 208452 12510
rect 208400 12446 208452 12452
rect 208412 4826 208440 12446
rect 208400 4820 208452 4826
rect 208400 4762 208452 4768
rect 208504 4282 208532 113834
rect 208584 99408 208636 99414
rect 208584 99350 208636 99356
rect 208596 12510 208624 99350
rect 208584 12504 208636 12510
rect 208584 12446 208636 12452
rect 208688 4978 208716 120006
rect 208780 120006 208932 120034
rect 209240 120006 209576 120034
rect 209976 120006 210220 120034
rect 210436 120006 210772 120034
rect 211264 120006 211416 120034
rect 211724 120006 212060 120034
rect 208780 99482 208808 120006
rect 209240 113898 209268 120006
rect 209228 113892 209280 113898
rect 209228 113834 209280 113840
rect 209872 113892 209924 113898
rect 209872 113834 209924 113840
rect 208768 99476 208820 99482
rect 208768 99418 208820 99424
rect 208596 4950 208716 4978
rect 209884 4962 209912 113834
rect 209872 4956 209924 4962
rect 208492 4276 208544 4282
rect 208492 4218 208544 4224
rect 207480 3528 207532 3534
rect 207480 3470 207532 3476
rect 208308 3528 208360 3534
rect 208308 3470 208360 3476
rect 206284 2984 206336 2990
rect 206284 2926 206336 2932
rect 206296 480 206324 2926
rect 207492 480 207520 3470
rect 208596 3466 208624 4950
rect 209872 4898 209924 4904
rect 208676 4820 208728 4826
rect 208676 4762 208728 4768
rect 208584 3460 208636 3466
rect 208584 3402 208636 3408
rect 208688 480 208716 4762
rect 209872 3528 209924 3534
rect 209872 3470 209924 3476
rect 209884 480 209912 3470
rect 209976 2854 210004 120006
rect 210436 113898 210464 120006
rect 211068 117428 211120 117434
rect 211068 117370 211120 117376
rect 210424 113892 210476 113898
rect 210424 113834 210476 113840
rect 211080 3534 211108 117370
rect 211160 113892 211212 113898
rect 211160 113834 211212 113840
rect 211172 5506 211200 113834
rect 211264 5574 211292 120006
rect 211724 113898 211752 120006
rect 212598 119762 212626 120020
rect 212920 120006 213256 120034
rect 212598 119734 212672 119762
rect 211712 113892 211764 113898
rect 211712 113834 211764 113840
rect 211252 5568 211304 5574
rect 211252 5510 211304 5516
rect 211160 5500 211212 5506
rect 211160 5442 211212 5448
rect 212644 5030 212672 119734
rect 212920 117366 212948 120006
rect 213886 119762 213914 120020
rect 214024 120006 214452 120034
rect 214576 120006 215096 120034
rect 215312 120006 215740 120034
rect 215956 120006 216292 120034
rect 216692 120006 216936 120034
rect 217336 120006 217580 120034
rect 213886 119734 213960 119762
rect 213828 118312 213880 118318
rect 213828 118254 213880 118260
rect 212908 117360 212960 117366
rect 212908 117302 212960 117308
rect 212632 5024 212684 5030
rect 212632 4966 212684 4972
rect 212264 4888 212316 4894
rect 212264 4830 212316 4836
rect 211068 3528 211120 3534
rect 211068 3470 211120 3476
rect 211068 3256 211120 3262
rect 211068 3198 211120 3204
rect 209964 2848 210016 2854
rect 209964 2790 210016 2796
rect 211080 480 211108 3198
rect 212276 480 212304 4830
rect 213840 626 213868 118254
rect 213932 5098 213960 119734
rect 213920 5092 213972 5098
rect 213920 5034 213972 5040
rect 214024 4418 214052 120006
rect 214576 117450 214604 120006
rect 214208 117422 214604 117450
rect 214208 99482 214236 117422
rect 214564 117360 214616 117366
rect 214564 117302 214616 117308
rect 214196 99476 214248 99482
rect 214196 99418 214248 99424
rect 214104 99408 214156 99414
rect 214104 99350 214156 99356
rect 214116 96626 214144 99350
rect 214104 96620 214156 96626
rect 214104 96562 214156 96568
rect 214288 96620 214340 96626
rect 214288 96562 214340 96568
rect 214300 87009 214328 96562
rect 214102 87000 214158 87009
rect 214102 86935 214158 86944
rect 214286 87000 214342 87009
rect 214286 86935 214342 86944
rect 214116 85542 214144 86935
rect 214104 85536 214156 85542
rect 214104 85478 214156 85484
rect 214104 75948 214156 75954
rect 214104 75890 214156 75896
rect 214116 66230 214144 75890
rect 214104 66224 214156 66230
rect 214104 66166 214156 66172
rect 214104 56636 214156 56642
rect 214104 56578 214156 56584
rect 214116 46918 214144 56578
rect 214104 46912 214156 46918
rect 214104 46854 214156 46860
rect 214104 37324 214156 37330
rect 214104 37266 214156 37272
rect 214116 27606 214144 37266
rect 214104 27600 214156 27606
rect 214104 27542 214156 27548
rect 214196 9716 214248 9722
rect 214196 9658 214248 9664
rect 214208 6186 214236 9658
rect 214196 6180 214248 6186
rect 214196 6122 214248 6128
rect 214012 4412 214064 4418
rect 214012 4354 214064 4360
rect 214576 3466 214604 117302
rect 215312 5166 215340 120006
rect 215956 114578 215984 120006
rect 216692 118114 216720 120006
rect 216680 118108 216732 118114
rect 216680 118050 216732 118056
rect 217336 115977 217364 120006
rect 218118 119762 218146 120020
rect 218440 120006 218776 120034
rect 219420 120006 219664 120034
rect 218118 119734 218192 119762
rect 216954 115968 217010 115977
rect 216954 115903 217010 115912
rect 217322 115968 217378 115977
rect 217322 115903 217378 115912
rect 215392 114572 215444 114578
rect 215392 114514 215444 114520
rect 215944 114572 215996 114578
rect 215944 114514 215996 114520
rect 215404 104854 215432 114514
rect 215392 104848 215444 104854
rect 215392 104790 215444 104796
rect 216968 99362 216996 115903
rect 216784 99334 216996 99362
rect 216784 96626 216812 99334
rect 216772 96620 216824 96626
rect 216772 96562 216824 96568
rect 215392 95260 215444 95266
rect 215392 95202 215444 95208
rect 215404 46918 215432 95202
rect 216864 89548 216916 89554
rect 216864 89490 216916 89496
rect 216876 80170 216904 89490
rect 216864 80164 216916 80170
rect 216864 80106 216916 80112
rect 216864 79960 216916 79966
rect 216864 79902 216916 79908
rect 216876 67590 216904 79902
rect 216864 67584 216916 67590
rect 216864 67526 216916 67532
rect 216864 61056 216916 61062
rect 216864 60998 216916 61004
rect 215392 46912 215444 46918
rect 215392 46854 215444 46860
rect 216876 41426 216904 60998
rect 216784 41398 216904 41426
rect 216784 41290 216812 41398
rect 216784 41262 216904 41290
rect 215392 37324 215444 37330
rect 215392 37266 215444 37272
rect 215404 27606 215432 37266
rect 215392 27600 215444 27606
rect 215392 27542 215444 27548
rect 216876 22114 216904 41262
rect 216784 22086 216904 22114
rect 216784 21978 216812 22086
rect 216784 21950 216904 21978
rect 215484 9716 215536 9722
rect 215484 9658 215536 9664
rect 215496 9602 215524 9658
rect 215496 9574 215616 9602
rect 215300 5160 215352 5166
rect 215300 5102 215352 5108
rect 215588 4350 215616 9574
rect 215852 4956 215904 4962
rect 215852 4898 215904 4904
rect 215576 4344 215628 4350
rect 215576 4286 215628 4292
rect 214564 3460 214616 3466
rect 214564 3402 214616 3408
rect 214656 2916 214708 2922
rect 214656 2858 214708 2864
rect 213472 598 213868 626
rect 213472 480 213500 598
rect 214668 480 214696 2858
rect 215864 480 215892 4898
rect 216876 3602 216904 21950
rect 218164 5234 218192 119734
rect 218440 118658 218468 120006
rect 218428 118652 218480 118658
rect 218428 118594 218480 118600
rect 219256 118108 219308 118114
rect 219256 118050 219308 118056
rect 218152 5228 218204 5234
rect 218152 5170 218204 5176
rect 219268 4078 219296 118050
rect 219532 113892 219584 113898
rect 219532 113834 219584 113840
rect 219544 5302 219572 113834
rect 219532 5296 219584 5302
rect 219532 5238 219584 5244
rect 219348 5024 219400 5030
rect 219348 4966 219400 4972
rect 218152 4072 218204 4078
rect 218152 4014 218204 4020
rect 219256 4072 219308 4078
rect 219256 4014 219308 4020
rect 216864 3596 216916 3602
rect 216864 3538 216916 3544
rect 217048 3460 217100 3466
rect 217048 3402 217100 3408
rect 217060 480 217088 3402
rect 218164 480 218192 4014
rect 219360 480 219388 4966
rect 219636 3670 219664 120006
rect 219728 120006 219972 120034
rect 220280 120006 220616 120034
rect 220832 120006 221260 120034
rect 221476 120006 221812 120034
rect 222212 120006 222456 120034
rect 222764 120006 223008 120034
rect 219728 113898 219756 120006
rect 220280 118522 220308 120006
rect 220268 118516 220320 118522
rect 220268 118458 220320 118464
rect 219992 118244 220044 118250
rect 219992 118186 220044 118192
rect 220004 118130 220032 118186
rect 220004 118102 220124 118130
rect 220096 118046 220124 118102
rect 220084 118040 220136 118046
rect 220084 117982 220136 117988
rect 219716 113892 219768 113898
rect 219716 113834 219768 113840
rect 220728 58676 220780 58682
rect 220728 58618 220780 58624
rect 220740 53961 220768 58618
rect 220726 53952 220782 53961
rect 220726 53887 220782 53896
rect 220832 3738 220860 120006
rect 221476 115977 221504 120006
rect 222212 118250 222240 120006
rect 222764 119354 222792 120006
rect 223638 119762 223666 120020
rect 223960 120006 224296 120034
rect 224512 120006 224848 120034
rect 225156 120006 225492 120034
rect 225800 120006 226136 120034
rect 226444 120006 226688 120034
rect 226996 120006 227332 120034
rect 227732 120006 227976 120034
rect 228100 120006 228528 120034
rect 223638 119734 223712 119762
rect 222396 119326 222792 119354
rect 222200 118244 222252 118250
rect 222200 118186 222252 118192
rect 221002 115968 221058 115977
rect 221002 115903 221058 115912
rect 221462 115968 221518 115977
rect 221462 115903 221518 115912
rect 221016 106282 221044 115903
rect 221004 106276 221056 106282
rect 221004 106218 221056 106224
rect 222396 104904 222424 119326
rect 223684 118318 223712 119734
rect 223672 118312 223724 118318
rect 223672 118254 223724 118260
rect 223960 118182 223988 120006
rect 223948 118176 224000 118182
rect 223948 118118 224000 118124
rect 223488 117972 223540 117978
rect 223488 117914 223540 117920
rect 222304 104876 222424 104904
rect 222304 100706 222332 104876
rect 222292 100700 222344 100706
rect 222292 100642 222344 100648
rect 221004 96688 221056 96694
rect 221004 96630 221056 96636
rect 221016 58682 221044 96630
rect 222568 82884 222620 82890
rect 222568 82826 222620 82832
rect 222580 79506 222608 82826
rect 222488 79478 222608 79506
rect 222488 73234 222516 79478
rect 222384 73228 222436 73234
rect 222384 73170 222436 73176
rect 222476 73228 222528 73234
rect 222476 73170 222528 73176
rect 222396 60738 222424 73170
rect 222304 60710 222424 60738
rect 222304 60602 222332 60710
rect 222304 60574 222424 60602
rect 221004 58676 221056 58682
rect 221004 58618 221056 58624
rect 221002 53952 221058 53961
rect 221002 53887 221058 53896
rect 221016 53825 221044 53887
rect 221002 53816 221058 53825
rect 221002 53751 221058 53760
rect 221186 53816 221242 53825
rect 221186 53751 221242 53760
rect 221200 44198 221228 53751
rect 221004 44192 221056 44198
rect 221004 44134 221056 44140
rect 221188 44192 221240 44198
rect 221188 44134 221240 44140
rect 221016 34513 221044 44134
rect 222396 41426 222424 60574
rect 222304 41398 222424 41426
rect 222304 41290 222332 41398
rect 222304 41262 222424 41290
rect 221002 34504 221058 34513
rect 221002 34439 221058 34448
rect 221186 34504 221242 34513
rect 221186 34439 221242 34448
rect 221200 24886 221228 34439
rect 222396 24954 222424 41262
rect 222384 24948 222436 24954
rect 222384 24890 222436 24896
rect 221004 24880 221056 24886
rect 221004 24822 221056 24828
rect 221188 24880 221240 24886
rect 221188 24822 221240 24828
rect 221016 20126 221044 24822
rect 222292 23520 222344 23526
rect 222292 23462 222344 23468
rect 221004 20120 221056 20126
rect 221004 20062 221056 20068
rect 221004 19984 221056 19990
rect 221004 19926 221056 19932
rect 221016 5370 221044 19926
rect 222304 15230 222332 23462
rect 222292 15224 222344 15230
rect 222292 15166 222344 15172
rect 222384 15156 222436 15162
rect 222384 15098 222436 15104
rect 221004 5364 221056 5370
rect 221004 5306 221056 5312
rect 222396 3874 222424 15098
rect 223500 4078 223528 117914
rect 224512 113150 224540 120006
rect 225156 117910 225184 120006
rect 225800 118046 225828 120006
rect 226248 118176 226300 118182
rect 226248 118118 226300 118124
rect 225788 118040 225840 118046
rect 225788 117982 225840 117988
rect 225144 117904 225196 117910
rect 225144 117846 225196 117852
rect 225604 117428 225656 117434
rect 225604 117370 225656 117376
rect 223672 113144 223724 113150
rect 223672 113086 223724 113092
rect 224500 113144 224552 113150
rect 224500 113086 224552 113092
rect 223684 112010 223712 113086
rect 223638 111982 223712 112010
rect 223638 111874 223666 111982
rect 223638 111846 223712 111874
rect 223684 102134 223712 111846
rect 223672 102128 223724 102134
rect 223672 102070 223724 102076
rect 223764 92540 223816 92546
rect 223764 92482 223816 92488
rect 223776 80170 223804 92482
rect 223764 80164 223816 80170
rect 223764 80106 223816 80112
rect 223672 74588 223724 74594
rect 223672 74530 223724 74536
rect 223684 70394 223712 74530
rect 223592 70366 223712 70394
rect 223592 70258 223620 70366
rect 223592 70230 223712 70258
rect 223684 51202 223712 70230
rect 223672 51196 223724 51202
rect 223672 51138 223724 51144
rect 223672 51060 223724 51066
rect 223672 51002 223724 51008
rect 223684 31890 223712 51002
rect 223672 31884 223724 31890
rect 223672 31826 223724 31832
rect 223580 31748 223632 31754
rect 223580 31690 223632 31696
rect 222936 4072 222988 4078
rect 222936 4014 222988 4020
rect 223488 4072 223540 4078
rect 223488 4014 223540 4020
rect 222384 3868 222436 3874
rect 222384 3810 222436 3816
rect 220820 3732 220872 3738
rect 220820 3674 220872 3680
rect 221740 3732 221792 3738
rect 221740 3674 221792 3680
rect 219624 3664 219676 3670
rect 219624 3606 219676 3612
rect 220544 3256 220596 3262
rect 220544 3198 220596 3204
rect 220556 480 220584 3198
rect 221752 480 221780 3674
rect 222948 480 222976 4014
rect 223592 3602 223620 31690
rect 224132 3664 224184 3670
rect 224132 3606 224184 3612
rect 223580 3596 223632 3602
rect 223580 3538 223632 3544
rect 224144 480 224172 3606
rect 225328 3392 225380 3398
rect 225328 3334 225380 3340
rect 225340 480 225368 3334
rect 225616 3058 225644 117370
rect 226260 3398 226288 118118
rect 226444 3942 226472 120006
rect 226996 117366 227024 120006
rect 227732 118522 227760 120006
rect 228100 119354 228128 120006
rect 229158 119762 229186 120020
rect 229480 120006 229816 120034
rect 230032 120006 230368 120034
rect 230584 120006 231012 120034
rect 231320 120006 231656 120034
rect 231964 120006 232208 120034
rect 232608 120006 232852 120034
rect 233252 120006 233496 120034
rect 233620 120006 234048 120034
rect 229158 119734 229232 119762
rect 227916 119326 228128 119354
rect 227720 118516 227772 118522
rect 227720 118458 227772 118464
rect 227628 118312 227680 118318
rect 227628 118254 227680 118260
rect 226984 117360 227036 117366
rect 226984 117302 227036 117308
rect 227640 4146 227668 118254
rect 227916 104990 227944 119326
rect 229008 118040 229060 118046
rect 229008 117982 229060 117988
rect 227904 104984 227956 104990
rect 227904 104926 227956 104932
rect 227812 104916 227864 104922
rect 227812 104858 227864 104864
rect 227824 99414 227852 104858
rect 227812 99408 227864 99414
rect 227812 99350 227864 99356
rect 227904 99340 227956 99346
rect 227904 99282 227956 99288
rect 227916 92478 227944 99282
rect 227904 92472 227956 92478
rect 227904 92414 227956 92420
rect 228088 82884 228140 82890
rect 228088 82826 228140 82832
rect 228100 74610 228128 82826
rect 228008 74582 228128 74610
rect 228008 73234 228036 74582
rect 227904 73228 227956 73234
rect 227904 73170 227956 73176
rect 227996 73228 228048 73234
rect 227996 73170 228048 73176
rect 227916 60738 227944 73170
rect 227824 60710 227944 60738
rect 227824 60602 227852 60710
rect 227824 60574 227944 60602
rect 227916 41342 227944 60574
rect 227904 41336 227956 41342
rect 227904 41278 227956 41284
rect 228180 41336 228232 41342
rect 228180 41278 228232 41284
rect 228192 34649 228220 41278
rect 227902 34640 227958 34649
rect 227902 34575 227958 34584
rect 228178 34640 228234 34649
rect 228178 34575 228234 34584
rect 227916 34474 227944 34575
rect 227904 34468 227956 34474
rect 227904 34410 227956 34416
rect 227996 34468 228048 34474
rect 227996 34410 228048 34416
rect 228008 20058 228036 34410
rect 227996 20052 228048 20058
rect 227996 19994 228048 20000
rect 227812 6928 227864 6934
rect 227812 6870 227864 6876
rect 226524 4140 226576 4146
rect 226524 4082 226576 4088
rect 227628 4140 227680 4146
rect 227628 4082 227680 4088
rect 227720 4140 227772 4146
rect 227720 4082 227772 4088
rect 226432 3936 226484 3942
rect 226432 3878 226484 3884
rect 226248 3392 226300 3398
rect 226248 3334 226300 3340
rect 225604 3052 225656 3058
rect 225604 2994 225656 3000
rect 226536 480 226564 4082
rect 227732 480 227760 4082
rect 227824 4010 227852 6870
rect 229020 4146 229048 117982
rect 229204 117910 229232 119734
rect 229480 118386 229508 120006
rect 229468 118380 229520 118386
rect 229468 118322 229520 118328
rect 229192 117904 229244 117910
rect 229192 117846 229244 117852
rect 230032 113898 230060 120006
rect 230388 117496 230440 117502
rect 230388 117438 230440 117444
rect 230400 114510 230428 117438
rect 230388 114504 230440 114510
rect 230388 114446 230440 114452
rect 229192 113892 229244 113898
rect 229192 113834 229244 113840
rect 230020 113892 230072 113898
rect 230020 113834 230072 113840
rect 229204 113150 229232 113834
rect 229192 113144 229244 113150
rect 229192 113086 229244 113092
rect 229192 103556 229244 103562
rect 229192 103498 229244 103504
rect 230388 103556 230440 103562
rect 230388 103498 230440 103504
rect 229204 93974 229232 103498
rect 229192 93968 229244 93974
rect 229192 93910 229244 93916
rect 229284 93900 229336 93906
rect 229284 93842 229336 93848
rect 229296 80170 229324 93842
rect 230400 84182 230428 103498
rect 230388 84176 230440 84182
rect 230388 84118 230440 84124
rect 229284 80164 229336 80170
rect 229284 80106 229336 80112
rect 229192 74588 229244 74594
rect 229192 74530 229244 74536
rect 230388 74588 230440 74594
rect 230388 74530 230440 74536
rect 229204 70394 229232 74530
rect 229112 70366 229232 70394
rect 229112 70258 229140 70366
rect 229112 70230 229232 70258
rect 229204 51202 229232 70230
rect 229192 51196 229244 51202
rect 229192 51138 229244 51144
rect 229192 51060 229244 51066
rect 229192 51002 229244 51008
rect 229204 31770 229232 51002
rect 230400 35873 230428 74530
rect 230386 35864 230442 35873
rect 230386 35799 230442 35808
rect 229112 31742 229232 31770
rect 229112 31634 229140 31742
rect 229112 31606 229232 31634
rect 229204 12458 229232 31606
rect 230478 26344 230534 26353
rect 230400 26302 230478 26330
rect 230400 24818 230428 26302
rect 230478 26279 230534 26288
rect 230388 24812 230440 24818
rect 230388 24754 230440 24760
rect 229112 12430 229232 12458
rect 229112 5438 229140 12430
rect 230112 6928 230164 6934
rect 230112 6870 230164 6876
rect 229100 5432 229152 5438
rect 229100 5374 229152 5380
rect 229008 4140 229060 4146
rect 229008 4082 229060 4088
rect 227812 4004 227864 4010
rect 227812 3946 227864 3952
rect 228916 3664 228968 3670
rect 228916 3606 228968 3612
rect 228928 480 228956 3606
rect 230124 480 230152 6870
rect 230584 3806 230612 120006
rect 231320 118590 231348 120006
rect 231308 118584 231360 118590
rect 231308 118526 231360 118532
rect 231768 118380 231820 118386
rect 231768 118322 231820 118328
rect 231124 118244 231176 118250
rect 231124 118186 231176 118192
rect 230662 35728 230718 35737
rect 230662 35663 230718 35672
rect 230676 26353 230704 35663
rect 230662 26344 230718 26353
rect 230662 26279 230718 26288
rect 230572 3800 230624 3806
rect 230572 3742 230624 3748
rect 231136 3126 231164 118186
rect 231780 4146 231808 118322
rect 231308 4140 231360 4146
rect 231308 4082 231360 4088
rect 231768 4140 231820 4146
rect 231768 4082 231820 4088
rect 231124 3120 231176 3126
rect 231124 3062 231176 3068
rect 231320 480 231348 4082
rect 231964 4078 231992 120006
rect 232504 118516 232556 118522
rect 232504 118458 232556 118464
rect 232228 114572 232280 114578
rect 232228 114514 232280 114520
rect 232240 99482 232268 114514
rect 232228 99476 232280 99482
rect 232228 99418 232280 99424
rect 232136 99408 232188 99414
rect 232136 99350 232188 99356
rect 232148 80170 232176 99350
rect 232136 80164 232188 80170
rect 232136 80106 232188 80112
rect 232136 79960 232188 79966
rect 232136 79902 232188 79908
rect 232148 60738 232176 79902
rect 232056 60710 232176 60738
rect 232056 60602 232084 60710
rect 232056 60574 232176 60602
rect 232148 41426 232176 60574
rect 232056 41398 232176 41426
rect 232056 41290 232084 41398
rect 232056 41262 232176 41290
rect 232148 22114 232176 41262
rect 232056 22086 232176 22114
rect 232056 21978 232084 22086
rect 232056 21950 232176 21978
rect 231952 4072 232004 4078
rect 231952 4014 232004 4020
rect 232148 3330 232176 21950
rect 232516 4298 232544 118458
rect 232608 114578 232636 120006
rect 233252 118454 233280 120006
rect 233620 119354 233648 120006
rect 234678 119762 234706 120020
rect 235000 120006 235336 120034
rect 235460 120006 235888 120034
rect 236196 120006 236532 120034
rect 236840 120006 237176 120034
rect 237484 120006 237728 120034
rect 238036 120006 238372 120034
rect 238864 120006 239016 120034
rect 239232 120006 239568 120034
rect 234678 119734 234752 119762
rect 233436 119326 233648 119354
rect 233240 118448 233292 118454
rect 233240 118390 233292 118396
rect 233148 117700 233200 117706
rect 233148 117642 233200 117648
rect 232596 114572 232648 114578
rect 232596 114514 232648 114520
rect 232424 4270 232544 4298
rect 232136 3324 232188 3330
rect 232136 3266 232188 3272
rect 232424 2990 232452 4270
rect 233160 4146 233188 117642
rect 233436 104938 233464 119326
rect 234528 118448 234580 118454
rect 234528 118390 234580 118396
rect 233884 117768 233936 117774
rect 233884 117710 233936 117716
rect 233344 104910 233464 104938
rect 233344 103494 233372 104910
rect 233332 103488 233384 103494
rect 233332 103430 233384 103436
rect 233424 93900 233476 93906
rect 233424 93842 233476 93848
rect 233436 90522 233464 93842
rect 233436 90494 233556 90522
rect 233528 85610 233556 90494
rect 233332 85604 233384 85610
rect 233332 85546 233384 85552
rect 233516 85604 233568 85610
rect 233516 85546 233568 85552
rect 233344 80186 233372 85546
rect 233344 80158 233464 80186
rect 233436 60738 233464 80158
rect 233344 60710 233464 60738
rect 233344 60602 233372 60710
rect 233344 60574 233464 60602
rect 233436 41426 233464 60574
rect 233344 41398 233464 41426
rect 233344 41290 233372 41398
rect 233344 41262 233464 41290
rect 233436 22114 233464 41262
rect 233344 22086 233464 22114
rect 233344 21978 233372 22086
rect 233344 21950 233464 21978
rect 232504 4140 232556 4146
rect 232504 4082 232556 4088
rect 233148 4140 233200 4146
rect 233148 4082 233200 4088
rect 232412 2984 232464 2990
rect 232412 2926 232464 2932
rect 232516 480 232544 4082
rect 233436 3874 233464 21950
rect 233700 4140 233752 4146
rect 233700 4082 233752 4088
rect 233424 3868 233476 3874
rect 233424 3810 233476 3816
rect 233712 480 233740 4082
rect 233896 3194 233924 117710
rect 234540 4146 234568 118390
rect 234724 117842 234752 119734
rect 234712 117836 234764 117842
rect 234712 117778 234764 117784
rect 235000 117638 235028 120006
rect 234988 117632 235040 117638
rect 234988 117574 235040 117580
rect 235460 116634 235488 120006
rect 236196 117910 236224 120006
rect 236184 117904 236236 117910
rect 236184 117846 236236 117852
rect 236840 117638 236868 120006
rect 237196 118584 237248 118590
rect 237196 118526 237248 118532
rect 236828 117632 236880 117638
rect 236828 117574 236880 117580
rect 236644 117564 236696 117570
rect 236644 117506 236696 117512
rect 234724 116606 235488 116634
rect 234724 99498 234752 116606
rect 234632 99470 234752 99498
rect 234632 99362 234660 99470
rect 234632 99334 234844 99362
rect 234816 89622 234844 99334
rect 234804 89616 234856 89622
rect 234804 89558 234856 89564
rect 234804 89480 234856 89486
rect 234804 89422 234856 89428
rect 234816 80170 234844 89422
rect 234804 80164 234856 80170
rect 234804 80106 234856 80112
rect 234712 80096 234764 80102
rect 234712 80038 234764 80044
rect 234724 70394 234752 80038
rect 234632 70366 234752 70394
rect 234632 70258 234660 70366
rect 234632 70230 234752 70258
rect 234724 51082 234752 70230
rect 234632 51054 234752 51082
rect 234632 50946 234660 51054
rect 234632 50918 234752 50946
rect 234724 31770 234752 50918
rect 234632 31742 234752 31770
rect 234632 31634 234660 31742
rect 234632 31606 234752 31634
rect 234724 12458 234752 31606
rect 234632 12430 234752 12458
rect 234632 4622 234660 12430
rect 234620 4616 234672 4622
rect 234620 4558 234672 4564
rect 234528 4140 234580 4146
rect 234528 4082 234580 4088
rect 236000 4140 236052 4146
rect 236000 4082 236052 4088
rect 234804 3800 234856 3806
rect 234804 3742 234856 3748
rect 233884 3188 233936 3194
rect 233884 3130 233936 3136
rect 234816 480 234844 3742
rect 236012 480 236040 4082
rect 236656 3942 236684 117506
rect 237208 12510 237236 118526
rect 237288 117904 237340 117910
rect 237288 117846 237340 117852
rect 237300 12578 237328 117846
rect 237288 12572 237340 12578
rect 237288 12514 237340 12520
rect 237196 12504 237248 12510
rect 237196 12446 237248 12452
rect 237104 12436 237156 12442
rect 237104 12378 237156 12384
rect 236644 3936 236696 3942
rect 236644 3878 236696 3884
rect 237116 3210 237144 12378
rect 237196 12368 237248 12374
rect 237196 12310 237248 12316
rect 237208 4146 237236 12310
rect 237484 4758 237512 120006
rect 238036 118250 238064 120006
rect 238024 118244 238076 118250
rect 238024 118186 238076 118192
rect 238668 117836 238720 117842
rect 238668 117778 238720 117784
rect 238024 117496 238076 117502
rect 238024 117438 238076 117444
rect 237472 4752 237524 4758
rect 237472 4694 237524 4700
rect 237196 4140 237248 4146
rect 237196 4082 237248 4088
rect 238036 3262 238064 117438
rect 238680 19310 238708 117778
rect 238864 117774 238892 120006
rect 238852 117768 238904 117774
rect 238852 117710 238904 117716
rect 239232 116634 239260 120006
rect 240198 119762 240226 120020
rect 240428 120006 240764 120034
rect 240888 120006 241408 120034
rect 241716 120006 242052 120034
rect 242268 120006 242604 120034
rect 243004 120006 243248 120034
rect 243556 120006 243892 120034
rect 244292 120006 244444 120034
rect 244568 120006 245088 120034
rect 240198 119734 240272 119762
rect 240244 118522 240272 119734
rect 240232 118516 240284 118522
rect 240232 118458 240284 118464
rect 240048 117700 240100 117706
rect 240048 117642 240100 117648
rect 239404 117360 239456 117366
rect 239404 117302 239456 117308
rect 238864 116606 239260 116634
rect 238864 113098 238892 116606
rect 238864 113070 238984 113098
rect 238956 80186 238984 113070
rect 238864 80158 238984 80186
rect 238864 80050 238892 80158
rect 238864 80022 238984 80050
rect 238956 67590 238984 80022
rect 238944 67584 238996 67590
rect 238944 67526 238996 67532
rect 238944 57996 238996 58002
rect 238944 57938 238996 57944
rect 238956 41426 238984 57938
rect 238864 41398 238984 41426
rect 238864 41290 238892 41398
rect 238864 41262 238984 41290
rect 238956 22234 238984 41262
rect 238944 22228 238996 22234
rect 238944 22170 238996 22176
rect 238944 19372 238996 19378
rect 238944 19314 238996 19320
rect 238668 19304 238720 19310
rect 238668 19246 238720 19252
rect 238392 9716 238444 9722
rect 238392 9658 238444 9664
rect 238024 3256 238076 3262
rect 237116 3182 237236 3210
rect 238024 3198 238076 3204
rect 237208 480 237236 3182
rect 238404 480 238432 9658
rect 238956 4690 238984 19314
rect 238944 4684 238996 4690
rect 238944 4626 238996 4632
rect 239416 2922 239444 117302
rect 240060 4146 240088 117642
rect 240428 117434 240456 120006
rect 240416 117428 240468 117434
rect 240416 117370 240468 117376
rect 240888 116634 240916 120006
rect 240968 118516 241020 118522
rect 240968 118458 241020 118464
rect 240244 116606 240916 116634
rect 240244 100094 240272 116606
rect 240980 116498 241008 118458
rect 241428 117564 241480 117570
rect 241428 117506 241480 117512
rect 240796 116470 241008 116498
rect 240232 100088 240284 100094
rect 240232 100030 240284 100036
rect 240324 95260 240376 95266
rect 240324 95202 240376 95208
rect 240336 80170 240364 95202
rect 240324 80164 240376 80170
rect 240324 80106 240376 80112
rect 240232 80096 240284 80102
rect 240232 80038 240284 80044
rect 240244 70394 240272 80038
rect 240152 70366 240272 70394
rect 240152 70258 240180 70366
rect 240152 70230 240272 70258
rect 240244 51082 240272 70230
rect 240152 51054 240272 51082
rect 240152 50946 240180 51054
rect 240152 50918 240272 50946
rect 240244 31770 240272 50918
rect 240152 31742 240272 31770
rect 240152 31634 240180 31742
rect 240152 31606 240272 31634
rect 240244 12458 240272 31606
rect 240152 12430 240272 12458
rect 240152 4826 240180 12430
rect 240140 4820 240192 4826
rect 240140 4762 240192 4768
rect 240796 4298 240824 116470
rect 240704 4270 240824 4298
rect 239588 4140 239640 4146
rect 239588 4082 239640 4088
rect 240048 4140 240100 4146
rect 240048 4082 240100 4088
rect 239404 2916 239456 2922
rect 239404 2858 239456 2864
rect 239600 480 239628 4082
rect 240704 3738 240732 4270
rect 241440 4146 241468 117506
rect 241716 117502 241744 120006
rect 242268 117638 242296 120006
rect 242256 117632 242308 117638
rect 242256 117574 242308 117580
rect 241704 117496 241756 117502
rect 241704 117438 241756 117444
rect 243004 4894 243032 120006
rect 243556 118658 243584 120006
rect 243544 118652 243596 118658
rect 243544 118594 243596 118600
rect 244188 117632 244240 117638
rect 244188 117574 244240 117580
rect 243544 117428 243596 117434
rect 243544 117370 243596 117376
rect 242992 4888 243044 4894
rect 242992 4830 243044 4836
rect 240784 4140 240836 4146
rect 240784 4082 240836 4088
rect 241428 4140 241480 4146
rect 241428 4082 241480 4088
rect 243176 4140 243228 4146
rect 243176 4082 243228 4088
rect 240692 3732 240744 3738
rect 240692 3674 240744 3680
rect 240796 480 240824 4082
rect 241980 4072 242032 4078
rect 241980 4014 242032 4020
rect 241992 480 242020 4014
rect 243188 480 243216 4082
rect 243556 4078 243584 117370
rect 243634 117328 243690 117337
rect 243634 117263 243690 117272
rect 243544 4072 243596 4078
rect 243544 4014 243596 4020
rect 243648 3466 243676 117263
rect 244200 4146 244228 117574
rect 244292 117366 244320 120006
rect 244568 119354 244596 120006
rect 245718 119762 245746 120020
rect 245948 120006 246284 120034
rect 246500 120006 246928 120034
rect 247236 120006 247572 120034
rect 247788 120006 248124 120034
rect 248524 120006 248768 120034
rect 245718 119734 245792 119762
rect 244476 119326 244596 119354
rect 244280 117360 244332 117366
rect 244280 117302 244332 117308
rect 244476 109138 244504 119326
rect 245476 117768 245528 117774
rect 245476 117710 245528 117716
rect 244464 109132 244516 109138
rect 244464 109074 244516 109080
rect 244464 108996 244516 109002
rect 244464 108938 244516 108944
rect 244476 106282 244504 108938
rect 244464 106276 244516 106282
rect 244464 106218 244516 106224
rect 244556 106276 244608 106282
rect 244556 106218 244608 106224
rect 244568 99362 244596 106218
rect 244476 99334 244596 99362
rect 244476 82090 244504 99334
rect 244292 82062 244504 82090
rect 244292 75886 244320 82062
rect 244280 75880 244332 75886
rect 244280 75822 244332 75828
rect 244372 70304 244424 70310
rect 244372 70246 244424 70252
rect 244384 60722 244412 70246
rect 244372 60716 244424 60722
rect 244372 60658 244424 60664
rect 244556 60716 244608 60722
rect 244556 60658 244608 60664
rect 244568 38690 244596 60658
rect 244280 38684 244332 38690
rect 244280 38626 244332 38632
rect 244556 38684 244608 38690
rect 244556 38626 244608 38632
rect 244292 37262 244320 38626
rect 244280 37256 244332 37262
rect 244280 37198 244332 37204
rect 244372 31680 244424 31686
rect 244372 31622 244424 31628
rect 244384 22098 244412 31622
rect 244372 22092 244424 22098
rect 244372 22034 244424 22040
rect 244556 22092 244608 22098
rect 244556 22034 244608 22040
rect 244568 4962 244596 22034
rect 244556 4956 244608 4962
rect 244556 4898 244608 4904
rect 244188 4140 244240 4146
rect 244188 4082 244240 4088
rect 243636 3460 243688 3466
rect 243636 3402 243688 3408
rect 245488 3330 245516 117710
rect 245568 117496 245620 117502
rect 245568 117438 245620 117444
rect 244372 3324 244424 3330
rect 244372 3266 244424 3272
rect 245476 3324 245528 3330
rect 245476 3266 245528 3272
rect 244384 480 244412 3266
rect 245580 480 245608 117438
rect 245764 117337 245792 119734
rect 245948 118114 245976 120006
rect 246500 119354 246528 120006
rect 246040 119326 246528 119354
rect 245936 118108 245988 118114
rect 245936 118050 245988 118056
rect 245750 117328 245806 117337
rect 245750 117263 245806 117272
rect 246040 113914 246068 119326
rect 247236 117434 247264 120006
rect 247788 118522 247816 120006
rect 247776 118516 247828 118522
rect 247776 118458 247828 118464
rect 248328 118108 248380 118114
rect 248328 118050 248380 118056
rect 247224 117428 247276 117434
rect 247224 117370 247276 117376
rect 247684 117428 247736 117434
rect 247684 117370 247736 117376
rect 245948 113886 246068 113914
rect 245948 77314 245976 113886
rect 245752 77308 245804 77314
rect 245752 77250 245804 77256
rect 245936 77308 245988 77314
rect 245936 77250 245988 77256
rect 245764 75886 245792 77250
rect 245752 75880 245804 75886
rect 245752 75822 245804 75828
rect 245844 70372 245896 70378
rect 245844 70314 245896 70320
rect 245856 60722 245884 70314
rect 245844 60716 245896 60722
rect 245844 60658 245896 60664
rect 246028 60716 246080 60722
rect 246028 60658 246080 60664
rect 246040 50674 246068 60658
rect 246040 50646 246160 50674
rect 246132 50402 246160 50646
rect 246040 50374 246160 50402
rect 246040 38690 246068 50374
rect 245752 38684 245804 38690
rect 245752 38626 245804 38632
rect 246028 38684 246080 38690
rect 246028 38626 246080 38632
rect 245764 37262 245792 38626
rect 245752 37256 245804 37262
rect 245752 37198 245804 37204
rect 245844 31680 245896 31686
rect 245844 31622 245896 31628
rect 245856 22098 245884 31622
rect 245844 22092 245896 22098
rect 245844 22034 245896 22040
rect 246028 22092 246080 22098
rect 246028 22034 246080 22040
rect 246040 12050 246068 22034
rect 246040 12022 246160 12050
rect 246132 11778 246160 12022
rect 246040 11750 246160 11778
rect 246040 5030 246068 11750
rect 246028 5024 246080 5030
rect 246028 4966 246080 4972
rect 247696 3670 247724 117370
rect 248340 115938 248368 118050
rect 248524 117978 248552 120006
rect 248892 119354 248920 120142
rect 248616 119326 248920 119354
rect 249812 120006 249964 120034
rect 250272 120006 250608 120034
rect 248512 117972 248564 117978
rect 248512 117914 248564 117920
rect 248328 115932 248380 115938
rect 248328 115874 248380 115880
rect 248420 115932 248472 115938
rect 248420 115874 248472 115880
rect 248432 114510 248460 115874
rect 248420 114504 248472 114510
rect 248420 114446 248472 114452
rect 248616 109018 248644 119326
rect 249812 118182 249840 120006
rect 250272 118318 250300 120006
rect 251238 119762 251266 120020
rect 251468 120006 251804 120034
rect 252112 120006 252448 120034
rect 252756 120006 253092 120034
rect 253308 120006 253644 120034
rect 253952 120006 254288 120034
rect 254596 120006 254932 120034
rect 255332 120006 255484 120034
rect 255792 120006 256128 120034
rect 251238 119734 251312 119762
rect 250260 118312 250312 118318
rect 250260 118254 250312 118260
rect 250536 118312 250588 118318
rect 250536 118254 250588 118260
rect 249800 118176 249852 118182
rect 249800 118118 249852 118124
rect 249708 117972 249760 117978
rect 249708 117914 249760 117920
rect 248524 108990 248644 109018
rect 248328 104916 248380 104922
rect 248328 104858 248380 104864
rect 248340 104802 248368 104858
rect 248340 104774 248460 104802
rect 248432 100094 248460 104774
rect 248420 100088 248472 100094
rect 248420 100030 248472 100036
rect 248524 99414 248552 108990
rect 248512 99408 248564 99414
rect 248512 99350 248564 99356
rect 248420 99340 248472 99346
rect 248420 99282 248472 99288
rect 248432 96665 248460 99282
rect 248418 96656 248474 96665
rect 248418 96591 248474 96600
rect 248602 96656 248658 96665
rect 248602 96591 248658 96600
rect 248328 95260 248380 95266
rect 248328 95202 248380 95208
rect 248340 57934 248368 95202
rect 248616 87038 248644 96591
rect 248604 87032 248656 87038
rect 248604 86974 248656 86980
rect 248788 86896 248840 86902
rect 248788 86838 248840 86844
rect 248800 84182 248828 86838
rect 248788 84176 248840 84182
rect 248788 84118 248840 84124
rect 248420 74588 248472 74594
rect 248420 74530 248472 74536
rect 248432 70258 248460 74530
rect 248432 70230 248552 70258
rect 248524 60738 248552 70230
rect 248432 60722 248552 60738
rect 248420 60716 248552 60722
rect 248472 60710 248552 60716
rect 248604 60716 248656 60722
rect 248420 60658 248472 60664
rect 248604 60658 248656 60664
rect 248236 57928 248288 57934
rect 248236 57870 248288 57876
rect 248328 57928 248380 57934
rect 248328 57870 248380 57876
rect 248248 48362 248276 57870
rect 248616 53122 248644 60658
rect 248616 53094 248920 53122
rect 248248 48334 248368 48362
rect 248340 46918 248368 48334
rect 248328 46912 248380 46918
rect 248328 46854 248380 46860
rect 248892 42090 248920 53094
rect 248696 42084 248748 42090
rect 248696 42026 248748 42032
rect 248880 42084 248932 42090
rect 248880 42026 248932 42032
rect 248328 37324 248380 37330
rect 248328 37266 248380 37272
rect 248340 12510 248368 37266
rect 248708 27674 248736 42026
rect 248512 27668 248564 27674
rect 248512 27610 248564 27616
rect 248696 27668 248748 27674
rect 248696 27610 248748 27616
rect 248524 22114 248552 27610
rect 248432 22098 248552 22114
rect 248420 22092 248552 22098
rect 248472 22086 248552 22092
rect 248604 22092 248656 22098
rect 248420 22034 248472 22040
rect 248604 22034 248656 22040
rect 248328 12504 248380 12510
rect 248328 12446 248380 12452
rect 247960 12436 248012 12442
rect 247960 12378 248012 12384
rect 247684 3664 247736 3670
rect 247684 3606 247736 3612
rect 246764 3256 246816 3262
rect 246764 3198 246816 3204
rect 246776 480 246804 3198
rect 247972 480 248000 12378
rect 248616 12050 248644 22034
rect 248616 12022 248736 12050
rect 248708 11778 248736 12022
rect 248616 11750 248736 11778
rect 248616 3602 248644 11750
rect 248604 3596 248656 3602
rect 248604 3538 248656 3544
rect 249720 3330 249748 117914
rect 250444 117360 250496 117366
rect 250444 117302 250496 117308
rect 250456 3806 250484 117302
rect 250444 3800 250496 3806
rect 250444 3742 250496 3748
rect 250352 3392 250404 3398
rect 250352 3334 250404 3340
rect 249156 3324 249208 3330
rect 249156 3266 249208 3272
rect 249708 3324 249760 3330
rect 249708 3266 249760 3272
rect 249168 480 249196 3266
rect 250364 480 250392 3334
rect 250548 3262 250576 118254
rect 251088 118176 251140 118182
rect 251088 118118 251140 118124
rect 251100 3398 251128 118118
rect 251284 118046 251312 119734
rect 251272 118040 251324 118046
rect 251272 117982 251324 117988
rect 251468 117434 251496 120006
rect 252112 118250 252140 120006
rect 252756 118386 252784 120006
rect 253308 118658 253336 120006
rect 253296 118652 253348 118658
rect 253296 118594 253348 118600
rect 253952 118454 253980 120006
rect 253940 118448 253992 118454
rect 253940 118390 253992 118396
rect 252744 118380 252796 118386
rect 252744 118322 252796 118328
rect 252100 118244 252152 118250
rect 252100 118186 252152 118192
rect 251456 117428 251508 117434
rect 251456 117370 251508 117376
rect 252468 117428 252520 117434
rect 252468 117370 252520 117376
rect 252480 4146 252508 117370
rect 254596 117366 254624 120006
rect 255332 118590 255360 120006
rect 255320 118584 255372 118590
rect 255320 118526 255372 118532
rect 254676 118244 254728 118250
rect 254676 118186 254728 118192
rect 254584 117360 254636 117366
rect 254584 117302 254636 117308
rect 254688 115682 254716 118186
rect 255228 118040 255280 118046
rect 255228 117982 255280 117988
rect 254596 115654 254716 115682
rect 251456 4140 251508 4146
rect 251456 4082 251508 4088
rect 252468 4140 252520 4146
rect 252468 4082 252520 4088
rect 251088 3392 251140 3398
rect 251088 3334 251140 3340
rect 250536 3256 250588 3262
rect 250536 3198 250588 3204
rect 251468 480 251496 4082
rect 253848 3324 253900 3330
rect 253848 3266 253900 3272
rect 252652 3052 252704 3058
rect 252652 2994 252704 3000
rect 252664 480 252692 2994
rect 253860 480 253888 3266
rect 254596 3058 254624 115654
rect 255240 3346 255268 117982
rect 255792 117910 255820 120006
rect 256758 119762 256786 120020
rect 256712 119734 256786 119762
rect 256988 120006 257324 120034
rect 257632 120006 257968 120034
rect 258276 120006 258520 120034
rect 258828 120006 259164 120034
rect 259472 120006 259808 120034
rect 260024 120006 260360 120034
rect 260852 120006 261004 120034
rect 261312 120006 261648 120034
rect 256608 118448 256660 118454
rect 256608 118390 256660 118396
rect 255780 117904 255832 117910
rect 255780 117846 255832 117852
rect 256620 3346 256648 118390
rect 256712 117842 256740 119734
rect 256700 117836 256752 117842
rect 256700 117778 256752 117784
rect 256988 117706 257016 120006
rect 257344 118584 257396 118590
rect 257344 118526 257396 118532
rect 256976 117700 257028 117706
rect 256976 117642 257028 117648
rect 255056 3318 255268 3346
rect 256252 3318 256648 3346
rect 257356 3330 257384 118526
rect 257632 117570 257660 120006
rect 258276 118658 258304 120006
rect 258264 118652 258316 118658
rect 258264 118594 258316 118600
rect 257988 118380 258040 118386
rect 257988 118322 258040 118328
rect 257620 117564 257672 117570
rect 257620 117506 257672 117512
rect 258000 3534 258028 118322
rect 258828 117638 258856 120006
rect 259472 117774 259500 120006
rect 259460 117768 259512 117774
rect 259460 117710 259512 117716
rect 258816 117632 258868 117638
rect 258816 117574 258868 117580
rect 260024 117502 260052 120006
rect 260852 118318 260880 120006
rect 260840 118312 260892 118318
rect 260840 118254 260892 118260
rect 261312 118114 261340 120006
rect 262186 119762 262214 120020
rect 262508 120006 262844 120034
rect 263152 120006 263488 120034
rect 263704 120006 264040 120034
rect 264348 120006 264684 120034
rect 264992 120006 265328 120034
rect 265544 120006 265880 120034
rect 266372 120006 266524 120034
rect 266832 120006 267168 120034
rect 262186 119734 262260 119762
rect 261300 118108 261352 118114
rect 261300 118050 261352 118056
rect 262128 118040 262180 118046
rect 262128 117982 262180 117988
rect 261484 117700 261536 117706
rect 261484 117642 261536 117648
rect 260012 117496 260064 117502
rect 260012 117438 260064 117444
rect 259368 117360 259420 117366
rect 259368 117302 259420 117308
rect 257436 3528 257488 3534
rect 257436 3470 257488 3476
rect 257988 3528 258040 3534
rect 257988 3470 258040 3476
rect 257344 3324 257396 3330
rect 254584 3052 254636 3058
rect 254584 2994 254636 3000
rect 255056 480 255084 3318
rect 256252 480 256280 3318
rect 257344 3266 257396 3272
rect 257448 480 257476 3470
rect 259380 3126 259408 117302
rect 261496 3534 261524 117642
rect 259828 3528 259880 3534
rect 259828 3470 259880 3476
rect 261484 3528 261536 3534
rect 261484 3470 261536 3476
rect 258632 3120 258684 3126
rect 258632 3062 258684 3068
rect 259368 3120 259420 3126
rect 259368 3062 259420 3068
rect 258644 480 258672 3062
rect 259840 480 259868 3470
rect 262140 3262 262168 117982
rect 262232 117978 262260 119734
rect 262508 118182 262536 120006
rect 262496 118176 262548 118182
rect 262496 118118 262548 118124
rect 262220 117972 262272 117978
rect 262220 117914 262272 117920
rect 263152 117434 263180 120006
rect 263704 118250 263732 120006
rect 264348 118590 264376 120006
rect 264336 118584 264388 118590
rect 264336 118526 264388 118532
rect 263692 118244 263744 118250
rect 263692 118186 263744 118192
rect 264992 118114 265020 120006
rect 265544 118454 265572 120006
rect 265532 118448 265584 118454
rect 265532 118390 265584 118396
rect 266372 118386 266400 120006
rect 266360 118380 266412 118386
rect 266360 118322 266412 118328
rect 264980 118108 265032 118114
rect 264980 118050 265032 118056
rect 263508 117972 263560 117978
rect 263508 117914 263560 117920
rect 263416 117904 263468 117910
rect 263416 117846 263468 117852
rect 263140 117428 263192 117434
rect 263140 117370 263192 117376
rect 262220 3528 262272 3534
rect 262220 3470 262272 3476
rect 261024 3256 261076 3262
rect 261024 3198 261076 3204
rect 262128 3256 262180 3262
rect 262128 3198 262180 3204
rect 261036 480 261064 3198
rect 262232 480 262260 3470
rect 263428 480 263456 117846
rect 263520 3534 263548 117914
rect 266268 117564 266320 117570
rect 266268 117506 266320 117512
rect 266280 4146 266308 117506
rect 266832 117366 266860 120006
rect 267706 119762 267734 120020
rect 268028 120006 268364 120034
rect 268672 120006 269008 120034
rect 269224 120006 269560 120034
rect 269868 120006 270204 120034
rect 270512 120006 270848 120034
rect 271064 120006 271400 120034
rect 271892 120006 272044 120034
rect 272444 120006 272688 120034
rect 273240 120006 273392 120034
rect 267706 119734 267780 119762
rect 267752 117706 267780 119734
rect 268028 118046 268056 120006
rect 268016 118040 268068 118046
rect 268016 117982 268068 117988
rect 268672 117978 268700 120006
rect 268660 117972 268712 117978
rect 268660 117914 268712 117920
rect 269224 117910 269252 120006
rect 269212 117904 269264 117910
rect 269212 117846 269264 117852
rect 267740 117700 267792 117706
rect 267740 117642 267792 117648
rect 267648 117496 267700 117502
rect 267648 117438 267700 117444
rect 266820 117360 266872 117366
rect 266820 117302 266872 117308
rect 265808 4140 265860 4146
rect 265808 4082 265860 4088
rect 266268 4140 266320 4146
rect 266268 4082 266320 4088
rect 263508 3528 263560 3534
rect 263508 3470 263560 3476
rect 264612 3120 264664 3126
rect 264612 3062 264664 3068
rect 264624 480 264652 3062
rect 265820 480 265848 4082
rect 267660 3330 267688 117438
rect 269764 117428 269816 117434
rect 269764 117370 269816 117376
rect 268384 117360 268436 117366
rect 268384 117302 268436 117308
rect 268108 4140 268160 4146
rect 268108 4082 268160 4088
rect 267004 3324 267056 3330
rect 267004 3266 267056 3272
rect 267648 3324 267700 3330
rect 267648 3266 267700 3272
rect 267016 480 267044 3266
rect 268120 480 268148 4082
rect 268396 3126 268424 117302
rect 269776 4146 269804 117370
rect 269868 117366 269896 120006
rect 270512 117570 270540 120006
rect 270500 117564 270552 117570
rect 270500 117506 270552 117512
rect 271064 117502 271092 120006
rect 271052 117496 271104 117502
rect 271052 117438 271104 117444
rect 271892 117434 271920 120006
rect 271880 117428 271932 117434
rect 271880 117370 271932 117376
rect 269856 117360 269908 117366
rect 269856 117302 269908 117308
rect 272444 116006 272472 120006
rect 272524 117428 272576 117434
rect 272524 117370 272576 117376
rect 272248 116000 272300 116006
rect 272248 115942 272300 115948
rect 272432 116000 272484 116006
rect 272432 115942 272484 115948
rect 272260 109018 272288 115942
rect 272076 108990 272288 109018
rect 272076 95282 272104 108990
rect 271984 95254 272104 95282
rect 271984 95198 272012 95254
rect 271972 95192 272024 95198
rect 271972 95134 272024 95140
rect 272064 85604 272116 85610
rect 272064 85546 272116 85552
rect 272076 85490 272104 85546
rect 272076 85462 272196 85490
rect 272168 80782 272196 85462
rect 271880 80776 271932 80782
rect 271880 80718 271932 80724
rect 272156 80776 272208 80782
rect 272156 80718 272208 80724
rect 271892 75886 271920 80718
rect 271880 75880 271932 75886
rect 271880 75822 271932 75828
rect 271972 66292 272024 66298
rect 271972 66234 272024 66240
rect 271984 60722 272012 66234
rect 271972 60716 272024 60722
rect 271972 60658 272024 60664
rect 272156 60716 272208 60722
rect 272156 60658 272208 60664
rect 272168 51134 272196 60658
rect 272156 51128 272208 51134
rect 272156 51070 272208 51076
rect 272064 51060 272116 51066
rect 272064 51002 272116 51008
rect 272076 48210 272104 51002
rect 272064 48204 272116 48210
rect 272064 48146 272116 48152
rect 271880 41336 271932 41342
rect 271880 41278 271932 41284
rect 271892 38622 271920 41278
rect 271880 38616 271932 38622
rect 271880 38558 271932 38564
rect 271972 29028 272024 29034
rect 271972 28970 272024 28976
rect 271984 28914 272012 28970
rect 271984 28886 272196 28914
rect 269764 4140 269816 4146
rect 269764 4082 269816 4088
rect 271696 4140 271748 4146
rect 271696 4082 271748 4088
rect 269304 4004 269356 4010
rect 269304 3946 269356 3952
rect 268384 3120 268436 3126
rect 268384 3062 268436 3068
rect 269316 480 269344 3946
rect 270500 3460 270552 3466
rect 270500 3402 270552 3408
rect 270512 480 270540 3402
rect 271708 480 271736 4082
rect 272168 4010 272196 28886
rect 272536 4146 272564 117370
rect 273168 117360 273220 117366
rect 273168 117302 273220 117308
rect 272524 4140 272576 4146
rect 272524 4082 272576 4088
rect 272156 4004 272208 4010
rect 272156 3946 272208 3952
rect 273180 610 273208 117302
rect 273364 3466 273392 120006
rect 273548 120006 273884 120034
rect 274192 120006 274528 120034
rect 274652 120006 275080 120034
rect 275388 120006 275724 120034
rect 276124 120006 276276 120034
rect 276920 120006 277348 120034
rect 277564 120006 277900 120034
rect 278116 120006 278452 120034
rect 278760 120006 279096 120034
rect 279404 120006 279740 120034
rect 279956 120006 280108 120034
rect 280600 120006 280936 120034
rect 281244 120006 281488 120034
rect 281796 120006 282132 120034
rect 282440 120006 282776 120034
rect 283084 120006 283420 120034
rect 283636 120006 283972 120034
rect 284280 120006 284616 120034
rect 284924 120006 285260 120034
rect 273548 117434 273576 120006
rect 273536 117428 273588 117434
rect 273536 117370 273588 117376
rect 274192 117366 274220 120006
rect 274180 117360 274232 117366
rect 274652 117314 274680 120006
rect 274180 117302 274232 117308
rect 274560 117286 274680 117314
rect 274560 4146 274588 117286
rect 275388 106321 275416 120006
rect 276124 115938 276152 120006
rect 276020 115932 276072 115938
rect 276020 115874 276072 115880
rect 276112 115932 276164 115938
rect 276112 115874 276164 115880
rect 276032 106457 276060 115874
rect 276018 106448 276074 106457
rect 276018 106383 276074 106392
rect 275006 106312 275062 106321
rect 275006 106247 275062 106256
rect 275374 106312 275430 106321
rect 275374 106247 275430 106256
rect 276110 106312 276166 106321
rect 276110 106247 276166 106256
rect 275020 96665 275048 106247
rect 276124 104854 276152 106247
rect 276112 104848 276164 104854
rect 276112 104790 276164 104796
rect 274730 96656 274786 96665
rect 274730 96591 274786 96600
rect 275006 96656 275062 96665
rect 275006 96591 275062 96600
rect 274744 89706 274772 96591
rect 276112 95260 276164 95266
rect 276112 95202 276164 95208
rect 274744 89678 274864 89706
rect 274836 15910 274864 89678
rect 276124 66230 276152 95202
rect 276112 66224 276164 66230
rect 276112 66166 276164 66172
rect 276296 66224 276348 66230
rect 276296 66166 276348 66172
rect 276308 48385 276336 66166
rect 276110 48376 276166 48385
rect 276110 48311 276166 48320
rect 276294 48376 276350 48385
rect 276294 48311 276350 48320
rect 276124 46918 276152 48311
rect 276112 46912 276164 46918
rect 276112 46854 276164 46860
rect 276112 29096 276164 29102
rect 276112 29038 276164 29044
rect 276124 27606 276152 29038
rect 276112 27600 276164 27606
rect 276112 27542 276164 27548
rect 276112 18012 276164 18018
rect 276112 17954 276164 17960
rect 274824 15904 274876 15910
rect 274824 15846 274876 15852
rect 276124 12510 276152 17954
rect 276112 12504 276164 12510
rect 276112 12446 276164 12452
rect 276480 12368 276532 12374
rect 276480 12310 276532 12316
rect 275284 9716 275336 9722
rect 275284 9658 275336 9664
rect 274088 4140 274140 4146
rect 274088 4082 274140 4088
rect 274548 4140 274600 4146
rect 274548 4082 274600 4088
rect 273352 3460 273404 3466
rect 273352 3402 273404 3408
rect 272892 604 272944 610
rect 272892 546 272944 552
rect 273168 604 273220 610
rect 273168 546 273220 552
rect 272904 480 272932 546
rect 274100 480 274128 4082
rect 275296 480 275324 9658
rect 276492 480 276520 12310
rect 277320 3890 277348 120006
rect 277872 117366 277900 120006
rect 278424 117434 278452 120006
rect 278412 117428 278464 117434
rect 278412 117370 278464 117376
rect 279068 117366 279096 120006
rect 279712 119354 279740 120006
rect 279712 119326 280016 119354
rect 279148 117428 279200 117434
rect 279148 117370 279200 117376
rect 277860 117360 277912 117366
rect 277860 117302 277912 117308
rect 278872 117360 278924 117366
rect 278872 117302 278924 117308
rect 279056 117360 279108 117366
rect 279056 117302 279108 117308
rect 277320 3862 277716 3890
rect 277688 480 277716 3862
rect 278884 480 278912 117302
rect 279160 4026 279188 117370
rect 279988 109018 280016 119326
rect 280080 117570 280108 120006
rect 280068 117564 280120 117570
rect 280068 117506 280120 117512
rect 280908 117366 280936 120006
rect 280344 117360 280396 117366
rect 280344 117302 280396 117308
rect 280896 117360 280948 117366
rect 280896 117302 280948 117308
rect 281356 117360 281408 117366
rect 281356 117302 281408 117308
rect 279804 108990 280016 109018
rect 279804 103494 279832 108990
rect 279792 103488 279844 103494
rect 279792 103430 279844 103436
rect 279700 93900 279752 93906
rect 279700 93842 279752 93848
rect 279712 84182 279740 93842
rect 279700 84176 279752 84182
rect 279700 84118 279752 84124
rect 279792 66292 279844 66298
rect 279792 66234 279844 66240
rect 279804 60738 279832 66234
rect 279804 60722 279924 60738
rect 279804 60716 279936 60722
rect 279804 60710 279884 60716
rect 279884 60658 279936 60664
rect 280068 60716 280120 60722
rect 280068 60658 280120 60664
rect 280080 57934 280108 60658
rect 280068 57928 280120 57934
rect 280068 57870 280120 57876
rect 280068 51060 280120 51066
rect 280068 51002 280120 51008
rect 280080 38690 280108 51002
rect 279884 38684 279936 38690
rect 279884 38626 279936 38632
rect 280068 38684 280120 38690
rect 280068 38626 280120 38632
rect 279896 31754 279924 38626
rect 279884 31748 279936 31754
rect 279884 31690 279936 31696
rect 280068 31748 280120 31754
rect 280068 31690 280120 31696
rect 280080 28966 280108 31690
rect 280068 28960 280120 28966
rect 280068 28902 280120 28908
rect 279976 19372 280028 19378
rect 279976 19314 280028 19320
rect 279988 12458 280016 19314
rect 280356 14498 280384 117302
rect 280356 14470 280476 14498
rect 279988 12430 280108 12458
rect 280080 4146 280108 12430
rect 280448 9722 280476 14470
rect 280436 9716 280488 9722
rect 280436 9658 280488 9664
rect 281264 9716 281316 9722
rect 281264 9658 281316 9664
rect 280068 4140 280120 4146
rect 280068 4082 280120 4088
rect 279160 3998 280108 4026
rect 280080 480 280108 3998
rect 281276 480 281304 9658
rect 281368 3194 281396 117302
rect 281460 3262 281488 120006
rect 282104 117434 282132 120006
rect 282748 117502 282776 120006
rect 283012 117564 283064 117570
rect 283012 117506 283064 117512
rect 282736 117496 282788 117502
rect 282736 117438 282788 117444
rect 282092 117428 282144 117434
rect 282092 117370 282144 117376
rect 283024 14498 283052 117506
rect 283392 117366 283420 120006
rect 283944 118182 283972 120006
rect 283932 118176 283984 118182
rect 283932 118118 283984 118124
rect 284588 118114 284616 120006
rect 284576 118108 284628 118114
rect 284576 118050 284628 118056
rect 284944 117496 284996 117502
rect 284944 117438 284996 117444
rect 283564 117428 283616 117434
rect 283564 117370 283616 117376
rect 283380 117360 283432 117366
rect 283380 117302 283432 117308
rect 282932 14470 283052 14498
rect 282932 9722 282960 14470
rect 282920 9716 282972 9722
rect 282920 9658 282972 9664
rect 283380 9716 283432 9722
rect 283380 9658 283432 9664
rect 282460 4140 282512 4146
rect 282460 4082 282512 4088
rect 281448 3256 281500 3262
rect 281448 3198 281500 3204
rect 281356 3188 281408 3194
rect 281356 3130 281408 3136
rect 282472 480 282500 4082
rect 283392 3890 283420 9658
rect 283576 4078 283604 117370
rect 284208 117360 284260 117366
rect 284208 117302 284260 117308
rect 283564 4072 283616 4078
rect 283564 4014 283616 4020
rect 283392 3862 283696 3890
rect 283668 480 283696 3862
rect 284220 3670 284248 117302
rect 284956 4146 284984 117438
rect 285232 117366 285260 120006
rect 285462 119762 285490 120020
rect 286120 120006 286456 120034
rect 286764 120006 286916 120034
rect 287316 120006 287652 120034
rect 287960 120006 288296 120034
rect 288604 120006 288940 120034
rect 289156 120006 289492 120034
rect 289800 120006 290044 120034
rect 290444 120006 290780 120034
rect 285462 119734 285536 119762
rect 285220 117360 285272 117366
rect 285220 117302 285272 117308
rect 284944 4140 284996 4146
rect 284944 4082 284996 4088
rect 284208 3664 284260 3670
rect 284208 3606 284260 3612
rect 285508 3466 285536 119734
rect 286428 117366 286456 120006
rect 285588 117360 285640 117366
rect 285588 117302 285640 117308
rect 286416 117360 286468 117366
rect 286416 117302 286468 117308
rect 285600 3942 285628 117302
rect 285588 3936 285640 3942
rect 285588 3878 285640 3884
rect 286888 3738 286916 120006
rect 287624 117366 287652 120006
rect 286968 117360 287020 117366
rect 286968 117302 287020 117308
rect 287612 117360 287664 117366
rect 287612 117302 287664 117308
rect 286980 3874 287008 117302
rect 288268 8378 288296 120006
rect 288912 117910 288940 120006
rect 288900 117904 288952 117910
rect 288900 117846 288952 117852
rect 289464 117434 289492 120006
rect 289452 117428 289504 117434
rect 289452 117370 289504 117376
rect 290016 117366 290044 120006
rect 290096 118176 290148 118182
rect 290096 118118 290148 118124
rect 288348 117360 288400 117366
rect 288348 117302 288400 117308
rect 290004 117360 290056 117366
rect 290004 117302 290056 117308
rect 288084 8350 288296 8378
rect 287152 4072 287204 4078
rect 287152 4014 287204 4020
rect 286968 3868 287020 3874
rect 286968 3810 287020 3816
rect 286876 3732 286928 3738
rect 286876 3674 286928 3680
rect 285496 3460 285548 3466
rect 285496 3402 285548 3408
rect 285956 3256 286008 3262
rect 285956 3198 286008 3204
rect 284760 3188 284812 3194
rect 284760 3130 284812 3136
rect 284772 480 284800 3130
rect 285968 480 285996 3198
rect 287164 480 287192 4014
rect 288084 3806 288112 8350
rect 288360 8242 288388 117302
rect 288268 8214 288388 8242
rect 288268 3942 288296 8214
rect 288348 4140 288400 4146
rect 288348 4082 288400 4088
rect 288256 3936 288308 3942
rect 288256 3878 288308 3884
rect 288072 3800 288124 3806
rect 288072 3742 288124 3748
rect 288360 480 288388 4082
rect 289544 3664 289596 3670
rect 289544 3606 289596 3612
rect 289556 480 289584 3606
rect 290108 610 290136 118118
rect 290752 116634 290780 120006
rect 290982 119762 291010 120020
rect 291640 120006 291976 120034
rect 292284 120006 292436 120034
rect 292836 120006 293172 120034
rect 293480 120006 293816 120034
rect 294032 120006 294368 120034
rect 294676 120006 295012 120034
rect 295320 120006 295656 120034
rect 295872 120006 296208 120034
rect 296516 120006 296668 120034
rect 297160 120006 297496 120034
rect 297712 120006 297956 120034
rect 298356 120006 298692 120034
rect 299000 120006 299428 120034
rect 299552 120006 299888 120034
rect 300196 120006 300532 120034
rect 300840 120006 301176 120034
rect 290982 119734 291056 119762
rect 290752 116606 290964 116634
rect 290936 113098 290964 116606
rect 290844 113070 290964 113098
rect 290844 109018 290872 113070
rect 290660 108990 290872 109018
rect 290660 99521 290688 108990
rect 290646 99512 290702 99521
rect 290646 99447 290702 99456
rect 290554 96656 290610 96665
rect 290554 96591 290556 96600
rect 290608 96591 290610 96600
rect 290556 96562 290608 96568
rect 290556 89412 290608 89418
rect 290556 89354 290608 89360
rect 290568 86970 290596 89354
rect 290556 86964 290608 86970
rect 290556 86906 290608 86912
rect 290556 79960 290608 79966
rect 290556 79902 290608 79908
rect 290568 67697 290596 79902
rect 290554 67688 290610 67697
rect 290554 67623 290610 67632
rect 290462 66328 290518 66337
rect 290462 66263 290518 66272
rect 290476 64870 290504 66263
rect 290464 64864 290516 64870
rect 290464 64806 290516 64812
rect 290556 55276 290608 55282
rect 290556 55218 290608 55224
rect 290568 51202 290596 55218
rect 290556 51196 290608 51202
rect 290556 51138 290608 51144
rect 290372 47048 290424 47054
rect 290372 46990 290424 46996
rect 290384 46918 290412 46990
rect 290372 46912 290424 46918
rect 290372 46854 290424 46860
rect 290648 38548 290700 38554
rect 290648 38490 290700 38496
rect 290660 31822 290688 38490
rect 290648 31816 290700 31822
rect 290648 31758 290700 31764
rect 290648 31680 290700 31686
rect 290648 31622 290700 31628
rect 290660 22114 290688 31622
rect 290660 22098 290780 22114
rect 290660 22092 290792 22098
rect 290660 22086 290740 22092
rect 290740 22034 290792 22040
rect 290924 22092 290976 22098
rect 290924 22034 290976 22040
rect 290936 19310 290964 22034
rect 290924 19304 290976 19310
rect 290924 19246 290976 19252
rect 290924 9716 290976 9722
rect 290924 9658 290976 9664
rect 290936 3670 290964 9658
rect 290924 3664 290976 3670
rect 290924 3606 290976 3612
rect 291028 3534 291056 119734
rect 291384 118108 291436 118114
rect 291384 118050 291436 118056
rect 291108 117360 291160 117366
rect 291108 117302 291160 117308
rect 291120 3602 291148 117302
rect 291108 3596 291160 3602
rect 291108 3538 291160 3544
rect 291016 3528 291068 3534
rect 291016 3470 291068 3476
rect 291396 610 291424 118050
rect 291948 117366 291976 120006
rect 291936 117360 291988 117366
rect 291936 117302 291988 117308
rect 292408 4146 292436 120006
rect 293144 117910 293172 120006
rect 293788 118250 293816 120006
rect 293776 118244 293828 118250
rect 293776 118186 293828 118192
rect 294340 117978 294368 120006
rect 294328 117972 294380 117978
rect 294328 117914 294380 117920
rect 293132 117904 293184 117910
rect 293132 117846 293184 117852
rect 293868 117904 293920 117910
rect 293868 117846 293920 117852
rect 292488 117360 292540 117366
rect 292488 117302 292540 117308
rect 292396 4140 292448 4146
rect 292396 4082 292448 4088
rect 292500 3330 292528 117302
rect 293132 4004 293184 4010
rect 293132 3946 293184 3952
rect 292488 3324 292540 3330
rect 292488 3266 292540 3272
rect 290096 604 290148 610
rect 290096 546 290148 552
rect 290740 604 290792 610
rect 290740 546 290792 552
rect 291384 604 291436 610
rect 291384 546 291436 552
rect 291936 604 291988 610
rect 291936 546 291988 552
rect 290752 480 290780 546
rect 291948 480 291976 546
rect 293144 480 293172 3946
rect 293880 3398 293908 117846
rect 294984 117638 295012 120006
rect 295628 118182 295656 120006
rect 296180 118318 296208 120006
rect 296168 118312 296220 118318
rect 296168 118254 296220 118260
rect 295616 118176 295668 118182
rect 295616 118118 295668 118124
rect 296640 118114 296668 120006
rect 296628 118108 296680 118114
rect 296628 118050 296680 118056
rect 297468 117978 297496 120006
rect 295248 117972 295300 117978
rect 295248 117914 295300 117920
rect 297456 117972 297508 117978
rect 297456 117914 297508 117920
rect 294972 117632 295024 117638
rect 294972 117574 295024 117580
rect 294604 117428 294656 117434
rect 294604 117370 294656 117376
rect 294328 3460 294380 3466
rect 294328 3402 294380 3408
rect 293868 3392 293920 3398
rect 293868 3334 293920 3340
rect 294340 480 294368 3402
rect 294616 3262 294644 117370
rect 295260 3466 295288 117914
rect 297364 117836 297416 117842
rect 297364 117778 297416 117784
rect 295524 3868 295576 3874
rect 295524 3810 295576 3816
rect 295248 3460 295300 3466
rect 295248 3402 295300 3408
rect 294604 3256 294656 3262
rect 294604 3198 294656 3204
rect 295536 480 295564 3810
rect 296720 3732 296772 3738
rect 296720 3674 296772 3680
rect 296732 480 296760 3674
rect 297376 3194 297404 117778
rect 297928 4078 297956 120006
rect 298664 118046 298692 120006
rect 298652 118040 298704 118046
rect 298652 117982 298704 117988
rect 298008 117972 298060 117978
rect 298008 117914 298060 117920
rect 298020 4078 298048 117914
rect 297916 4072 297968 4078
rect 297916 4014 297968 4020
rect 298008 4072 298060 4078
rect 298008 4014 298060 4020
rect 297916 3936 297968 3942
rect 297916 3878 297968 3884
rect 297364 3188 297416 3194
rect 297364 3130 297416 3136
rect 297928 480 297956 3878
rect 299400 3874 299428 120006
rect 299860 117570 299888 120006
rect 300504 117978 300532 120006
rect 300492 117972 300544 117978
rect 300492 117914 300544 117920
rect 299848 117564 299900 117570
rect 299848 117506 299900 117512
rect 301148 117366 301176 120006
rect 301378 119762 301406 120020
rect 302036 120006 302188 120034
rect 302680 120006 303016 120034
rect 303232 120006 303476 120034
rect 303876 120006 304212 120034
rect 304520 120006 304856 120034
rect 305072 120006 305408 120034
rect 305716 120006 306052 120034
rect 306360 120006 306696 120034
rect 306912 120006 307248 120034
rect 307556 120006 307708 120034
rect 308200 120006 308536 120034
rect 308752 120006 309088 120034
rect 309396 120006 309732 120034
rect 310040 120006 310468 120034
rect 310592 120006 310928 120034
rect 311236 120006 311572 120034
rect 301378 119734 301452 119762
rect 301136 117360 301188 117366
rect 301136 117302 301188 117308
rect 301424 116113 301452 119734
rect 302160 117774 302188 120006
rect 302884 118244 302936 118250
rect 302884 118186 302936 118192
rect 302148 117768 302200 117774
rect 302148 117710 302200 117716
rect 302148 117360 302200 117366
rect 302148 117302 302200 117308
rect 301410 116104 301466 116113
rect 301410 116039 301466 116048
rect 301778 115968 301834 115977
rect 301700 115938 301778 115954
rect 301688 115932 301778 115938
rect 301740 115926 301778 115932
rect 301778 115903 301834 115912
rect 301964 115932 302016 115938
rect 301688 115874 301740 115880
rect 301964 115874 302016 115880
rect 301700 115843 301728 115874
rect 301976 106282 302004 115874
rect 301964 106276 302016 106282
rect 301964 106218 302016 106224
rect 301964 99340 302016 99346
rect 301964 99282 302016 99288
rect 301976 96642 302004 99282
rect 301976 96614 302096 96642
rect 302068 89706 302096 96614
rect 301884 89678 302096 89706
rect 301884 77382 301912 89678
rect 301872 77376 301924 77382
rect 301872 77318 301924 77324
rect 302056 77376 302108 77382
rect 302056 77318 302108 77324
rect 302068 77178 302096 77318
rect 302056 77172 302108 77178
rect 302056 77114 302108 77120
rect 301964 67652 302016 67658
rect 301964 67594 302016 67600
rect 301976 60738 302004 67594
rect 301792 60710 302004 60738
rect 301792 57934 301820 60710
rect 301780 57928 301832 57934
rect 301780 57870 301832 57876
rect 301872 48340 301924 48346
rect 301872 48282 301924 48288
rect 301884 41426 301912 48282
rect 301884 41398 302004 41426
rect 301976 31890 302004 41398
rect 301964 31884 302016 31890
rect 301964 31826 302016 31832
rect 302056 31748 302108 31754
rect 302056 31690 302108 31696
rect 302068 26353 302096 31690
rect 301870 26344 301926 26353
rect 301870 26279 301926 26288
rect 302054 26344 302110 26353
rect 302054 26279 302110 26288
rect 301884 26246 301912 26279
rect 301872 26240 301924 26246
rect 301872 26182 301924 26188
rect 302056 8356 302108 8362
rect 302056 8298 302108 8304
rect 299388 3868 299440 3874
rect 299388 3810 299440 3816
rect 302068 3806 302096 8298
rect 302160 3942 302188 117302
rect 302148 3936 302200 3942
rect 302148 3878 302200 3884
rect 299112 3800 299164 3806
rect 299112 3742 299164 3748
rect 302056 3800 302108 3806
rect 302056 3742 302108 3748
rect 299124 480 299152 3742
rect 302608 3596 302660 3602
rect 302608 3538 302660 3544
rect 301412 3256 301464 3262
rect 301412 3198 301464 3204
rect 300308 3188 300360 3194
rect 300308 3130 300360 3136
rect 300320 480 300348 3130
rect 301424 480 301452 3198
rect 302620 480 302648 3538
rect 302896 3194 302924 118186
rect 302988 117366 303016 120006
rect 302976 117360 303028 117366
rect 302976 117302 303028 117308
rect 303448 3602 303476 120006
rect 304184 117706 304212 120006
rect 304828 117910 304856 120006
rect 304816 117904 304868 117910
rect 304816 117846 304868 117852
rect 304172 117700 304224 117706
rect 304172 117642 304224 117648
rect 305380 117366 305408 120006
rect 306024 118658 306052 120006
rect 306012 118652 306064 118658
rect 306012 118594 306064 118600
rect 305644 118312 305696 118318
rect 305644 118254 305696 118260
rect 303528 117360 303580 117366
rect 303528 117302 303580 117308
rect 305368 117360 305420 117366
rect 305368 117302 305420 117308
rect 303540 3738 303568 117302
rect 303528 3732 303580 3738
rect 303528 3674 303580 3680
rect 303804 3664 303856 3670
rect 303804 3606 303856 3612
rect 303436 3596 303488 3602
rect 303436 3538 303488 3544
rect 302884 3188 302936 3194
rect 302884 3130 302936 3136
rect 303816 480 303844 3606
rect 305656 3534 305684 118254
rect 306668 117842 306696 120006
rect 307220 118318 307248 120006
rect 307208 118312 307260 118318
rect 307208 118254 307260 118260
rect 307680 118250 307708 120006
rect 308508 118590 308536 120006
rect 308496 118584 308548 118590
rect 308496 118526 308548 118532
rect 307668 118244 307720 118250
rect 307668 118186 307720 118192
rect 308404 118176 308456 118182
rect 308404 118118 308456 118124
rect 306656 117836 306708 117842
rect 306656 117778 306708 117784
rect 306288 117360 306340 117366
rect 306288 117302 306340 117308
rect 306300 3670 306328 117302
rect 307392 4140 307444 4146
rect 307392 4082 307444 4088
rect 306288 3664 306340 3670
rect 306288 3606 306340 3612
rect 305000 3528 305052 3534
rect 305000 3470 305052 3476
rect 305644 3528 305696 3534
rect 305644 3470 305696 3476
rect 306288 3528 306340 3534
rect 306288 3470 306340 3476
rect 305012 480 305040 3470
rect 306300 3330 306328 3470
rect 306196 3324 306248 3330
rect 306196 3266 306248 3272
rect 306288 3324 306340 3330
rect 306288 3266 306340 3272
rect 306208 480 306236 3266
rect 307404 480 307432 4082
rect 308416 2990 308444 118118
rect 309060 3534 309088 120006
rect 309704 118454 309732 120006
rect 309692 118448 309744 118454
rect 309692 118390 309744 118396
rect 310440 4962 310468 120006
rect 310900 118522 310928 120006
rect 310888 118516 310940 118522
rect 310888 118458 310940 118464
rect 311544 118386 311572 120006
rect 311774 119762 311802 120020
rect 312432 120006 312768 120034
rect 311728 119734 311802 119762
rect 311532 118380 311584 118386
rect 311532 118322 311584 118328
rect 311728 118182 311756 119734
rect 311716 118176 311768 118182
rect 311716 118118 311768 118124
rect 311900 117632 311952 117638
rect 311900 117574 311952 117580
rect 310428 4956 310480 4962
rect 310428 4898 310480 4904
rect 309048 3528 309100 3534
rect 309048 3470 309100 3476
rect 310980 3460 311032 3466
rect 310980 3402 311032 3408
rect 308588 3392 308640 3398
rect 308588 3334 308640 3340
rect 308404 2984 308456 2990
rect 308404 2926 308456 2932
rect 308600 480 308628 3334
rect 309784 3188 309836 3194
rect 309784 3130 309836 3136
rect 309796 480 309824 3130
rect 310992 480 311020 3402
rect 311912 626 311940 117574
rect 312740 117366 312768 120006
rect 313062 119762 313090 120020
rect 313628 120006 313964 120034
rect 314272 120006 314608 120034
rect 314916 120006 315252 120034
rect 315468 120006 315988 120034
rect 316112 120006 316448 120034
rect 316756 120006 317184 120034
rect 313062 119734 313136 119762
rect 312728 117360 312780 117366
rect 312728 117302 312780 117308
rect 313108 4826 313136 119734
rect 313936 117366 313964 120006
rect 314580 117638 314608 120006
rect 314844 118108 314896 118114
rect 314844 118050 314896 118056
rect 314568 117632 314620 117638
rect 314568 117574 314620 117580
rect 313188 117360 313240 117366
rect 313188 117302 313240 117308
rect 313924 117360 313976 117366
rect 313924 117302 313976 117308
rect 314568 117360 314620 117366
rect 314568 117302 314620 117308
rect 313096 4820 313148 4826
rect 313096 4762 313148 4768
rect 313200 3466 313228 117302
rect 314580 4894 314608 117302
rect 314568 4888 314620 4894
rect 314568 4830 314620 4836
rect 313188 3460 313240 3466
rect 313188 3402 313240 3408
rect 314856 3346 314884 118050
rect 315224 117366 315252 120006
rect 315304 117564 315356 117570
rect 315304 117506 315356 117512
rect 315212 117360 315264 117366
rect 315212 117302 315264 117308
rect 315316 4146 315344 117506
rect 315856 117360 315908 117366
rect 315856 117302 315908 117308
rect 315868 5914 315896 117302
rect 315960 5982 315988 120006
rect 316420 117366 316448 120006
rect 316408 117360 316460 117366
rect 316408 117302 316460 117308
rect 317156 6050 317184 120006
rect 317294 119762 317322 120020
rect 317952 120006 318288 120034
rect 318596 120006 318748 120034
rect 319148 120006 319484 120034
rect 319792 120006 320128 120034
rect 320436 120006 320772 120034
rect 320988 120006 321508 120034
rect 321632 120006 321968 120034
rect 322276 120006 322428 120034
rect 317248 119734 317322 119762
rect 317248 6866 317276 119734
rect 318260 117434 318288 120006
rect 318248 117428 318300 117434
rect 318248 117370 318300 117376
rect 317328 117360 317380 117366
rect 317328 117302 317380 117308
rect 317236 6860 317288 6866
rect 317236 6802 317288 6808
rect 317144 6044 317196 6050
rect 317144 5986 317196 5992
rect 315948 5976 316000 5982
rect 315948 5918 316000 5924
rect 315856 5908 315908 5914
rect 315856 5850 315908 5856
rect 315304 4140 315356 4146
rect 315304 4082 315356 4088
rect 315856 4140 315908 4146
rect 315856 4082 315908 4088
rect 314568 3324 314620 3330
rect 314856 3318 315804 3346
rect 314568 3266 314620 3272
rect 313372 2984 313424 2990
rect 313372 2926 313424 2932
rect 311912 598 312216 626
rect 312188 480 312216 598
rect 313384 480 313412 2926
rect 314580 480 314608 3266
rect 315776 480 315804 3318
rect 315868 3262 315896 4082
rect 316960 4072 317012 4078
rect 316960 4014 317012 4020
rect 315856 3256 315908 3262
rect 315856 3198 315908 3204
rect 316972 480 317000 4014
rect 317340 3330 317368 117302
rect 318720 6118 318748 120006
rect 318984 118040 319036 118046
rect 318984 117982 319036 117988
rect 318708 6112 318760 6118
rect 318708 6054 318760 6060
rect 318064 4004 318116 4010
rect 318064 3946 318116 3952
rect 317328 3324 317380 3330
rect 317328 3266 317380 3272
rect 318076 480 318104 3946
rect 318996 610 319024 117982
rect 319456 117366 319484 120006
rect 320100 117502 320128 120006
rect 320088 117496 320140 117502
rect 320088 117438 320140 117444
rect 320744 117366 320772 120006
rect 320824 117632 320876 117638
rect 320824 117574 320876 117580
rect 319444 117360 319496 117366
rect 319444 117302 319496 117308
rect 320088 117360 320140 117366
rect 320088 117302 320140 117308
rect 320732 117360 320784 117366
rect 320732 117302 320784 117308
rect 320100 3398 320128 117302
rect 320456 3868 320508 3874
rect 320456 3810 320508 3816
rect 320088 3392 320140 3398
rect 320088 3334 320140 3340
rect 318984 604 319036 610
rect 318984 546 319036 552
rect 319260 604 319312 610
rect 319260 546 319312 552
rect 319272 480 319300 546
rect 320468 480 320496 3810
rect 320836 3194 320864 117574
rect 321376 117360 321428 117366
rect 321376 117302 321428 117308
rect 321388 4214 321416 117302
rect 321376 4208 321428 4214
rect 321376 4150 321428 4156
rect 321480 4146 321508 120006
rect 321940 118046 321968 120006
rect 321928 118040 321980 118046
rect 321928 117982 321980 117988
rect 321744 117972 321796 117978
rect 321744 117914 321796 117920
rect 321756 12442 321784 117914
rect 322204 117428 322256 117434
rect 322204 117370 322256 117376
rect 321744 12436 321796 12442
rect 321744 12378 321796 12384
rect 321468 4140 321520 4146
rect 321468 4082 321520 4088
rect 322216 3262 322244 117370
rect 322400 116006 322428 120006
rect 322814 119762 322842 120020
rect 323472 120006 323808 120034
rect 322814 119734 322888 119762
rect 322388 116000 322440 116006
rect 322388 115942 322440 115948
rect 322572 116000 322624 116006
rect 322572 115942 322624 115948
rect 322584 109018 322612 115942
rect 322584 108990 322704 109018
rect 322676 106282 322704 108990
rect 322664 106276 322716 106282
rect 322664 106218 322716 106224
rect 322664 99340 322716 99346
rect 322664 99282 322716 99288
rect 322676 96642 322704 99282
rect 322676 96614 322796 96642
rect 322768 89758 322796 96614
rect 322572 89752 322624 89758
rect 322756 89752 322808 89758
rect 322624 89700 322704 89706
rect 322572 89694 322704 89700
rect 322756 89694 322808 89700
rect 322584 89678 322704 89694
rect 322676 86970 322704 89678
rect 322664 86964 322716 86970
rect 322664 86906 322716 86912
rect 322756 77308 322808 77314
rect 322756 77250 322808 77256
rect 322768 66298 322796 77250
rect 322664 66292 322716 66298
rect 322664 66234 322716 66240
rect 322756 66292 322808 66298
rect 322756 66234 322808 66240
rect 322676 60738 322704 66234
rect 322676 60710 322796 60738
rect 322768 57934 322796 60710
rect 322756 57928 322808 57934
rect 322756 57870 322808 57876
rect 322664 48340 322716 48346
rect 322664 48282 322716 48288
rect 322676 41426 322704 48282
rect 322676 41398 322796 41426
rect 322768 38622 322796 41398
rect 322756 38616 322808 38622
rect 322756 38558 322808 38564
rect 322664 29028 322716 29034
rect 322664 28970 322716 28976
rect 322676 22114 322704 28970
rect 322676 22086 322796 22114
rect 322768 12458 322796 22086
rect 322584 12430 322796 12458
rect 322584 4282 322612 12430
rect 322756 12368 322808 12374
rect 322756 12310 322808 12316
rect 322572 4276 322624 4282
rect 322572 4218 322624 4224
rect 322768 3890 322796 12310
rect 322860 4010 322888 119734
rect 323780 117366 323808 120006
rect 324102 119762 324130 120020
rect 324668 120006 325004 120034
rect 325312 120006 325464 120034
rect 325956 120006 326292 120034
rect 326508 120006 326936 120034
rect 327152 120006 327488 120034
rect 327796 120006 328132 120034
rect 324102 119734 324176 119762
rect 323768 117360 323820 117366
rect 323768 117302 323820 117308
rect 324148 4350 324176 119734
rect 324976 117502 325004 120006
rect 325436 117978 325464 120006
rect 325424 117972 325476 117978
rect 325424 117914 325476 117920
rect 324964 117496 325016 117502
rect 324964 117438 325016 117444
rect 326264 117366 326292 120006
rect 326344 117496 326396 117502
rect 326344 117438 326396 117444
rect 324228 117360 324280 117366
rect 324228 117302 324280 117308
rect 326252 117360 326304 117366
rect 326252 117302 326304 117308
rect 324136 4344 324188 4350
rect 324136 4286 324188 4292
rect 324240 4078 324268 117302
rect 325700 114572 325752 114578
rect 325700 114514 325752 114520
rect 325712 104854 325740 114514
rect 325700 104848 325752 104854
rect 325700 104790 325752 104796
rect 325700 95260 325752 95266
rect 325700 95202 325752 95208
rect 325712 85542 325740 95202
rect 325700 85536 325752 85542
rect 325700 85478 325752 85484
rect 325700 75948 325752 75954
rect 325700 75890 325752 75896
rect 325712 66230 325740 75890
rect 325700 66224 325752 66230
rect 325700 66166 325752 66172
rect 325516 56636 325568 56642
rect 325516 56578 325568 56584
rect 325528 48385 325556 56578
rect 325514 48376 325570 48385
rect 325514 48311 325570 48320
rect 325698 48376 325754 48385
rect 325698 48311 325754 48320
rect 325712 46918 325740 48311
rect 325700 46912 325752 46918
rect 325700 46854 325752 46860
rect 325700 29096 325752 29102
rect 325700 29038 325752 29044
rect 325712 27606 325740 29038
rect 325700 27600 325752 27606
rect 325700 27542 325752 27548
rect 326252 9716 326304 9722
rect 326252 9658 326304 9664
rect 326264 9602 326292 9658
rect 326172 9574 326292 9602
rect 324228 4072 324280 4078
rect 324228 4014 324280 4020
rect 322848 4004 322900 4010
rect 322848 3946 322900 3952
rect 324044 3936 324096 3942
rect 322768 3862 322888 3890
rect 324044 3878 324096 3884
rect 321652 3256 321704 3262
rect 321652 3198 321704 3204
rect 322204 3256 322256 3262
rect 322204 3198 322256 3204
rect 320824 3188 320876 3194
rect 320824 3130 320876 3136
rect 321664 480 321692 3198
rect 322860 480 322888 3862
rect 324056 480 324084 3878
rect 326172 3806 326200 9574
rect 326356 3942 326384 117438
rect 326908 6798 326936 120006
rect 327460 117366 327488 120006
rect 328104 117502 328132 120006
rect 328196 120006 328348 120034
rect 328992 120006 329328 120034
rect 329544 120006 329788 120034
rect 330188 120006 330524 120034
rect 330832 120006 331168 120034
rect 331384 120006 331720 120034
rect 332028 120006 332456 120034
rect 332672 120006 333008 120034
rect 333224 120006 333560 120034
rect 328092 117496 328144 117502
rect 328092 117438 328144 117444
rect 326988 117360 327040 117366
rect 326988 117302 327040 117308
rect 327448 117360 327500 117366
rect 327448 117302 327500 117308
rect 326896 6792 326948 6798
rect 326896 6734 326948 6740
rect 327000 4418 327028 117302
rect 328196 6730 328224 120006
rect 329300 117774 329328 120006
rect 329288 117768 329340 117774
rect 329288 117710 329340 117716
rect 328276 117496 328328 117502
rect 328276 117438 328328 117444
rect 328184 6724 328236 6730
rect 328184 6666 328236 6672
rect 328288 4486 328316 117438
rect 328368 117360 328420 117366
rect 328368 117302 328420 117308
rect 328276 4480 328328 4486
rect 328276 4422 328328 4428
rect 326988 4412 327040 4418
rect 326988 4354 327040 4360
rect 326344 3936 326396 3942
rect 326344 3878 326396 3884
rect 328380 3874 328408 117302
rect 329760 4554 329788 120006
rect 329840 117700 329892 117706
rect 329840 117642 329892 117648
rect 329748 4548 329800 4554
rect 329748 4490 329800 4496
rect 328368 3868 328420 3874
rect 328368 3810 328420 3816
rect 325240 3800 325292 3806
rect 325240 3742 325292 3748
rect 326160 3800 326212 3806
rect 326160 3742 326212 3748
rect 325252 480 325280 3742
rect 327632 3732 327684 3738
rect 327632 3674 327684 3680
rect 326436 604 326488 610
rect 326436 546 326488 552
rect 326448 480 326476 546
rect 327644 480 327672 3674
rect 328828 3596 328880 3602
rect 328828 3538 328880 3544
rect 328840 480 328868 3538
rect 329852 626 329880 117642
rect 330496 117638 330524 120006
rect 330484 117632 330536 117638
rect 330484 117574 330536 117580
rect 331036 117632 331088 117638
rect 331036 117574 331088 117580
rect 331048 6662 331076 117574
rect 331036 6656 331088 6662
rect 331036 6598 331088 6604
rect 331140 3602 331168 120006
rect 331312 117904 331364 117910
rect 331312 117846 331364 117852
rect 331128 3596 331180 3602
rect 331128 3538 331180 3544
rect 331324 626 331352 117846
rect 331692 117366 331720 120006
rect 331680 117360 331732 117366
rect 331680 117302 331732 117308
rect 332428 6594 332456 120006
rect 332876 118652 332928 118658
rect 332876 118594 332928 118600
rect 332508 117360 332560 117366
rect 332508 117302 332560 117308
rect 332416 6588 332468 6594
rect 332416 6530 332468 6536
rect 332520 4622 332548 117302
rect 332508 4616 332560 4622
rect 332508 4558 332560 4564
rect 332416 3664 332468 3670
rect 332416 3606 332468 3612
rect 329852 598 330064 626
rect 330036 480 330064 598
rect 331232 598 331352 626
rect 331232 480 331260 598
rect 332428 480 332456 3606
rect 332888 610 332916 118594
rect 332980 117434 333008 120006
rect 332968 117428 333020 117434
rect 332968 117370 333020 117376
rect 333532 117366 333560 120006
rect 333716 120006 333868 120034
rect 334512 120006 334848 120034
rect 335064 120006 335216 120034
rect 335708 120006 336044 120034
rect 336352 120006 336688 120034
rect 336904 120006 337240 120034
rect 337548 120006 337976 120034
rect 338192 120006 338528 120034
rect 338744 120006 339080 120034
rect 333520 117360 333572 117366
rect 333520 117302 333572 117308
rect 333716 6458 333744 120006
rect 334624 118312 334676 118318
rect 334624 118254 334676 118260
rect 333980 117836 334032 117842
rect 333980 117778 334032 117784
rect 333888 117428 333940 117434
rect 333888 117370 333940 117376
rect 333796 117360 333848 117366
rect 333796 117302 333848 117308
rect 333704 6452 333756 6458
rect 333704 6394 333756 6400
rect 333808 4690 333836 117302
rect 333796 4684 333848 4690
rect 333796 4626 333848 4632
rect 333900 3738 333928 117370
rect 333888 3732 333940 3738
rect 333888 3674 333940 3680
rect 333992 3346 334020 117778
rect 334636 3806 334664 118254
rect 334820 117366 334848 120006
rect 334808 117360 334860 117366
rect 334808 117302 334860 117308
rect 335188 5506 335216 120006
rect 336016 117366 336044 120006
rect 336660 118318 336688 120006
rect 336648 118312 336700 118318
rect 336648 118254 336700 118260
rect 336924 118244 336976 118250
rect 336924 118186 336976 118192
rect 335268 117360 335320 117366
rect 335268 117302 335320 117308
rect 336004 117360 336056 117366
rect 336004 117302 336056 117308
rect 336648 117360 336700 117366
rect 336648 117302 336700 117308
rect 335176 5500 335228 5506
rect 335176 5442 335228 5448
rect 334624 3800 334676 3806
rect 334624 3742 334676 3748
rect 335280 3670 335308 117302
rect 336660 6526 336688 117302
rect 336648 6520 336700 6526
rect 336648 6462 336700 6468
rect 335912 3800 335964 3806
rect 335912 3742 335964 3748
rect 335268 3664 335320 3670
rect 335268 3606 335320 3612
rect 333992 3318 334756 3346
rect 332876 604 332928 610
rect 332876 546 332928 552
rect 333612 604 333664 610
rect 333612 546 333664 552
rect 333624 480 333652 546
rect 334728 480 334756 3318
rect 335924 480 335952 3742
rect 336936 610 336964 118186
rect 337212 117366 337240 120006
rect 337200 117360 337252 117366
rect 337200 117302 337252 117308
rect 337948 6390 337976 120006
rect 338396 118584 338448 118590
rect 338396 118526 338448 118532
rect 338028 117360 338080 117366
rect 338028 117302 338080 117308
rect 337936 6384 337988 6390
rect 337936 6326 337988 6332
rect 338040 4758 338068 117302
rect 338028 4752 338080 4758
rect 338028 4694 338080 4700
rect 338408 626 338436 118526
rect 338500 118250 338528 120006
rect 338488 118244 338540 118250
rect 338488 118186 338540 118192
rect 339052 117366 339080 120006
rect 339374 119762 339402 120020
rect 340032 120006 340368 120034
rect 340584 120006 340736 120034
rect 341228 120006 341564 120034
rect 341872 120006 342208 120034
rect 342424 120006 342760 120034
rect 343068 120006 343496 120034
rect 343712 120006 344048 120034
rect 344264 120006 344600 120034
rect 339328 119734 339402 119762
rect 339040 117360 339092 117366
rect 339040 117302 339092 117308
rect 339328 6254 339356 119734
rect 339592 118448 339644 118454
rect 339592 118390 339644 118396
rect 339408 117360 339460 117366
rect 339408 117302 339460 117308
rect 339316 6248 339368 6254
rect 339316 6190 339368 6196
rect 339420 5438 339448 117302
rect 339408 5432 339460 5438
rect 339408 5374 339460 5380
rect 339500 3528 339552 3534
rect 339500 3470 339552 3476
rect 336924 604 336976 610
rect 336924 546 336976 552
rect 337108 604 337160 610
rect 337108 546 337160 552
rect 338316 598 338436 626
rect 337120 480 337148 546
rect 338316 480 338344 598
rect 339512 480 339540 3470
rect 339604 3346 339632 118390
rect 340340 117366 340368 120006
rect 340328 117360 340380 117366
rect 340328 117302 340380 117308
rect 340708 5370 340736 120006
rect 341432 118516 341484 118522
rect 341432 118458 341484 118464
rect 340788 117360 340840 117366
rect 340788 117302 340840 117308
rect 340696 5364 340748 5370
rect 340696 5306 340748 5312
rect 339604 3318 340736 3346
rect 340708 480 340736 3318
rect 340800 2854 340828 117302
rect 341444 117178 341472 118458
rect 341536 117366 341564 120006
rect 342180 118454 342208 120006
rect 342168 118448 342220 118454
rect 342168 118390 342220 118396
rect 342732 117366 342760 120006
rect 341524 117360 341576 117366
rect 341524 117302 341576 117308
rect 342168 117360 342220 117366
rect 342168 117302 342220 117308
rect 342720 117360 342772 117366
rect 342720 117302 342772 117308
rect 341444 117150 341564 117178
rect 341536 109018 341564 117150
rect 341444 108990 341564 109018
rect 341444 99521 341472 108990
rect 341430 99512 341486 99521
rect 341430 99447 341486 99456
rect 341338 96656 341394 96665
rect 341064 96620 341116 96626
rect 341338 96591 341340 96600
rect 341064 96562 341116 96568
rect 341392 96591 341394 96600
rect 341340 96562 341392 96568
rect 341076 87009 341104 96562
rect 341062 87000 341118 87009
rect 341062 86935 341118 86944
rect 341246 87000 341302 87009
rect 341246 86935 341302 86944
rect 341260 79914 341288 86935
rect 341260 79886 341380 79914
rect 341352 77178 341380 79886
rect 341340 77172 341392 77178
rect 341340 77114 341392 77120
rect 341432 67652 341484 67658
rect 341432 67594 341484 67600
rect 341444 60738 341472 67594
rect 341444 60710 341564 60738
rect 341536 51202 341564 60710
rect 341524 51196 341576 51202
rect 341524 51138 341576 51144
rect 341524 45620 341576 45626
rect 341524 45562 341576 45568
rect 341536 45490 341564 45562
rect 341524 45484 341576 45490
rect 341524 45426 341576 45432
rect 341432 38276 341484 38282
rect 341432 38218 341484 38224
rect 341444 31686 341472 38218
rect 341432 31680 341484 31686
rect 341432 31622 341484 31628
rect 341524 31680 341576 31686
rect 341524 31622 341576 31628
rect 341536 12458 341564 31622
rect 341536 12430 341656 12458
rect 341628 3602 341656 12430
rect 342180 6322 342208 117302
rect 342168 6316 342220 6322
rect 342168 6258 342220 6264
rect 343468 6186 343496 120006
rect 343916 118380 343968 118386
rect 343916 118322 343968 118328
rect 343548 117360 343600 117366
rect 343548 117302 343600 117308
rect 343456 6180 343508 6186
rect 343456 6122 343508 6128
rect 343560 5302 343588 117302
rect 343548 5296 343600 5302
rect 343548 5238 343600 5244
rect 341892 4956 341944 4962
rect 341892 4898 341944 4904
rect 341616 3596 341668 3602
rect 341616 3538 341668 3544
rect 340788 2848 340840 2854
rect 340788 2790 340840 2796
rect 341904 480 341932 4898
rect 343088 3596 343140 3602
rect 343088 3538 343140 3544
rect 343100 480 343128 3538
rect 343928 610 343956 118322
rect 344020 117842 344048 120006
rect 344008 117836 344060 117842
rect 344008 117778 344060 117784
rect 344572 117366 344600 120006
rect 344756 120006 344908 120034
rect 345552 120006 345888 120034
rect 346104 120006 346348 120034
rect 346748 120006 347084 120034
rect 347300 120006 347636 120034
rect 347944 120006 348280 120034
rect 348588 120006 349016 120034
rect 349140 120006 349476 120034
rect 349784 120006 350120 120034
rect 344560 117360 344612 117366
rect 344560 117302 344612 117308
rect 344756 7750 344784 120006
rect 345204 118176 345256 118182
rect 345204 118118 345256 118124
rect 344928 117836 344980 117842
rect 344928 117778 344980 117784
rect 344836 117360 344888 117366
rect 344836 117302 344888 117308
rect 344744 7744 344796 7750
rect 344744 7686 344796 7692
rect 344848 5234 344876 117302
rect 344836 5228 344888 5234
rect 344836 5170 344888 5176
rect 344940 3534 344968 117778
rect 344928 3528 344980 3534
rect 344928 3470 344980 3476
rect 345216 626 345244 118118
rect 345860 117842 345888 120006
rect 345848 117836 345900 117842
rect 345848 117778 345900 117784
rect 346320 5166 346348 120006
rect 347056 117366 347084 120006
rect 347608 118522 347636 120006
rect 347596 118516 347648 118522
rect 347596 118458 347648 118464
rect 348252 117366 348280 120006
rect 347044 117360 347096 117366
rect 347044 117302 347096 117308
rect 347688 117360 347740 117366
rect 347688 117302 347740 117308
rect 348240 117360 348292 117366
rect 348240 117302 348292 117308
rect 347700 7682 347728 117302
rect 347688 7676 347740 7682
rect 347688 7618 347740 7624
rect 348988 7614 349016 120006
rect 349448 118182 349476 120006
rect 349436 118176 349488 118182
rect 349436 118118 349488 118124
rect 350092 117366 350120 120006
rect 350414 119762 350442 120020
rect 350980 120006 351316 120034
rect 351624 120006 351776 120034
rect 352268 120006 352604 120034
rect 352820 120006 353156 120034
rect 353464 120006 353800 120034
rect 354108 120006 354536 120034
rect 354660 120006 354996 120034
rect 355304 120006 355640 120034
rect 350368 119734 350442 119762
rect 349068 117360 349120 117366
rect 349068 117302 349120 117308
rect 350080 117360 350132 117366
rect 350080 117302 350132 117308
rect 348976 7608 349028 7614
rect 348976 7550 349028 7556
rect 346308 5160 346360 5166
rect 346308 5102 346360 5108
rect 349080 5098 349108 117302
rect 350368 9178 350396 119734
rect 351288 117366 351316 120006
rect 350448 117360 350500 117366
rect 350448 117302 350500 117308
rect 351276 117360 351328 117366
rect 351276 117302 351328 117308
rect 350356 9172 350408 9178
rect 350356 9114 350408 9120
rect 349068 5092 349120 5098
rect 349068 5034 349120 5040
rect 350460 5030 350488 117302
rect 351368 5908 351420 5914
rect 351368 5850 351420 5856
rect 350448 5024 350500 5030
rect 350448 4966 350500 4972
rect 349068 4888 349120 4894
rect 349068 4830 349120 4836
rect 347872 4820 347924 4826
rect 347872 4762 347924 4768
rect 346676 3460 346728 3466
rect 346676 3402 346728 3408
rect 343916 604 343968 610
rect 343916 546 343968 552
rect 344284 604 344336 610
rect 345216 598 345520 626
rect 344284 546 344336 552
rect 344296 480 344324 546
rect 345492 480 345520 598
rect 346688 480 346716 3402
rect 347884 480 347912 4762
rect 349080 480 349108 4830
rect 350264 3188 350316 3194
rect 350264 3130 350316 3136
rect 350276 480 350304 3130
rect 351380 480 351408 5850
rect 351748 4962 351776 120006
rect 352576 117366 352604 120006
rect 353128 118658 353156 120006
rect 353116 118652 353168 118658
rect 353116 118594 353168 118600
rect 353772 117366 353800 120006
rect 351828 117360 351880 117366
rect 351828 117302 351880 117308
rect 352564 117360 352616 117366
rect 352564 117302 352616 117308
rect 353208 117360 353260 117366
rect 353208 117302 353260 117308
rect 353760 117360 353812 117366
rect 353760 117302 353812 117308
rect 351736 4956 351788 4962
rect 351736 4898 351788 4904
rect 351840 3466 351868 117302
rect 353220 9110 353248 117302
rect 353208 9104 353260 9110
rect 353208 9046 353260 9052
rect 354508 9042 354536 120006
rect 354968 117570 354996 120006
rect 354956 117564 355008 117570
rect 354956 117506 355008 117512
rect 355612 117366 355640 120006
rect 355934 119762 355962 120020
rect 356500 120006 356836 120034
rect 357144 120006 357388 120034
rect 357788 120006 358124 120034
rect 358340 120006 358768 120034
rect 358984 120006 359320 120034
rect 359628 120006 360056 120034
rect 360180 120006 360516 120034
rect 360824 120006 361160 120034
rect 355888 119734 355962 119762
rect 354588 117360 354640 117366
rect 354588 117302 354640 117308
rect 355600 117360 355652 117366
rect 355600 117302 355652 117308
rect 354496 9036 354548 9042
rect 354496 8978 354548 8984
rect 352564 5976 352616 5982
rect 352564 5918 352616 5924
rect 351828 3460 351880 3466
rect 351828 3402 351880 3408
rect 352576 480 352604 5918
rect 354600 4894 354628 117302
rect 355888 8974 355916 119734
rect 356808 117638 356836 120006
rect 356796 117632 356848 117638
rect 356796 117574 356848 117580
rect 355968 117360 356020 117366
rect 355968 117302 356020 117308
rect 355876 8968 355928 8974
rect 355876 8910 355928 8916
rect 354956 6044 355008 6050
rect 354956 5986 355008 5992
rect 354588 4888 354640 4894
rect 354588 4830 354640 4836
rect 353760 3324 353812 3330
rect 353760 3266 353812 3272
rect 353772 480 353800 3266
rect 354968 480 354996 5986
rect 355980 4826 356008 117302
rect 356152 6860 356204 6866
rect 356152 6802 356204 6808
rect 355968 4820 356020 4826
rect 355968 4762 356020 4768
rect 356164 480 356192 6802
rect 357360 4865 357388 120006
rect 357992 118108 358044 118114
rect 357992 118050 358044 118056
rect 358004 117178 358032 118050
rect 358096 117366 358124 120006
rect 358176 117768 358228 117774
rect 358176 117710 358228 117716
rect 358084 117360 358136 117366
rect 358084 117302 358136 117308
rect 358004 117150 358124 117178
rect 357346 4856 357402 4865
rect 357346 4791 357402 4800
rect 358096 4146 358124 117150
rect 358084 4140 358136 4146
rect 358084 4082 358136 4088
rect 358188 3330 358216 117710
rect 358636 117360 358688 117366
rect 358636 117302 358688 117308
rect 358648 8498 358676 117302
rect 358636 8492 358688 8498
rect 358636 8434 358688 8440
rect 358740 7138 358768 120006
rect 359292 117366 359320 120006
rect 359280 117360 359332 117366
rect 359280 117302 359332 117308
rect 360028 8566 360056 120006
rect 360488 117706 360516 120006
rect 360476 117700 360528 117706
rect 360476 117642 360528 117648
rect 361132 117366 361160 120006
rect 361454 119762 361482 120020
rect 362020 120006 362356 120034
rect 362664 120006 362908 120034
rect 363308 120006 363644 120034
rect 363860 120006 364104 120034
rect 364504 120006 364840 120034
rect 365056 120006 365576 120034
rect 365700 120006 366036 120034
rect 366344 120006 366680 120034
rect 361408 119734 361482 119762
rect 360108 117360 360160 117366
rect 360108 117302 360160 117308
rect 361120 117360 361172 117366
rect 361120 117302 361172 117308
rect 360016 8560 360068 8566
rect 360016 8502 360068 8508
rect 360120 7206 360148 117302
rect 361408 8702 361436 119734
rect 362328 118590 362356 120006
rect 362316 118584 362368 118590
rect 362316 118526 362368 118532
rect 361488 117360 361540 117366
rect 361488 117302 361540 117308
rect 361396 8696 361448 8702
rect 361396 8638 361448 8644
rect 361500 7274 361528 117302
rect 362880 7342 362908 120006
rect 363512 118040 363564 118046
rect 363512 117982 363564 117988
rect 363524 117178 363552 117982
rect 363616 117366 363644 120006
rect 364076 117774 364104 120006
rect 364064 117768 364116 117774
rect 364064 117710 364116 117716
rect 364812 117366 364840 120006
rect 363604 117360 363656 117366
rect 363604 117302 363656 117308
rect 364248 117360 364300 117366
rect 364248 117302 364300 117308
rect 364800 117360 364852 117366
rect 364800 117302 364852 117308
rect 363524 117150 363644 117178
rect 362868 7336 362920 7342
rect 362868 7278 362920 7284
rect 361488 7268 361540 7274
rect 361488 7210 361540 7216
rect 360108 7200 360160 7206
rect 360108 7142 360160 7148
rect 358728 7132 358780 7138
rect 358728 7074 358780 7080
rect 358544 6112 358596 6118
rect 358544 6054 358596 6060
rect 358176 3324 358228 3330
rect 358176 3266 358228 3272
rect 357348 3256 357400 3262
rect 357348 3198 357400 3204
rect 357360 480 357388 3198
rect 358556 480 358584 6054
rect 362132 4208 362184 4214
rect 362132 4150 362184 4156
rect 360936 4140 360988 4146
rect 360936 4082 360988 4088
rect 359740 3392 359792 3398
rect 359740 3334 359792 3340
rect 359752 480 359780 3334
rect 360948 480 360976 4082
rect 362144 480 362172 4150
rect 363616 4146 363644 117150
rect 364260 8634 364288 117302
rect 365548 8770 365576 120006
rect 366008 118386 366036 120006
rect 365996 118380 366048 118386
rect 365996 118322 366048 118328
rect 366652 117366 366680 120006
rect 366882 119762 366910 120020
rect 367540 120006 367876 120034
rect 368184 120006 368428 120034
rect 368736 120006 369072 120034
rect 369380 120006 369716 120034
rect 370024 120006 370360 120034
rect 370576 120006 371096 120034
rect 371220 120006 371556 120034
rect 371864 120006 372200 120034
rect 366882 119734 366956 119762
rect 365628 117360 365680 117366
rect 365628 117302 365680 117308
rect 366640 117360 366692 117366
rect 366640 117302 366692 117308
rect 365536 8764 365588 8770
rect 365536 8706 365588 8712
rect 364248 8628 364300 8634
rect 364248 8570 364300 8576
rect 365640 7410 365668 117302
rect 366928 8838 366956 119734
rect 367848 117502 367876 120006
rect 367836 117496 367888 117502
rect 367836 117438 367888 117444
rect 367008 117360 367060 117366
rect 367008 117302 367060 117308
rect 366916 8832 366968 8838
rect 366916 8774 366968 8780
rect 367020 7478 367048 117302
rect 368400 9654 368428 120006
rect 369044 117366 369072 120006
rect 369688 118182 369716 120006
rect 369676 118176 369728 118182
rect 369676 118118 369728 118124
rect 369124 117972 369176 117978
rect 369124 117914 369176 117920
rect 369032 117360 369084 117366
rect 369032 117302 369084 117308
rect 368388 9648 368440 9654
rect 368388 9590 368440 9596
rect 367008 7472 367060 7478
rect 367008 7414 367060 7420
rect 365628 7404 365680 7410
rect 365628 7346 365680 7352
rect 365720 4276 365772 4282
rect 365720 4218 365772 4224
rect 363604 4140 363656 4146
rect 363604 4082 363656 4088
rect 364524 4140 364576 4146
rect 364524 4082 364576 4088
rect 363328 4004 363380 4010
rect 363328 3946 363380 3952
rect 363340 480 363368 3946
rect 364536 480 364564 4082
rect 365732 480 365760 4218
rect 368020 4072 368072 4078
rect 368020 4014 368072 4020
rect 366916 3596 366968 3602
rect 366916 3538 366968 3544
rect 366928 480 366956 3538
rect 368032 480 368060 4014
rect 369136 2990 369164 117914
rect 369216 117564 369268 117570
rect 369216 117506 369268 117512
rect 369228 4842 369256 117506
rect 370332 117366 370360 120006
rect 369768 117360 369820 117366
rect 369768 117302 369820 117308
rect 370320 117360 370372 117366
rect 370320 117302 370372 117308
rect 369780 8906 369808 117302
rect 371068 10742 371096 120006
rect 371528 117434 371556 120006
rect 371516 117428 371568 117434
rect 371516 117370 371568 117376
rect 372172 117366 372200 120006
rect 372402 119762 372430 120020
rect 373060 120006 373396 120034
rect 373704 120006 373948 120034
rect 374256 120006 374592 120034
rect 374900 120006 375328 120034
rect 375544 120006 375880 120034
rect 376096 120006 376616 120034
rect 376740 120006 377076 120034
rect 377384 120006 377720 120034
rect 372356 119734 372430 119762
rect 371148 117360 371200 117366
rect 371148 117302 371200 117308
rect 372160 117360 372212 117366
rect 372160 117302 372212 117308
rect 371056 10736 371108 10742
rect 371056 10678 371108 10684
rect 371160 9586 371188 117302
rect 372356 10674 372384 119734
rect 373368 118114 373396 120006
rect 373356 118108 373408 118114
rect 373356 118050 373408 118056
rect 372528 117428 372580 117434
rect 372528 117370 372580 117376
rect 372436 117360 372488 117366
rect 372436 117302 372488 117308
rect 372344 10668 372396 10674
rect 372344 10610 372396 10616
rect 371148 9580 371200 9586
rect 371148 9522 371200 9528
rect 372448 9518 372476 117302
rect 372436 9512 372488 9518
rect 372436 9454 372488 9460
rect 369768 8900 369820 8906
rect 369768 8842 369820 8848
rect 369228 4814 369440 4842
rect 369216 4344 369268 4350
rect 369216 4286 369268 4292
rect 369124 2984 369176 2990
rect 369124 2926 369176 2932
rect 369228 480 369256 4286
rect 369412 2922 369440 4814
rect 370412 3936 370464 3942
rect 370412 3878 370464 3884
rect 369400 2916 369452 2922
rect 369400 2858 369452 2864
rect 370424 480 370452 3878
rect 372540 3126 372568 117370
rect 373920 5642 373948 120006
rect 374564 117366 374592 120006
rect 374644 118312 374696 118318
rect 374644 118254 374696 118260
rect 374552 117360 374604 117366
rect 374552 117302 374604 117308
rect 374000 6792 374052 6798
rect 374000 6734 374052 6740
rect 373908 5636 373960 5642
rect 373908 5578 373960 5584
rect 372804 4412 372856 4418
rect 372804 4354 372856 4360
rect 372528 3120 372580 3126
rect 372528 3062 372580 3068
rect 371608 2984 371660 2990
rect 371608 2926 371660 2932
rect 371620 480 371648 2926
rect 372816 480 372844 4354
rect 374012 480 374040 6734
rect 374656 3942 374684 118254
rect 375196 117360 375248 117366
rect 375196 117302 375248 117308
rect 375208 10606 375236 117302
rect 375196 10600 375248 10606
rect 375196 10542 375248 10548
rect 374644 3936 374696 3942
rect 374644 3878 374696 3884
rect 375196 3868 375248 3874
rect 375196 3810 375248 3816
rect 375208 480 375236 3810
rect 375300 3194 375328 120006
rect 375852 117366 375880 120006
rect 376024 118516 376076 118522
rect 376024 118458 376076 118464
rect 375840 117360 375892 117366
rect 375840 117302 375892 117308
rect 375288 3188 375340 3194
rect 375288 3130 375340 3136
rect 376036 2990 376064 118458
rect 376588 10538 376616 120006
rect 377048 118318 377076 120006
rect 377036 118312 377088 118318
rect 377036 118254 377088 118260
rect 377404 117496 377456 117502
rect 377404 117438 377456 117444
rect 376668 117360 376720 117366
rect 376668 117302 376720 117308
rect 376576 10532 376628 10538
rect 376576 10474 376628 10480
rect 376680 5574 376708 117302
rect 376668 5568 376720 5574
rect 376668 5510 376720 5516
rect 376392 4480 376444 4486
rect 376392 4422 376444 4428
rect 376024 2984 376076 2990
rect 376024 2926 376076 2932
rect 376404 480 376432 4422
rect 377416 3058 377444 117438
rect 377692 117366 377720 120006
rect 377922 119762 377950 120020
rect 378580 120006 378916 120034
rect 379224 120006 379376 120034
rect 379776 120006 380112 120034
rect 380420 120006 380756 120034
rect 381064 120006 381400 120034
rect 381616 120006 382136 120034
rect 382260 120006 382596 120034
rect 382812 120006 382964 120034
rect 377922 119734 377996 119762
rect 377680 117360 377732 117366
rect 377680 117302 377732 117308
rect 377968 10470 377996 119734
rect 378888 117366 378916 120006
rect 378048 117360 378100 117366
rect 378048 117302 378100 117308
rect 378876 117360 378928 117366
rect 378876 117302 378928 117308
rect 377956 10464 378008 10470
rect 377956 10406 378008 10412
rect 377588 6724 377640 6730
rect 377588 6666 377640 6672
rect 377404 3052 377456 3058
rect 377404 2994 377456 3000
rect 377600 480 377628 6666
rect 378060 5710 378088 117302
rect 379348 5846 379376 120006
rect 380084 117366 380112 120006
rect 380728 117978 380756 120006
rect 380716 117972 380768 117978
rect 380716 117914 380768 117920
rect 381372 117366 381400 120006
rect 379428 117360 379480 117366
rect 379428 117302 379480 117308
rect 380072 117360 380124 117366
rect 380072 117302 380124 117308
rect 380808 117360 380860 117366
rect 380808 117302 380860 117308
rect 381360 117360 381412 117366
rect 381360 117302 381412 117308
rect 379336 5840 379388 5846
rect 379336 5782 379388 5788
rect 378048 5704 378100 5710
rect 378048 5646 378100 5652
rect 378784 3324 378836 3330
rect 378784 3266 378836 3272
rect 378796 480 378824 3266
rect 379440 3262 379468 117302
rect 380820 10402 380848 117302
rect 380808 10396 380860 10402
rect 380808 10338 380860 10344
rect 382108 10334 382136 120006
rect 382568 117366 382596 120006
rect 382188 117360 382240 117366
rect 382188 117302 382240 117308
rect 382556 117360 382608 117366
rect 382556 117302 382608 117308
rect 382096 10328 382148 10334
rect 382096 10270 382148 10276
rect 381176 6656 381228 6662
rect 381176 6598 381228 6604
rect 379980 4548 380032 4554
rect 379980 4490 380032 4496
rect 379428 3256 379480 3262
rect 379428 3198 379480 3204
rect 379992 480 380020 4490
rect 381188 480 381216 6598
rect 382200 5778 382228 117302
rect 382936 116006 382964 120006
rect 383442 119762 383470 120020
rect 384100 120006 384436 120034
rect 384652 120006 384988 120034
rect 385296 120006 385632 120034
rect 385940 120006 386276 120034
rect 386492 120006 386828 120034
rect 387136 120006 387656 120034
rect 387780 120006 388116 120034
rect 383442 119734 383516 119762
rect 382924 116000 382976 116006
rect 382924 115942 382976 115948
rect 383108 116000 383160 116006
rect 383108 115942 383160 115948
rect 383120 109018 383148 115942
rect 383120 108990 383332 109018
rect 383304 99482 383332 108990
rect 383292 99476 383344 99482
rect 383292 99418 383344 99424
rect 383200 99340 383252 99346
rect 383200 99282 383252 99288
rect 383212 96626 383240 99282
rect 383200 96620 383252 96626
rect 383200 96562 383252 96568
rect 383108 87032 383160 87038
rect 383108 86974 383160 86980
rect 383120 79914 383148 86974
rect 383120 79886 383240 79914
rect 383212 77178 383240 79886
rect 383200 77172 383252 77178
rect 383200 77114 383252 77120
rect 383292 67652 383344 67658
rect 383292 67594 383344 67600
rect 383304 60858 383332 67594
rect 383292 60852 383344 60858
rect 383292 60794 383344 60800
rect 383200 60716 383252 60722
rect 383200 60658 383252 60664
rect 383212 57934 383240 60658
rect 383200 57928 383252 57934
rect 383200 57870 383252 57876
rect 383292 48340 383344 48346
rect 383292 48282 383344 48288
rect 383304 43466 383332 48282
rect 383212 43438 383332 43466
rect 383212 38622 383240 43438
rect 383200 38616 383252 38622
rect 383200 38558 383252 38564
rect 383292 29028 383344 29034
rect 383292 28970 383344 28976
rect 383304 28914 383332 28970
rect 383304 28886 383424 28914
rect 383396 25294 383424 28886
rect 383384 25288 383436 25294
rect 383384 25230 383436 25236
rect 383384 19372 383436 19378
rect 383384 19314 383436 19320
rect 383396 19258 383424 19314
rect 383304 19230 383424 19258
rect 383304 12578 383332 19230
rect 383292 12572 383344 12578
rect 383292 12514 383344 12520
rect 383292 9716 383344 9722
rect 383292 9658 383344 9664
rect 383304 7546 383332 9658
rect 383292 7540 383344 7546
rect 383292 7482 383344 7488
rect 383488 5982 383516 119734
rect 384212 118244 384264 118250
rect 384212 118186 384264 118192
rect 384224 118130 384252 118186
rect 384224 118102 384344 118130
rect 383568 117360 383620 117366
rect 383568 117302 383620 117308
rect 383476 5976 383528 5982
rect 383476 5918 383528 5924
rect 383580 5828 383608 117302
rect 383488 5800 383608 5828
rect 382188 5772 382240 5778
rect 382188 5714 382240 5720
rect 382372 3732 382424 3738
rect 382372 3674 382424 3680
rect 382384 480 382412 3674
rect 383488 3330 383516 5800
rect 383568 4616 383620 4622
rect 383568 4558 383620 4564
rect 383476 3324 383528 3330
rect 383476 3266 383528 3272
rect 383580 480 383608 4558
rect 384316 3738 384344 118102
rect 384408 117570 384436 120006
rect 384396 117564 384448 117570
rect 384396 117506 384448 117512
rect 384960 8294 384988 120006
rect 385604 117366 385632 120006
rect 386248 118250 386276 120006
rect 386236 118244 386288 118250
rect 386236 118186 386288 118192
rect 386800 117366 386828 120006
rect 387628 118674 387656 120006
rect 387536 118646 387656 118674
rect 385592 117360 385644 117366
rect 385592 117302 385644 117308
rect 386328 117360 386380 117366
rect 386328 117302 386380 117308
rect 386788 117360 386840 117366
rect 386788 117302 386840 117308
rect 384948 8288 385000 8294
rect 384948 8230 385000 8236
rect 384672 6588 384724 6594
rect 384672 6530 384724 6536
rect 384304 3732 384356 3738
rect 384304 3674 384356 3680
rect 384684 480 384712 6530
rect 386340 5914 386368 117302
rect 387536 109070 387564 118646
rect 388088 117366 388116 120006
rect 388318 119762 388346 120020
rect 388962 119762 388990 120020
rect 389620 120006 389956 120034
rect 390172 120006 390508 120034
rect 390816 120006 391152 120034
rect 391460 120006 391888 120034
rect 392012 120006 392348 120034
rect 392656 120006 393176 120034
rect 393300 120006 393636 120034
rect 388318 119734 388392 119762
rect 388962 119734 389036 119762
rect 387616 117360 387668 117366
rect 387616 117302 387668 117308
rect 388076 117360 388128 117366
rect 388076 117302 388128 117308
rect 387524 109064 387576 109070
rect 387524 109006 387576 109012
rect 387628 8226 387656 117302
rect 388364 116113 388392 119734
rect 388350 116104 388406 116113
rect 388350 116039 388406 116048
rect 388718 115968 388774 115977
rect 388718 115903 388720 115912
rect 388772 115903 388774 115912
rect 388904 115932 388956 115938
rect 388720 115874 388772 115880
rect 388904 115874 388956 115880
rect 387708 109064 387760 109070
rect 387708 109006 387760 109012
rect 387616 8220 387668 8226
rect 387616 8162 387668 8168
rect 387720 6050 387748 109006
rect 388916 106321 388944 115874
rect 388718 106312 388774 106321
rect 388902 106312 388958 106321
rect 388718 106247 388720 106256
rect 388772 106247 388774 106256
rect 388812 106276 388864 106282
rect 388720 106218 388772 106224
rect 388902 106247 388958 106256
rect 388812 106218 388864 106224
rect 388824 96642 388852 106218
rect 388732 96626 388852 96642
rect 388720 96620 388852 96626
rect 388772 96614 388852 96620
rect 388720 96562 388772 96568
rect 388732 96531 388760 96562
rect 388628 87032 388680 87038
rect 388628 86974 388680 86980
rect 388640 82090 388668 86974
rect 388640 82062 388852 82090
rect 388824 79914 388852 82062
rect 388732 79886 388852 79914
rect 388732 77178 388760 79886
rect 388720 77172 388772 77178
rect 388720 77114 388772 77120
rect 388812 67652 388864 67658
rect 388812 67594 388864 67600
rect 388824 60858 388852 67594
rect 388812 60852 388864 60858
rect 388812 60794 388864 60800
rect 388720 60716 388772 60722
rect 388720 60658 388772 60664
rect 388732 57934 388760 60658
rect 388720 57928 388772 57934
rect 388720 57870 388772 57876
rect 388812 48340 388864 48346
rect 388812 48282 388864 48288
rect 388824 43466 388852 48282
rect 388732 43438 388852 43466
rect 388732 31754 388760 43438
rect 388720 31748 388772 31754
rect 388720 31690 388772 31696
rect 388904 31748 388956 31754
rect 388904 31690 388956 31696
rect 388916 24206 388944 31690
rect 388720 24200 388772 24206
rect 388720 24142 388772 24148
rect 388904 24200 388956 24206
rect 388904 24142 388956 24148
rect 388732 12458 388760 24142
rect 388732 12430 388944 12458
rect 388916 8158 388944 12430
rect 388904 8152 388956 8158
rect 388904 8094 388956 8100
rect 388260 6452 388312 6458
rect 388260 6394 388312 6400
rect 387708 6044 387760 6050
rect 387708 5986 387760 5992
rect 386328 5908 386380 5914
rect 386328 5850 386380 5856
rect 387064 4684 387116 4690
rect 387064 4626 387116 4632
rect 385868 3800 385920 3806
rect 385868 3742 385920 3748
rect 385880 480 385908 3742
rect 387076 480 387104 4626
rect 388272 480 388300 6394
rect 389008 6118 389036 119734
rect 389824 118448 389876 118454
rect 389824 118390 389876 118396
rect 389088 117360 389140 117366
rect 389088 117302 389140 117308
rect 388996 6112 389048 6118
rect 388996 6054 389048 6060
rect 389100 3398 389128 117302
rect 389836 3806 389864 118390
rect 389928 118318 389956 120006
rect 389916 118312 389968 118318
rect 389916 118254 389968 118260
rect 390480 8090 390508 120006
rect 391124 117638 391152 120006
rect 391112 117632 391164 117638
rect 391112 117574 391164 117580
rect 391756 117632 391808 117638
rect 391756 117574 391808 117580
rect 390468 8084 390520 8090
rect 390468 8026 390520 8032
rect 391768 6866 391796 117574
rect 391756 6860 391808 6866
rect 391756 6802 391808 6808
rect 391860 6746 391888 120006
rect 392320 117366 392348 120006
rect 393148 118674 393176 120006
rect 393056 118646 393176 118674
rect 392308 117360 392360 117366
rect 392308 117302 392360 117308
rect 393056 109070 393084 118646
rect 393608 118522 393636 120006
rect 393596 118516 393648 118522
rect 393596 118458 393648 118464
rect 393964 117496 394016 117502
rect 393964 117438 394016 117444
rect 393136 117360 393188 117366
rect 393136 117302 393188 117308
rect 393044 109064 393096 109070
rect 393044 109006 393096 109012
rect 393148 8022 393176 117302
rect 393228 109064 393280 109070
rect 393228 109006 393280 109012
rect 393136 8016 393188 8022
rect 393136 7958 393188 7964
rect 393240 6798 393268 109006
rect 391768 6718 391888 6746
rect 393228 6792 393280 6798
rect 393228 6734 393280 6740
rect 390652 5500 390704 5506
rect 390652 5442 390704 5448
rect 389824 3800 389876 3806
rect 389824 3742 389876 3748
rect 389456 3664 389508 3670
rect 389456 3606 389508 3612
rect 389088 3392 389140 3398
rect 389088 3334 389140 3340
rect 389468 480 389496 3606
rect 390664 480 390692 5442
rect 391768 4146 391796 6718
rect 391848 6520 391900 6526
rect 391848 6462 391900 6468
rect 391756 4140 391808 4146
rect 391756 4082 391808 4088
rect 391860 480 391888 6462
rect 393044 3868 393096 3874
rect 393044 3810 393096 3816
rect 393056 480 393084 3810
rect 393976 3670 394004 117438
rect 394160 109018 394188 120278
rect 403696 120142 404124 120170
rect 414736 120142 414888 120170
rect 420164 120142 420408 120170
rect 394496 120006 394648 120034
rect 394160 108990 394372 109018
rect 394344 108882 394372 108990
rect 394344 108854 394464 108882
rect 394436 106282 394464 108854
rect 394424 106276 394476 106282
rect 394424 106218 394476 106224
rect 394424 99340 394476 99346
rect 394424 99282 394476 99288
rect 394436 96642 394464 99282
rect 394436 96614 394556 96642
rect 394528 89758 394556 96614
rect 394332 89752 394384 89758
rect 394516 89752 394568 89758
rect 394384 89700 394464 89706
rect 394332 89694 394464 89700
rect 394516 89694 394568 89700
rect 394344 89678 394464 89694
rect 394436 86970 394464 89678
rect 394424 86964 394476 86970
rect 394424 86906 394476 86912
rect 394516 77308 394568 77314
rect 394516 77250 394568 77256
rect 394528 67658 394556 77250
rect 394424 67652 394476 67658
rect 394424 67594 394476 67600
rect 394516 67652 394568 67658
rect 394516 67594 394568 67600
rect 394436 60738 394464 67594
rect 394436 60710 394556 60738
rect 394528 48346 394556 60710
rect 394424 48340 394476 48346
rect 394424 48282 394476 48288
rect 394516 48340 394568 48346
rect 394516 48282 394568 48288
rect 394436 41426 394464 48282
rect 394436 41398 394556 41426
rect 394528 29034 394556 41398
rect 394424 29028 394476 29034
rect 394424 28970 394476 28976
rect 394516 29028 394568 29034
rect 394516 28970 394568 28976
rect 394436 19394 394464 28970
rect 394344 19366 394464 19394
rect 394344 12510 394372 19366
rect 394332 12504 394384 12510
rect 394332 12446 394384 12452
rect 394424 12368 394476 12374
rect 394424 12310 394476 12316
rect 394436 9602 394464 12310
rect 394344 9574 394464 9602
rect 394344 7954 394372 9574
rect 394332 7948 394384 7954
rect 394332 7890 394384 7896
rect 394620 6730 394648 120006
rect 395126 119814 395154 120020
rect 395692 120006 395936 120034
rect 396336 120006 396672 120034
rect 396980 120006 397316 120034
rect 397532 120006 397868 120034
rect 398176 120006 398696 120034
rect 398820 120006 399156 120034
rect 399372 120006 399708 120034
rect 395114 119808 395166 119814
rect 395114 119750 395166 119756
rect 395908 7886 395936 120006
rect 395988 119808 396040 119814
rect 395988 119750 396040 119756
rect 395896 7880 395948 7886
rect 395896 7822 395948 7828
rect 394608 6724 394660 6730
rect 394608 6666 394660 6672
rect 395436 6384 395488 6390
rect 395436 6326 395488 6332
rect 394240 4752 394292 4758
rect 394240 4694 394292 4700
rect 393964 3664 394016 3670
rect 393964 3606 394016 3612
rect 394252 480 394280 4694
rect 395448 480 395476 6326
rect 396000 4078 396028 119750
rect 396644 117366 396672 120006
rect 397288 118454 397316 120006
rect 397276 118448 397328 118454
rect 397276 118390 397328 118396
rect 396724 117836 396776 117842
rect 396724 117778 396776 117784
rect 396632 117360 396684 117366
rect 396632 117302 396684 117308
rect 395988 4072 396040 4078
rect 395988 4014 396040 4020
rect 396736 3738 396764 117778
rect 397840 117366 397868 120006
rect 398104 117700 398156 117706
rect 398104 117642 398156 117648
rect 397368 117360 397420 117366
rect 397368 117302 397420 117308
rect 397828 117360 397880 117366
rect 397828 117302 397880 117308
rect 397380 6662 397408 117302
rect 397368 6656 397420 6662
rect 397368 6598 397420 6604
rect 397828 5432 397880 5438
rect 397828 5374 397880 5380
rect 396632 3732 396684 3738
rect 396632 3674 396684 3680
rect 396724 3732 396776 3738
rect 396724 3674 396776 3680
rect 396644 480 396672 3674
rect 397840 480 397868 5374
rect 398116 3602 398144 117642
rect 398668 6594 398696 120006
rect 399128 117366 399156 120006
rect 399680 117502 399708 120006
rect 400002 119762 400030 120020
rect 400568 120006 400904 120034
rect 401212 120006 401548 120034
rect 401856 120006 402192 120034
rect 402408 120006 402928 120034
rect 403052 120006 403388 120034
rect 399956 119734 400030 119762
rect 399668 117496 399720 117502
rect 399668 117438 399720 117444
rect 398748 117360 398800 117366
rect 398748 117302 398800 117308
rect 399116 117360 399168 117366
rect 399116 117302 399168 117308
rect 398656 6588 398708 6594
rect 398656 6530 398708 6536
rect 398760 4214 398788 117302
rect 399956 6526 399984 119734
rect 400876 117774 400904 120006
rect 400864 117768 400916 117774
rect 400864 117710 400916 117716
rect 400036 117496 400088 117502
rect 400036 117438 400088 117444
rect 399944 6520 399996 6526
rect 399944 6462 399996 6468
rect 399024 6248 399076 6254
rect 399024 6190 399076 6196
rect 398748 4208 398800 4214
rect 398748 4150 398800 4156
rect 398104 3596 398156 3602
rect 398104 3538 398156 3544
rect 399036 480 399064 6190
rect 400048 4282 400076 117438
rect 400128 117360 400180 117366
rect 400128 117302 400180 117308
rect 400036 4276 400088 4282
rect 400036 4218 400088 4224
rect 400140 4010 400168 117302
rect 401324 5364 401376 5370
rect 401324 5306 401376 5312
rect 400128 4004 400180 4010
rect 400128 3946 400180 3952
rect 400220 2848 400272 2854
rect 400220 2790 400272 2796
rect 400232 480 400260 2790
rect 401336 480 401364 5306
rect 401520 4418 401548 120006
rect 402164 117366 402192 120006
rect 402152 117360 402204 117366
rect 402152 117302 402204 117308
rect 402796 117360 402848 117366
rect 402796 117302 402848 117308
rect 402244 117292 402296 117298
rect 402244 117234 402296 117240
rect 401508 4412 401560 4418
rect 401508 4354 401560 4360
rect 402256 2854 402284 117234
rect 402808 6458 402836 117302
rect 402796 6452 402848 6458
rect 402796 6394 402848 6400
rect 402520 6316 402572 6322
rect 402520 6258 402572 6264
rect 402244 2848 402296 2854
rect 402244 2790 402296 2796
rect 402532 480 402560 6258
rect 402900 3942 402928 120006
rect 403360 117366 403388 120006
rect 403348 117360 403400 117366
rect 403348 117302 403400 117308
rect 404096 115938 404124 120142
rect 404234 119762 404262 120020
rect 404892 120006 405228 120034
rect 404234 119734 404308 119762
rect 404280 117638 404308 119734
rect 404268 117632 404320 117638
rect 404268 117574 404320 117580
rect 405200 117434 405228 120006
rect 405522 119762 405550 120020
rect 406088 120006 406424 120034
rect 406732 120006 406976 120034
rect 407376 120006 407712 120034
rect 407928 120006 408264 120034
rect 408572 120006 408908 120034
rect 409216 120006 409644 120034
rect 405522 119734 405596 119762
rect 405188 117428 405240 117434
rect 405188 117370 405240 117376
rect 404268 117360 404320 117366
rect 404268 117302 404320 117308
rect 404084 115932 404136 115938
rect 404084 115874 404136 115880
rect 403900 106344 403952 106350
rect 403900 106286 403952 106292
rect 403912 99414 403940 106286
rect 403900 99408 403952 99414
rect 403900 99350 403952 99356
rect 403992 99340 404044 99346
rect 403992 99282 404044 99288
rect 404004 96626 404032 99282
rect 403992 96620 404044 96626
rect 403992 96562 404044 96568
rect 403900 87032 403952 87038
rect 403900 86974 403952 86980
rect 403912 79914 403940 86974
rect 403912 79886 404032 79914
rect 404004 77178 404032 79886
rect 403992 77172 404044 77178
rect 403992 77114 404044 77120
rect 404084 67652 404136 67658
rect 404084 67594 404136 67600
rect 404096 60858 404124 67594
rect 404084 60852 404136 60858
rect 404084 60794 404136 60800
rect 403992 60716 404044 60722
rect 403992 60658 404044 60664
rect 404004 57934 404032 60658
rect 403992 57928 404044 57934
rect 403992 57870 404044 57876
rect 404084 48340 404136 48346
rect 404084 48282 404136 48288
rect 404096 43466 404124 48282
rect 404004 43438 404124 43466
rect 404004 38622 404032 43438
rect 403992 38616 404044 38622
rect 403992 38558 404044 38564
rect 404084 29028 404136 29034
rect 404084 28970 404136 28976
rect 404096 22166 404124 28970
rect 404084 22160 404136 22166
rect 404084 22102 404136 22108
rect 403992 22092 404044 22098
rect 403992 22034 404044 22040
rect 404004 12458 404032 22034
rect 404004 12430 404216 12458
rect 404188 6390 404216 12430
rect 404176 6384 404228 6390
rect 404176 6326 404228 6332
rect 404280 4350 404308 117302
rect 405568 6254 405596 119734
rect 405648 117428 405700 117434
rect 405648 117370 405700 117376
rect 405556 6248 405608 6254
rect 405556 6190 405608 6196
rect 404912 5296 404964 5302
rect 404912 5238 404964 5244
rect 404268 4344 404320 4350
rect 404268 4286 404320 4292
rect 402888 3936 402940 3942
rect 402888 3878 402940 3884
rect 403716 3800 403768 3806
rect 403716 3742 403768 3748
rect 403728 480 403756 3742
rect 404924 480 404952 5238
rect 405660 4486 405688 117370
rect 406396 117366 406424 120006
rect 406384 117360 406436 117366
rect 406384 117302 406436 117308
rect 406108 6180 406160 6186
rect 406108 6122 406160 6128
rect 405648 4480 405700 4486
rect 405648 4422 405700 4428
rect 406120 480 406148 6122
rect 406948 4554 406976 120006
rect 407684 117366 407712 120006
rect 408236 117434 408264 120006
rect 408224 117428 408276 117434
rect 408224 117370 408276 117376
rect 408880 117366 408908 120006
rect 407028 117360 407080 117366
rect 407028 117302 407080 117308
rect 407672 117360 407724 117366
rect 407672 117302 407724 117308
rect 408408 117360 408460 117366
rect 408408 117302 408460 117308
rect 408868 117360 408920 117366
rect 408868 117302 408920 117308
rect 406936 4548 406988 4554
rect 406936 4490 406988 4496
rect 407040 3874 407068 117302
rect 408420 6322 408448 117302
rect 409512 9240 409564 9246
rect 409512 9182 409564 9188
rect 408408 6316 408460 6322
rect 408408 6258 408460 6264
rect 408684 5228 408736 5234
rect 408684 5170 408736 5176
rect 407028 3868 407080 3874
rect 407028 3810 407080 3816
rect 408314 3768 408370 3777
rect 408314 3703 408370 3712
rect 408498 3768 408554 3777
rect 408498 3703 408554 3712
rect 408328 3602 408356 3703
rect 408512 3602 408540 3703
rect 408316 3596 408368 3602
rect 408316 3538 408368 3544
rect 408500 3596 408552 3602
rect 408500 3538 408552 3544
rect 407304 3528 407356 3534
rect 408696 3482 408724 5170
rect 409524 3806 409552 9182
rect 409616 6186 409644 120006
rect 409754 119762 409782 120020
rect 410412 120006 410748 120034
rect 409754 119734 409828 119762
rect 409696 117360 409748 117366
rect 409696 117302 409748 117308
rect 409708 8514 409736 117302
rect 409800 9246 409828 119734
rect 410720 117366 410748 120006
rect 411042 119762 411070 120020
rect 411608 120006 411944 120034
rect 412252 120006 412588 120034
rect 412896 120006 413232 120034
rect 413448 120006 413784 120034
rect 414092 120006 414428 120034
rect 411042 119734 411116 119762
rect 410708 117360 410760 117366
rect 410708 117302 410760 117308
rect 409788 9240 409840 9246
rect 409788 9182 409840 9188
rect 409708 8486 409828 8514
rect 409696 7744 409748 7750
rect 409696 7686 409748 7692
rect 409604 6180 409656 6186
rect 409604 6122 409656 6128
rect 409512 3800 409564 3806
rect 409512 3742 409564 3748
rect 407304 3470 407356 3476
rect 407316 480 407344 3470
rect 408512 3454 408724 3482
rect 408512 480 408540 3454
rect 409708 480 409736 7686
rect 409800 4622 409828 8486
rect 411088 6225 411116 119734
rect 411916 117706 411944 120006
rect 411904 117700 411956 117706
rect 411904 117642 411956 117648
rect 411168 117360 411220 117366
rect 411168 117302 411220 117308
rect 411074 6216 411130 6225
rect 411074 6151 411130 6160
rect 411180 4690 411208 117302
rect 412088 5160 412140 5166
rect 412088 5102 412140 5108
rect 411168 4684 411220 4690
rect 411168 4626 411220 4632
rect 409788 4616 409840 4622
rect 409788 4558 409840 4564
rect 410892 3732 410944 3738
rect 410892 3674 410944 3680
rect 410904 480 410932 3674
rect 412100 480 412128 5102
rect 412560 4758 412588 120006
rect 413204 117366 413232 120006
rect 413284 117564 413336 117570
rect 413284 117506 413336 117512
rect 413192 117360 413244 117366
rect 413192 117302 413244 117308
rect 413296 10690 413324 117506
rect 413756 117502 413784 120006
rect 413744 117496 413796 117502
rect 413744 117438 413796 117444
rect 414400 117366 414428 120006
rect 413928 117360 413980 117366
rect 413928 117302 413980 117308
rect 414388 117360 414440 117366
rect 414388 117302 414440 117308
rect 413204 10662 413324 10690
rect 412548 4752 412600 4758
rect 412548 4694 412600 4700
rect 413204 3670 413232 10662
rect 413940 7818 413968 117302
rect 414860 115938 414888 120142
rect 415274 119762 415302 120020
rect 415932 120006 416268 120034
rect 415274 119734 415348 119762
rect 415320 117774 415348 119734
rect 415308 117768 415360 117774
rect 415308 117710 415360 117716
rect 416044 117496 416096 117502
rect 416044 117438 416096 117444
rect 415308 117360 415360 117366
rect 415308 117302 415360 117308
rect 414848 115932 414900 115938
rect 414848 115874 414900 115880
rect 414940 115932 414992 115938
rect 414940 115874 414992 115880
rect 414952 108882 414980 115874
rect 414952 108854 415072 108882
rect 415044 104854 415072 108854
rect 415032 104848 415084 104854
rect 415032 104790 415084 104796
rect 415216 95260 415268 95266
rect 415216 95202 415268 95208
rect 415228 89826 415256 95202
rect 415216 89820 415268 89826
rect 415216 89762 415268 89768
rect 415124 89684 415176 89690
rect 415124 89626 415176 89632
rect 415136 75954 415164 89626
rect 415032 75948 415084 75954
rect 415032 75890 415084 75896
rect 415124 75948 415176 75954
rect 415124 75890 415176 75896
rect 415044 66230 415072 75890
rect 415032 66224 415084 66230
rect 415032 66166 415084 66172
rect 415032 56636 415084 56642
rect 415032 56578 415084 56584
rect 415044 51338 415072 56578
rect 415032 51332 415084 51338
rect 415032 51274 415084 51280
rect 415216 51332 415268 51338
rect 415216 51274 415268 51280
rect 415228 48385 415256 51274
rect 415030 48376 415086 48385
rect 414952 48334 415030 48362
rect 414952 45558 414980 48334
rect 415030 48311 415086 48320
rect 415214 48376 415270 48385
rect 415214 48311 415270 48320
rect 414940 45552 414992 45558
rect 414940 45494 414992 45500
rect 415032 35964 415084 35970
rect 415032 35906 415084 35912
rect 415044 26246 415072 35906
rect 415032 26240 415084 26246
rect 415032 26182 415084 26188
rect 415032 16652 415084 16658
rect 415032 16594 415084 16600
rect 415044 12510 415072 16594
rect 415032 12504 415084 12510
rect 415032 12446 415084 12452
rect 414940 12436 414992 12442
rect 414940 12378 414992 12384
rect 413928 7812 413980 7818
rect 413928 7754 413980 7760
rect 414952 7750 414980 12378
rect 414940 7744 414992 7750
rect 414940 7686 414992 7692
rect 413284 7676 413336 7682
rect 413284 7618 413336 7624
rect 413192 3664 413244 3670
rect 413192 3606 413244 3612
rect 413296 480 413324 7618
rect 415320 5506 415348 117302
rect 415308 5500 415360 5506
rect 415308 5442 415360 5448
rect 415676 5092 415728 5098
rect 415676 5034 415728 5040
rect 414480 2984 414532 2990
rect 414480 2926 414532 2932
rect 414492 480 414520 2926
rect 415688 480 415716 5034
rect 416056 2990 416084 117438
rect 416240 117366 416268 120006
rect 416562 119762 416590 120020
rect 417128 120006 417464 120034
rect 417772 120006 418108 120034
rect 418324 120006 418660 120034
rect 418968 120006 419304 120034
rect 419612 120006 419948 120034
rect 416562 119734 416636 119762
rect 416228 117360 416280 117366
rect 416228 117302 416280 117308
rect 416608 7682 416636 119734
rect 416780 117904 416832 117910
rect 416780 117846 416832 117852
rect 416688 117360 416740 117366
rect 416688 117302 416740 117308
rect 416596 7676 416648 7682
rect 416596 7618 416648 7624
rect 416700 5438 416728 117302
rect 416792 7614 416820 117846
rect 417436 117706 417464 120006
rect 417424 117700 417476 117706
rect 417424 117642 417476 117648
rect 416780 7608 416832 7614
rect 416780 7550 416832 7556
rect 417976 7608 418028 7614
rect 417976 7550 418028 7556
rect 416872 7064 416924 7070
rect 416872 7006 416924 7012
rect 416688 5432 416740 5438
rect 416688 5374 416740 5380
rect 416044 2984 416096 2990
rect 416044 2926 416096 2932
rect 416884 480 416912 7006
rect 417882 3632 417938 3641
rect 417882 3567 417938 3576
rect 417896 3534 417924 3567
rect 417884 3528 417936 3534
rect 417884 3470 417936 3476
rect 417988 480 418016 7550
rect 418080 5370 418108 120006
rect 418160 117768 418212 117774
rect 418158 117736 418160 117745
rect 418212 117736 418214 117745
rect 418158 117671 418214 117680
rect 418632 117502 418660 120006
rect 419276 117570 419304 120006
rect 419264 117564 419316 117570
rect 419264 117506 419316 117512
rect 419920 117502 419948 120006
rect 420380 117994 420408 120142
rect 420794 119762 420822 120020
rect 421452 120006 421788 120034
rect 422004 120006 422156 120034
rect 422648 120006 422984 120034
rect 423292 120006 423628 120034
rect 423844 120006 424180 120034
rect 424488 120006 424824 120034
rect 425132 120006 425468 120034
rect 420794 119734 420868 119762
rect 420380 117966 420592 117994
rect 420184 117564 420236 117570
rect 420184 117506 420236 117512
rect 418620 117496 418672 117502
rect 418620 117438 418672 117444
rect 419448 117496 419500 117502
rect 419448 117438 419500 117444
rect 419908 117496 419960 117502
rect 419908 117438 419960 117444
rect 419460 9450 419488 117438
rect 419448 9444 419500 9450
rect 419448 9386 419500 9392
rect 418068 5364 418120 5370
rect 418068 5306 418120 5312
rect 419172 5024 419224 5030
rect 419172 4966 419224 4972
rect 418160 3732 418212 3738
rect 418160 3674 418212 3680
rect 418172 2990 418200 3674
rect 418342 3632 418398 3641
rect 418342 3567 418398 3576
rect 418356 3466 418384 3567
rect 418344 3460 418396 3466
rect 418344 3402 418396 3408
rect 418160 2984 418212 2990
rect 418160 2926 418212 2932
rect 419184 480 419212 4966
rect 420196 3670 420224 117506
rect 420564 115938 420592 117966
rect 420840 117910 420868 119734
rect 420828 117904 420880 117910
rect 420828 117846 420880 117852
rect 421760 117502 421788 120006
rect 420828 117496 420880 117502
rect 420828 117438 420880 117444
rect 421748 117496 421800 117502
rect 421748 117438 421800 117444
rect 420552 115932 420604 115938
rect 420552 115874 420604 115880
rect 420552 108996 420604 109002
rect 420552 108938 420604 108944
rect 420564 106298 420592 108938
rect 420564 106282 420684 106298
rect 420552 106276 420696 106282
rect 420604 106270 420644 106276
rect 420552 106218 420604 106224
rect 420644 106218 420696 106224
rect 420564 99362 420592 106218
rect 420564 99334 420684 99362
rect 420656 96642 420684 99334
rect 420656 96626 420776 96642
rect 420656 96620 420788 96626
rect 420656 96614 420736 96620
rect 420736 96562 420788 96568
rect 420748 96531 420776 96562
rect 420644 87032 420696 87038
rect 420644 86974 420696 86980
rect 420656 82142 420684 86974
rect 420276 82136 420328 82142
rect 420276 82078 420328 82084
rect 420644 82136 420696 82142
rect 420644 82078 420696 82084
rect 420288 77353 420316 82078
rect 420274 77344 420330 77353
rect 420274 77279 420330 77288
rect 420458 77344 420514 77353
rect 420514 77302 420592 77330
rect 420458 77279 420514 77288
rect 420564 66298 420592 77302
rect 420460 66292 420512 66298
rect 420460 66234 420512 66240
rect 420552 66292 420604 66298
rect 420552 66234 420604 66240
rect 420472 66162 420500 66234
rect 420460 66156 420512 66162
rect 420460 66098 420512 66104
rect 420644 66156 420696 66162
rect 420644 66098 420696 66104
rect 420656 61441 420684 66098
rect 420642 61432 420698 61441
rect 420642 61367 420698 61376
rect 420550 48376 420606 48385
rect 420472 48334 420550 48362
rect 420472 46918 420500 48334
rect 420550 48311 420606 48320
rect 420460 46912 420512 46918
rect 420460 46854 420512 46860
rect 420644 46912 420696 46918
rect 420644 46854 420696 46860
rect 420656 42129 420684 46854
rect 420642 42120 420698 42129
rect 420642 42055 420698 42064
rect 420550 29064 420606 29073
rect 420472 29022 420550 29050
rect 420472 27606 420500 29022
rect 420550 28999 420606 29008
rect 420460 27600 420512 27606
rect 420460 27542 420512 27548
rect 420552 18012 420604 18018
rect 420552 17954 420604 17960
rect 420564 12510 420592 17954
rect 420552 12504 420604 12510
rect 420552 12446 420604 12452
rect 420460 12436 420512 12442
rect 420460 12378 420512 12384
rect 420472 9382 420500 12378
rect 420460 9376 420512 9382
rect 420460 9318 420512 9324
rect 420368 9172 420420 9178
rect 420368 9114 420420 9120
rect 420184 3664 420236 3670
rect 420184 3606 420236 3612
rect 420380 480 420408 9114
rect 420840 5302 420868 117438
rect 422128 9314 422156 120006
rect 422956 117706 422984 120006
rect 422944 117700 422996 117706
rect 422944 117642 422996 117648
rect 422208 117496 422260 117502
rect 422208 117438 422260 117444
rect 422116 9308 422168 9314
rect 422116 9250 422168 9256
rect 420828 5296 420880 5302
rect 420828 5238 420880 5244
rect 422220 5234 422248 117438
rect 422208 5228 422260 5234
rect 422208 5170 422260 5176
rect 423600 5098 423628 120006
rect 424152 117502 424180 120006
rect 424796 118726 424824 120006
rect 424784 118720 424836 118726
rect 424784 118662 424836 118668
rect 425336 118652 425388 118658
rect 425336 118594 425388 118600
rect 424324 117700 424376 117706
rect 424324 117642 424376 117648
rect 424140 117496 424192 117502
rect 424140 117438 424192 117444
rect 423956 9104 424008 9110
rect 423956 9046 424008 9052
rect 423588 5092 423640 5098
rect 423588 5034 423640 5040
rect 422760 4956 422812 4962
rect 422760 4898 422812 4904
rect 421564 3528 421616 3534
rect 421564 3470 421616 3476
rect 421576 480 421604 3470
rect 422772 480 422800 4898
rect 423968 480 423996 9046
rect 424336 2990 424364 117642
rect 424968 117496 425020 117502
rect 424968 117438 425020 117444
rect 424980 9246 425008 117438
rect 424968 9240 425020 9246
rect 424968 9182 425020 9188
rect 424324 2984 424376 2990
rect 424324 2926 424376 2932
rect 425348 610 425376 118594
rect 425440 117502 425468 120006
rect 425428 117496 425480 117502
rect 425428 117438 425480 117444
rect 426084 115938 426112 120278
rect 426314 119762 426342 120020
rect 426972 120006 427308 120034
rect 427524 120006 427676 120034
rect 428168 120006 428504 120034
rect 428812 120006 429148 120034
rect 429364 120006 429700 120034
rect 430008 120006 430344 120034
rect 430652 120006 430988 120034
rect 431204 120006 431540 120034
rect 426314 119734 426388 119762
rect 426360 118658 426388 119734
rect 426348 118652 426400 118658
rect 426348 118594 426400 118600
rect 427280 117502 427308 120006
rect 426348 117496 426400 117502
rect 426348 117438 426400 117444
rect 427268 117496 427320 117502
rect 427268 117438 427320 117444
rect 426072 115932 426124 115938
rect 426072 115874 426124 115880
rect 426256 115932 426308 115938
rect 426256 115874 426308 115880
rect 426268 104854 426296 115874
rect 426256 104848 426308 104854
rect 426256 104790 426308 104796
rect 426256 95328 426308 95334
rect 426256 95270 426308 95276
rect 426268 87038 426296 95270
rect 426256 87032 426308 87038
rect 426256 86974 426308 86980
rect 426164 85604 426216 85610
rect 426164 85546 426216 85552
rect 426176 84182 426204 85546
rect 426164 84176 426216 84182
rect 426164 84118 426216 84124
rect 426072 69692 426124 69698
rect 426072 69634 426124 69640
rect 426084 53174 426112 69634
rect 426072 53168 426124 53174
rect 426072 53110 426124 53116
rect 426256 53168 426308 53174
rect 426256 53110 426308 53116
rect 426268 48385 426296 53110
rect 426070 48376 426126 48385
rect 425992 48334 426070 48362
rect 425992 46918 426020 48334
rect 426070 48311 426126 48320
rect 426254 48376 426310 48385
rect 426254 48311 426310 48320
rect 425980 46912 426032 46918
rect 425980 46854 426032 46860
rect 426072 37324 426124 37330
rect 426072 37266 426124 37272
rect 426084 19310 426112 37266
rect 425980 19304 426032 19310
rect 425980 19246 426032 19252
rect 426072 19304 426124 19310
rect 426072 19246 426124 19252
rect 425992 9178 426020 19246
rect 425980 9172 426032 9178
rect 425980 9114 426032 9120
rect 426360 5166 426388 117438
rect 427648 9110 427676 120006
rect 427726 117736 427782 117745
rect 427726 117671 427728 117680
rect 427780 117671 427782 117680
rect 427728 117642 427780 117648
rect 428476 117502 428504 120006
rect 427728 117496 427780 117502
rect 427728 117438 427780 117444
rect 428464 117496 428516 117502
rect 428464 117438 428516 117444
rect 427636 9104 427688 9110
rect 427636 9046 427688 9052
rect 427544 9036 427596 9042
rect 427544 8978 427596 8984
rect 426348 5160 426400 5166
rect 426348 5102 426400 5108
rect 426348 4888 426400 4894
rect 426348 4830 426400 4836
rect 425152 604 425204 610
rect 425152 546 425204 552
rect 425336 604 425388 610
rect 425336 546 425388 552
rect 425164 480 425192 546
rect 426360 480 426388 4830
rect 427556 480 427584 8978
rect 427740 5030 427768 117438
rect 427728 5024 427780 5030
rect 427728 4966 427780 4972
rect 429120 4962 429148 120006
rect 429672 117774 429700 120006
rect 429844 118652 429896 118658
rect 429844 118594 429896 118600
rect 429660 117768 429712 117774
rect 429660 117710 429712 117716
rect 429108 4956 429160 4962
rect 429108 4898 429160 4904
rect 427634 3632 427690 3641
rect 427634 3567 427636 3576
rect 427688 3567 427690 3576
rect 427818 3632 427874 3641
rect 427818 3567 427874 3576
rect 427636 3538 427688 3544
rect 427832 3534 427860 3567
rect 427820 3528 427872 3534
rect 427820 3470 427872 3476
rect 429856 2922 429884 118594
rect 430316 117502 430344 120006
rect 430960 117774 430988 120006
rect 430488 117768 430540 117774
rect 430488 117710 430540 117716
rect 430948 117768 431000 117774
rect 430948 117710 431000 117716
rect 430304 117496 430356 117502
rect 430304 117438 430356 117444
rect 430500 7614 430528 117710
rect 431224 117496 431276 117502
rect 431224 117438 431276 117444
rect 431132 8968 431184 8974
rect 431132 8910 431184 8916
rect 430488 7608 430540 7614
rect 430488 7550 430540 7556
rect 429936 4820 429988 4826
rect 429936 4762 429988 4768
rect 428740 2916 428792 2922
rect 428740 2858 428792 2864
rect 429844 2916 429896 2922
rect 429844 2858 429896 2864
rect 428752 480 428780 2858
rect 429948 480 429976 4762
rect 431144 480 431172 8910
rect 431236 3369 431264 117438
rect 431512 115938 431540 120006
rect 431834 119762 431862 120020
rect 432492 120006 432828 120034
rect 433044 120006 433196 120034
rect 433688 120006 434024 120034
rect 431788 119734 431862 119762
rect 431788 118658 431816 119734
rect 431776 118652 431828 118658
rect 431776 118594 431828 118600
rect 431868 117768 431920 117774
rect 431868 117710 431920 117716
rect 431500 115932 431552 115938
rect 431500 115874 431552 115880
rect 431684 108996 431736 109002
rect 431684 108938 431736 108944
rect 431696 106282 431724 108938
rect 431592 106276 431644 106282
rect 431592 106218 431644 106224
rect 431684 106276 431736 106282
rect 431684 106218 431736 106224
rect 431604 104854 431632 106218
rect 431592 104848 431644 104854
rect 431592 104790 431644 104796
rect 431592 87032 431644 87038
rect 431592 86974 431644 86980
rect 431604 80102 431632 86974
rect 431788 80102 431816 80133
rect 431592 80096 431644 80102
rect 431776 80096 431828 80102
rect 431644 80044 431776 80050
rect 431592 80038 431828 80044
rect 431604 80022 431816 80038
rect 431604 75886 431632 80022
rect 431592 75880 431644 75886
rect 431592 75822 431644 75828
rect 431592 66292 431644 66298
rect 431592 66234 431644 66240
rect 431604 56574 431632 66234
rect 431592 56568 431644 56574
rect 431592 56510 431644 56516
rect 431776 56568 431828 56574
rect 431776 56510 431828 56516
rect 431788 47025 431816 56510
rect 431590 47016 431646 47025
rect 431590 46951 431646 46960
rect 431774 47016 431830 47025
rect 431774 46951 431830 46960
rect 431604 46918 431632 46951
rect 431500 46912 431552 46918
rect 431500 46854 431552 46860
rect 431592 46912 431644 46918
rect 431592 46854 431644 46860
rect 431512 37346 431540 46854
rect 431512 37318 431632 37346
rect 431604 37262 431632 37318
rect 431592 37256 431644 37262
rect 431592 37198 431644 37204
rect 431684 31680 431736 31686
rect 431684 31622 431736 31628
rect 431696 26246 431724 31622
rect 431684 26240 431736 26246
rect 431684 26182 431736 26188
rect 431500 16652 431552 16658
rect 431500 16594 431552 16600
rect 431512 9042 431540 16594
rect 431500 9036 431552 9042
rect 431500 8978 431552 8984
rect 431880 4894 431908 117710
rect 432800 117502 432828 120006
rect 432788 117496 432840 117502
rect 432788 117438 432840 117444
rect 433168 8974 433196 120006
rect 433996 118017 434024 120006
rect 433982 118008 434038 118017
rect 433982 117943 434038 117952
rect 433248 117496 433300 117502
rect 433248 117438 433300 117444
rect 433156 8968 433208 8974
rect 433156 8910 433208 8916
rect 431868 4888 431920 4894
rect 431868 4830 431920 4836
rect 433260 4826 433288 117438
rect 435008 80034 435036 196143
rect 435100 188873 435128 251194
rect 435180 207052 435232 207058
rect 435180 206994 435232 207000
rect 435192 190233 435220 206994
rect 435178 190224 435234 190233
rect 435178 190159 435234 190168
rect 435086 188864 435142 188873
rect 435086 188799 435142 188808
rect 436112 180305 436140 385630
rect 436560 201136 436612 201142
rect 436560 201078 436612 201084
rect 436468 201068 436520 201074
rect 436468 201010 436520 201016
rect 436376 201000 436428 201006
rect 436376 200942 436428 200948
rect 436190 198928 436246 198937
rect 436190 198863 436246 198872
rect 436098 180296 436154 180305
rect 436098 180231 436154 180240
rect 436100 155236 436152 155242
rect 436100 155178 436152 155184
rect 436112 155145 436140 155178
rect 436098 155136 436154 155145
rect 436098 155071 436154 155080
rect 436100 149048 436152 149054
rect 436100 148990 436152 148996
rect 436112 148753 436140 148990
rect 436098 148744 436154 148753
rect 436098 148679 436154 148688
rect 436100 142112 436152 142118
rect 436098 142080 436100 142089
rect 436152 142080 436154 142089
rect 436098 142015 436154 142024
rect 434996 80028 435048 80034
rect 434996 79970 435048 79976
rect 436204 35902 436232 198863
rect 436282 194032 436338 194041
rect 436282 193967 436338 193976
rect 436296 120630 436324 193967
rect 436388 176225 436416 200942
rect 436480 177993 436508 201010
rect 436572 182073 436600 201078
rect 436652 200184 436704 200190
rect 436652 200126 436704 200132
rect 436664 193089 436692 200126
rect 436650 193080 436706 193089
rect 436650 193015 436706 193024
rect 436558 182064 436614 182073
rect 436558 181999 436614 182008
rect 436466 177984 436522 177993
rect 436466 177919 436522 177928
rect 436374 176216 436430 176225
rect 436374 176151 436430 176160
rect 436756 140457 436784 438874
rect 436836 157412 436888 157418
rect 436836 157354 436888 157360
rect 436742 140448 436798 140457
rect 436742 140383 436798 140392
rect 436848 127809 436876 157354
rect 438136 155242 438164 700402
rect 462332 700398 462360 703520
rect 478524 700505 478552 703520
rect 478510 700496 478566 700505
rect 494808 700466 494836 703520
rect 478510 700431 478566 700440
rect 494796 700460 494848 700466
rect 494796 700402 494848 700408
rect 462320 700392 462372 700398
rect 462320 700334 462372 700340
rect 447784 700324 447836 700330
rect 447784 700266 447836 700272
rect 446404 673532 446456 673538
rect 446404 673474 446456 673480
rect 445024 626612 445076 626618
rect 445024 626554 445076 626560
rect 442264 579692 442316 579698
rect 442264 579634 442316 579640
rect 438216 485852 438268 485858
rect 438216 485794 438268 485800
rect 438124 155236 438176 155242
rect 438124 155178 438176 155184
rect 437388 153196 437440 153202
rect 437388 153138 437440 153144
rect 437400 152833 437428 153138
rect 437386 152824 437442 152833
rect 437386 152759 437442 152768
rect 437388 150408 437440 150414
rect 437388 150350 437440 150356
rect 437400 150249 437428 150350
rect 437386 150240 437442 150249
rect 437386 150175 437442 150184
rect 437386 146296 437442 146305
rect 437386 146231 437442 146240
rect 437400 146198 437428 146231
rect 437388 146192 437440 146198
rect 437388 146134 437440 146140
rect 437020 144900 437072 144906
rect 437020 144842 437072 144848
rect 437032 144537 437060 144842
rect 437018 144528 437074 144537
rect 437018 144463 437074 144472
rect 438228 142118 438256 485794
rect 442276 146198 442304 579634
rect 445036 149054 445064 626554
rect 446416 150414 446444 673474
rect 447796 153202 447824 700266
rect 511264 556300 511316 556306
rect 511264 556242 511316 556248
rect 484400 556232 484452 556238
rect 484400 556174 484452 556180
rect 484412 554676 484440 556174
rect 511276 554676 511304 556242
rect 514024 532772 514076 532778
rect 514024 532714 514076 532720
rect 478892 520118 480010 520146
rect 506492 520118 506874 520146
rect 464252 389428 464304 389434
rect 464252 389370 464304 389376
rect 464264 387532 464292 389370
rect 475844 389360 475896 389366
rect 475844 389302 475896 389308
rect 475856 387532 475884 389302
rect 478892 387122 478920 520118
rect 487436 389292 487488 389298
rect 487436 389234 487488 389240
rect 487448 387532 487476 389234
rect 499028 389224 499080 389230
rect 499028 389166 499080 389172
rect 499040 387532 499068 389166
rect 478880 387116 478932 387122
rect 478880 387058 478932 387064
rect 504730 378448 504786 378457
rect 503732 378406 504730 378434
rect 456798 375184 456854 375193
rect 456798 375119 456854 375128
rect 456812 374066 456840 375119
rect 456800 374060 456852 374066
rect 456800 374002 456852 374008
rect 503732 361434 503760 378406
rect 504730 378383 504786 378392
rect 503640 361406 503760 361434
rect 503640 360074 503668 361406
rect 504730 360496 504786 360505
rect 504376 360454 504730 360482
rect 503640 360046 503760 360074
rect 503732 359938 503760 360046
rect 503732 359910 503852 359938
rect 457442 358048 457498 358057
rect 457442 357983 457498 357992
rect 457456 202502 457484 357983
rect 503824 350554 503852 359910
rect 504376 351914 504404 360454
rect 504730 360431 504786 360440
rect 504100 351886 504404 351914
rect 504100 350554 504128 351886
rect 503824 350526 504036 350554
rect 504100 350526 504220 350554
rect 504008 344978 504036 350526
rect 503916 344950 504036 344978
rect 503812 342032 503864 342038
rect 503812 341974 503864 341980
rect 503718 340912 503774 340921
rect 503718 340847 503774 340856
rect 460584 337618 460612 340068
rect 460572 337612 460624 337618
rect 460572 337554 460624 337560
rect 472176 337550 472204 340068
rect 472164 337544 472216 337550
rect 472164 337486 472216 337492
rect 483768 337482 483796 340068
rect 483756 337476 483808 337482
rect 483756 337418 483808 337424
rect 495360 337414 495388 340068
rect 495348 337408 495400 337414
rect 495348 337350 495400 337356
rect 503732 331378 503760 340847
rect 503640 331350 503760 331378
rect 503640 331226 503668 331350
rect 503824 331294 503852 341974
rect 503916 340921 503944 344950
rect 504192 342038 504220 350526
rect 504824 345092 504876 345098
rect 504824 345034 504876 345040
rect 504730 343632 504786 343641
rect 504730 343567 504786 343576
rect 504180 342032 504232 342038
rect 504180 341974 504232 341980
rect 503902 340912 503958 340921
rect 504744 340882 504772 343567
rect 503902 340847 503958 340856
rect 504732 340876 504784 340882
rect 504732 340818 504784 340824
rect 503904 340808 503956 340814
rect 503904 340750 503956 340756
rect 503812 331288 503864 331294
rect 503812 331230 503864 331236
rect 503628 331220 503680 331226
rect 503628 331162 503680 331168
rect 503720 328568 503772 328574
rect 503720 328510 503772 328516
rect 503732 321706 503760 328510
rect 503916 321774 503944 340750
rect 503996 331220 504048 331226
rect 503996 331162 504048 331168
rect 503904 321768 503956 321774
rect 503904 321710 503956 321716
rect 504008 321706 504036 331162
rect 504836 328681 504864 345034
rect 504822 328672 504878 328681
rect 504822 328607 504878 328616
rect 504362 328536 504418 328545
rect 504362 328471 504418 328480
rect 504376 328438 504404 328471
rect 504272 328432 504324 328438
rect 504272 328374 504324 328380
rect 504364 328432 504416 328438
rect 504364 328374 504416 328380
rect 504284 327078 504312 328374
rect 504272 327072 504324 327078
rect 504272 327014 504324 327020
rect 503720 321700 503772 321706
rect 503720 321642 503772 321648
rect 503996 321700 504048 321706
rect 503996 321642 504048 321648
rect 503904 321564 503956 321570
rect 503904 321506 503956 321512
rect 503720 317484 503772 317490
rect 503720 317426 503772 317432
rect 503628 311908 503680 311914
rect 503628 311850 503680 311856
rect 503640 311778 503668 311850
rect 503628 311772 503680 311778
rect 503628 311714 503680 311720
rect 503732 311658 503760 317426
rect 503640 311630 503760 311658
rect 503640 299538 503668 311630
rect 503628 299532 503680 299538
rect 503628 299474 503680 299480
rect 503812 299532 503864 299538
rect 503812 299474 503864 299480
rect 503824 292482 503852 299474
rect 503732 292454 503852 292482
rect 503732 283082 503760 292454
rect 503720 283076 503772 283082
rect 503720 283018 503772 283024
rect 503812 283008 503864 283014
rect 503812 282950 503864 282956
rect 503628 273352 503680 273358
rect 503628 273294 503680 273300
rect 503640 273222 503668 273294
rect 503628 273216 503680 273222
rect 503628 273158 503680 273164
rect 503720 263696 503772 263702
rect 503720 263638 503772 263644
rect 503732 263566 503760 263638
rect 503720 263560 503772 263566
rect 503720 263502 503772 263508
rect 503628 254040 503680 254046
rect 503628 253982 503680 253988
rect 503640 253910 503668 253982
rect 503628 253904 503680 253910
rect 503824 253858 503852 282950
rect 503628 253846 503680 253852
rect 503732 253830 503852 253858
rect 503732 244458 503760 253830
rect 503720 244452 503772 244458
rect 503720 244394 503772 244400
rect 503812 244384 503864 244390
rect 503812 244326 503864 244332
rect 503628 234728 503680 234734
rect 503628 234670 503680 234676
rect 503640 234598 503668 234670
rect 503628 234592 503680 234598
rect 503824 234546 503852 244326
rect 503628 234534 503680 234540
rect 503732 234518 503852 234546
rect 503732 225146 503760 234518
rect 503720 225140 503772 225146
rect 503720 225082 503772 225088
rect 503812 225072 503864 225078
rect 503812 225014 503864 225020
rect 503628 215416 503680 215422
rect 503628 215358 503680 215364
rect 503640 215286 503668 215358
rect 503628 215280 503680 215286
rect 503824 215234 503852 225014
rect 503628 215222 503680 215228
rect 503732 215206 503852 215234
rect 503732 205834 503760 215206
rect 503720 205828 503772 205834
rect 503720 205770 503772 205776
rect 503812 205760 503864 205766
rect 503812 205702 503864 205708
rect 503720 205692 503772 205698
rect 503720 205634 503772 205640
rect 457444 202496 457496 202502
rect 457444 202438 457496 202444
rect 503732 202230 503760 205634
rect 503824 202298 503852 205702
rect 503916 202366 503944 321506
rect 503996 318844 504048 318850
rect 503996 318786 504048 318792
rect 504008 311914 504036 318786
rect 504364 317484 504416 317490
rect 504364 317426 504416 317432
rect 504376 312662 504404 317426
rect 504364 312656 504416 312662
rect 504364 312598 504416 312604
rect 503996 311908 504048 311914
rect 503996 311850 504048 311856
rect 503996 311772 504048 311778
rect 503996 311714 504048 311720
rect 504008 273358 504036 311714
rect 504456 299532 504508 299538
rect 504456 299474 504508 299480
rect 504468 298110 504496 299474
rect 504456 298104 504508 298110
rect 504456 298046 504508 298052
rect 504548 288448 504600 288454
rect 504548 288390 504600 288396
rect 504560 280242 504588 288390
rect 504468 280214 504588 280242
rect 504468 278730 504496 280214
rect 504456 278724 504508 278730
rect 504456 278666 504508 278672
rect 503996 273352 504048 273358
rect 503996 273294 504048 273300
rect 503996 273216 504048 273222
rect 503996 273158 504048 273164
rect 504008 263702 504036 273158
rect 504640 269136 504692 269142
rect 504640 269078 504692 269084
rect 503996 263696 504048 263702
rect 503996 263638 504048 263644
rect 503996 263560 504048 263566
rect 503996 263502 504048 263508
rect 504008 254046 504036 263502
rect 504652 260953 504680 269078
rect 504270 260944 504326 260953
rect 504270 260879 504326 260888
rect 504638 260944 504694 260953
rect 504638 260879 504694 260888
rect 504284 260846 504312 260879
rect 504272 260840 504324 260846
rect 504272 260782 504324 260788
rect 503996 254040 504048 254046
rect 503996 253982 504048 253988
rect 503996 253904 504048 253910
rect 503996 253846 504048 253852
rect 504008 234734 504036 253846
rect 504272 253836 504324 253842
rect 504272 253778 504324 253784
rect 504284 251190 504312 253778
rect 504272 251184 504324 251190
rect 504272 251126 504324 251132
rect 504456 241528 504508 241534
rect 504456 241470 504508 241476
rect 504468 234734 504496 241470
rect 503996 234728 504048 234734
rect 503996 234670 504048 234676
rect 504456 234728 504508 234734
rect 504456 234670 504508 234676
rect 503996 234592 504048 234598
rect 503996 234534 504048 234540
rect 504364 234592 504416 234598
rect 504364 234534 504416 234540
rect 504008 215422 504036 234534
rect 504376 231810 504404 234534
rect 504364 231804 504416 231810
rect 504364 231746 504416 231752
rect 504456 222216 504508 222222
rect 504456 222158 504508 222164
rect 504468 215422 504496 222158
rect 503996 215416 504048 215422
rect 503996 215358 504048 215364
rect 504456 215416 504508 215422
rect 504456 215358 504508 215364
rect 503996 215280 504048 215286
rect 503996 215222 504048 215228
rect 504272 215280 504324 215286
rect 504272 215222 504324 215228
rect 504008 205698 504036 215222
rect 504284 212514 504312 215222
rect 504192 212486 504312 212514
rect 504192 205698 504220 212486
rect 503996 205692 504048 205698
rect 503996 205634 504048 205640
rect 504180 205692 504232 205698
rect 504180 205634 504232 205640
rect 504180 202904 504232 202910
rect 504180 202846 504232 202852
rect 503904 202360 503956 202366
rect 503904 202302 503956 202308
rect 503812 202292 503864 202298
rect 503812 202234 503864 202240
rect 503720 202224 503772 202230
rect 503720 202166 503772 202172
rect 504192 200462 504220 202846
rect 506492 202162 506520 520118
rect 506480 202156 506532 202162
rect 506480 202098 506532 202104
rect 504180 200456 504232 200462
rect 504180 200398 504232 200404
rect 504456 200456 504508 200462
rect 504456 200398 504508 200404
rect 504468 186266 504496 200398
rect 504376 186238 504496 186266
rect 504376 183569 504404 186238
rect 504362 183560 504418 183569
rect 504362 183495 504418 183504
rect 504638 183560 504694 183569
rect 504638 183495 504694 183504
rect 504652 173942 504680 183495
rect 504456 173936 504508 173942
rect 504456 173878 504508 173884
rect 504640 173936 504692 173942
rect 504640 173878 504692 173884
rect 504468 166954 504496 173878
rect 504376 166926 504496 166954
rect 504376 164218 504404 166926
rect 504180 164212 504232 164218
rect 504180 164154 504232 164160
rect 504364 164212 504416 164218
rect 504364 164154 504416 164160
rect 504192 154601 504220 164154
rect 504178 154592 504234 154601
rect 504178 154527 504234 154536
rect 504454 154592 504510 154601
rect 504454 154527 504510 154536
rect 447784 153196 447836 153202
rect 447784 153138 447836 153144
rect 446404 150408 446456 150414
rect 446404 150350 446456 150356
rect 445024 149048 445076 149054
rect 445024 148990 445076 148996
rect 442264 146192 442316 146198
rect 442264 146134 442316 146140
rect 438216 142112 438268 142118
rect 438216 142054 438268 142060
rect 437388 137964 437440 137970
rect 437388 137906 437440 137912
rect 437400 137873 437428 137906
rect 437386 137864 437442 137873
rect 437386 137799 437442 137808
rect 504468 136610 504496 154527
rect 514036 144906 514064 532714
rect 527192 200705 527220 703520
rect 543476 700369 543504 703520
rect 543462 700360 543518 700369
rect 559668 700330 559696 703520
rect 543462 700295 543518 700304
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 579698 580212 580751
rect 580172 579692 580224 579698
rect 580172 579634 580224 579640
rect 580262 557288 580318 557297
rect 580262 557223 580318 557232
rect 580170 533896 580226 533905
rect 580170 533831 580226 533840
rect 580184 532778 580212 533831
rect 580172 532772 580224 532778
rect 580172 532714 580224 532720
rect 580170 498672 580226 498681
rect 580170 498607 580226 498616
rect 580184 498234 580212 498607
rect 580172 498228 580224 498234
rect 580172 498170 580224 498176
rect 580170 486840 580226 486849
rect 580170 486775 580226 486784
rect 580184 485858 580212 486775
rect 580172 485852 580224 485858
rect 580172 485794 580224 485800
rect 579802 463448 579858 463457
rect 579802 463383 579858 463392
rect 579816 462398 579844 463383
rect 579804 462392 579856 462398
rect 579804 462334 579856 462340
rect 580170 451752 580226 451761
rect 580170 451687 580226 451696
rect 580184 451314 580212 451687
rect 580172 451308 580224 451314
rect 580172 451250 580224 451256
rect 580170 439920 580226 439929
rect 580170 439855 580226 439864
rect 580184 438938 580212 439855
rect 580172 438932 580224 438938
rect 580172 438874 580224 438880
rect 579802 416528 579858 416537
rect 579802 416463 579858 416472
rect 579816 415478 579844 416463
rect 579804 415472 579856 415478
rect 579804 415414 579856 415420
rect 579986 346080 580042 346089
rect 579986 346015 580042 346024
rect 580000 345098 580028 346015
rect 579988 345092 580040 345098
rect 579988 345034 580040 345040
rect 579618 322688 579674 322697
rect 579618 322623 579674 322632
rect 579632 321638 579660 322623
rect 579620 321632 579672 321638
rect 579620 321574 579672 321580
rect 579710 310856 579766 310865
rect 579710 310791 579766 310800
rect 579724 310554 579752 310791
rect 579712 310548 579764 310554
rect 579712 310490 579764 310496
rect 579618 275768 579674 275777
rect 579618 275703 579674 275712
rect 579632 274718 579660 275703
rect 579620 274712 579672 274718
rect 579620 274654 579672 274660
rect 580170 263936 580226 263945
rect 580170 263871 580226 263880
rect 580184 263634 580212 263871
rect 580172 263628 580224 263634
rect 580172 263570 580224 263576
rect 580170 228848 580226 228857
rect 580170 228783 580226 228792
rect 580184 227798 580212 228783
rect 580172 227792 580224 227798
rect 580172 227734 580224 227740
rect 579618 217016 579674 217025
rect 579618 216951 579674 216960
rect 579632 216714 579660 216951
rect 579620 216708 579672 216714
rect 579620 216650 579672 216656
rect 580276 200938 580304 557223
rect 580354 545592 580410 545601
rect 580354 545527 580410 545536
rect 580264 200932 580316 200938
rect 580264 200874 580316 200880
rect 580368 200802 580396 545527
rect 580446 510368 580502 510377
rect 580446 510303 580502 510312
rect 580460 200870 580488 510303
rect 580630 404832 580686 404841
rect 580630 404767 580686 404776
rect 580538 393000 580594 393009
rect 580538 392935 580594 392944
rect 580448 200864 580500 200870
rect 580448 200806 580500 200812
rect 580356 200796 580408 200802
rect 580356 200738 580408 200744
rect 527178 200696 527234 200705
rect 527178 200631 527234 200640
rect 580264 199844 580316 199850
rect 580264 199786 580316 199792
rect 580276 181937 580304 199786
rect 580262 181928 580318 181937
rect 580262 181863 580318 181872
rect 580262 170096 580318 170105
rect 580262 170031 580318 170040
rect 580170 158400 580226 158409
rect 580170 158335 580226 158344
rect 580184 157418 580212 158335
rect 580172 157412 580224 157418
rect 580172 157354 580224 157360
rect 514024 144900 514076 144906
rect 514024 144842 514076 144848
rect 437020 136604 437072 136610
rect 437020 136546 437072 136552
rect 504456 136604 504508 136610
rect 504456 136546 504508 136552
rect 437032 136105 437060 136546
rect 437018 136096 437074 136105
rect 437018 136031 437074 136040
rect 437388 133884 437440 133890
rect 437388 133826 437440 133832
rect 437400 133657 437428 133826
rect 437386 133648 437442 133657
rect 437386 133583 437442 133592
rect 437388 132456 437440 132462
rect 437388 132398 437440 132404
rect 437400 132025 437428 132398
rect 437386 132016 437442 132025
rect 437386 131951 437442 131960
rect 437388 129736 437440 129742
rect 437388 129678 437440 129684
rect 437400 129577 437428 129678
rect 437386 129568 437442 129577
rect 437386 129503 437442 129512
rect 436834 127800 436890 127809
rect 436834 127735 436890 127744
rect 436926 124536 436982 124545
rect 436926 124471 436982 124480
rect 436834 122904 436890 122913
rect 436834 122839 436890 122848
rect 436284 120624 436336 120630
rect 436284 120566 436336 120572
rect 436742 120456 436798 120465
rect 436742 120391 436798 120400
rect 436192 35896 436244 35902
rect 436192 35838 436244 35844
rect 436756 17950 436784 120391
rect 436848 64870 436876 122839
rect 436940 111790 436968 124471
rect 580276 120698 580304 170031
rect 580552 137970 580580 392935
rect 580644 341698 580672 404767
rect 580722 369608 580778 369617
rect 580722 369543 580778 369552
rect 580632 341692 580684 341698
rect 580632 341634 580684 341640
rect 580736 341562 580764 369543
rect 580814 357912 580870 357921
rect 580814 357847 580870 357856
rect 580828 341630 580856 357847
rect 580816 341624 580868 341630
rect 580816 341566 580868 341572
rect 580724 341556 580776 341562
rect 580724 341498 580776 341504
rect 580630 299160 580686 299169
rect 580630 299095 580686 299104
rect 580540 137964 580592 137970
rect 580540 137906 580592 137912
rect 580354 134872 580410 134881
rect 580354 134807 580410 134816
rect 580368 120766 580396 134807
rect 580644 133890 580672 299095
rect 580722 252240 580778 252249
rect 580722 252175 580778 252184
rect 580632 133884 580684 133890
rect 580632 133826 580684 133832
rect 580736 132462 580764 252175
rect 580814 205320 580870 205329
rect 580814 205255 580870 205264
rect 580724 132456 580776 132462
rect 580724 132398 580776 132404
rect 580828 129742 580856 205255
rect 580816 129736 580868 129742
rect 580816 129678 580868 129684
rect 580906 123176 580962 123185
rect 580906 123111 580962 123120
rect 580920 120834 580948 123111
rect 580908 120828 580960 120834
rect 580908 120770 580960 120776
rect 580356 120760 580408 120766
rect 580356 120702 580408 120708
rect 580264 120692 580316 120698
rect 580264 120634 580316 120640
rect 511264 118652 511316 118658
rect 511264 118594 511316 118600
rect 443000 118584 443052 118590
rect 443000 118526 443052 118532
rect 442262 118008 442318 118017
rect 442262 117943 442318 117952
rect 436928 111784 436980 111790
rect 436928 111726 436980 111732
rect 436836 64864 436888 64870
rect 436836 64806 436888 64812
rect 436744 17944 436796 17950
rect 436744 17886 436796 17892
rect 441804 8696 441856 8702
rect 441804 8638 441856 8644
rect 438216 8560 438268 8566
rect 438216 8502 438268 8508
rect 434628 8492 434680 8498
rect 434628 8434 434680 8440
rect 433522 4856 433578 4865
rect 433248 4820 433300 4826
rect 433522 4791 433578 4800
rect 433248 4762 433300 4768
rect 432328 3460 432380 3466
rect 432328 3402 432380 3408
rect 431222 3360 431278 3369
rect 431222 3295 431278 3304
rect 432340 480 432368 3402
rect 433536 480 433564 4791
rect 434640 480 434668 8434
rect 437020 7200 437072 7206
rect 437020 7142 437072 7148
rect 435824 7132 435876 7138
rect 435824 7074 435876 7080
rect 435836 480 435864 7074
rect 437032 480 437060 7142
rect 438228 480 438256 8502
rect 440608 7268 440660 7274
rect 440608 7210 440660 7216
rect 439412 3528 439464 3534
rect 439412 3470 439464 3476
rect 439424 480 439452 3470
rect 440620 480 440648 7210
rect 441816 480 441844 8638
rect 442276 7970 442304 117943
rect 442184 7942 442304 7970
rect 442184 3466 442212 7942
rect 442172 3460 442224 3466
rect 442172 3402 442224 3408
rect 443012 480 443040 118526
rect 475384 118516 475436 118522
rect 475384 118458 475436 118464
rect 449900 118380 449952 118386
rect 449900 118322 449952 118328
rect 448980 8764 449032 8770
rect 448980 8706 449032 8712
rect 445392 8628 445444 8634
rect 445392 8570 445444 8576
rect 444196 7336 444248 7342
rect 444196 7278 444248 7284
rect 444208 480 444236 7278
rect 445404 480 445432 8570
rect 447784 7404 447836 7410
rect 447784 7346 447836 7352
rect 446588 2848 446640 2854
rect 446588 2790 446640 2796
rect 446600 480 446628 2790
rect 447796 480 447824 7346
rect 448992 480 449020 8706
rect 449912 626 449940 118322
rect 474004 118312 474056 118318
rect 474004 118254 474056 118260
rect 469864 118244 469916 118250
rect 469864 118186 469916 118192
rect 456800 118176 456852 118182
rect 456800 118118 456852 118124
rect 454868 9648 454920 9654
rect 454868 9590 454920 9596
rect 452476 8832 452528 8838
rect 452476 8774 452528 8780
rect 451280 7472 451332 7478
rect 451280 7414 451332 7420
rect 449912 598 450216 626
rect 450188 480 450216 598
rect 451292 480 451320 7414
rect 452488 480 452516 8774
rect 453672 3052 453724 3058
rect 453672 2994 453724 3000
rect 453684 480 453712 2994
rect 454880 480 454908 9590
rect 456064 8900 456116 8906
rect 456064 8842 456116 8848
rect 456076 480 456104 8842
rect 456812 610 456840 118118
rect 463700 118108 463752 118114
rect 463700 118050 463752 118056
rect 463712 12442 463740 118050
rect 463700 12436 463752 12442
rect 463700 12378 463752 12384
rect 464344 12436 464396 12442
rect 464344 12378 464396 12384
rect 464356 12322 464384 12378
rect 464356 12294 464476 12322
rect 459652 10736 459704 10742
rect 459652 10678 459704 10684
rect 458456 9580 458508 9586
rect 458456 9522 458508 9528
rect 456800 604 456852 610
rect 456800 546 456852 552
rect 457260 604 457312 610
rect 457260 546 457312 552
rect 457272 480 457300 546
rect 458468 480 458496 9522
rect 459664 480 459692 10678
rect 463240 10668 463292 10674
rect 463240 10610 463292 10616
rect 462044 9512 462096 9518
rect 462044 9454 462096 9460
rect 460848 3120 460900 3126
rect 460848 3062 460900 3068
rect 460860 480 460888 3062
rect 462056 480 462084 9454
rect 463252 480 463280 10610
rect 464448 480 464476 12294
rect 466828 10600 466880 10606
rect 466828 10542 466880 10548
rect 465632 5636 465684 5642
rect 465632 5578 465684 5584
rect 465644 480 465672 5578
rect 466840 480 466868 10542
rect 469128 5568 469180 5574
rect 469128 5510 469180 5516
rect 467932 3188 467984 3194
rect 467932 3130 467984 3136
rect 467944 480 467972 3130
rect 469140 480 469168 5510
rect 469876 3126 469904 118186
rect 470600 118040 470652 118046
rect 470600 117982 470652 117988
rect 470324 10532 470376 10538
rect 470324 10474 470376 10480
rect 469864 3120 469916 3126
rect 469864 3062 469916 3068
rect 470336 480 470364 10474
rect 470612 610 470640 117982
rect 473360 10464 473412 10470
rect 473360 10406 473412 10412
rect 472716 5704 472768 5710
rect 472716 5646 472768 5652
rect 470600 604 470652 610
rect 470600 546 470652 552
rect 471520 604 471572 610
rect 471520 546 471572 552
rect 471532 480 471560 546
rect 472728 480 472756 5646
rect 473372 610 473400 10406
rect 474016 3194 474044 118254
rect 475396 3262 475424 118458
rect 478144 118448 478196 118454
rect 478144 118390 478196 118396
rect 477500 117972 477552 117978
rect 477500 117914 477552 117920
rect 477512 7546 477540 117914
rect 477684 10396 477736 10402
rect 477684 10338 477736 10344
rect 477500 7540 477552 7546
rect 477500 7482 477552 7488
rect 477696 7426 477724 10338
rect 477512 7398 477724 7426
rect 476304 5840 476356 5846
rect 476304 5782 476356 5788
rect 475108 3256 475160 3262
rect 475108 3198 475160 3204
rect 475384 3256 475436 3262
rect 475384 3198 475436 3204
rect 474004 3188 474056 3194
rect 474004 3130 474056 3136
rect 473360 604 473412 610
rect 473360 546 473412 552
rect 473912 604 473964 610
rect 473912 546 473964 552
rect 473924 480 473952 546
rect 475120 480 475148 3198
rect 476316 480 476344 5782
rect 477512 480 477540 7398
rect 478156 2990 478184 118390
rect 500224 117904 500276 117910
rect 500224 117846 500276 117852
rect 480904 117836 480956 117842
rect 480904 117778 480956 117784
rect 478696 7540 478748 7546
rect 478696 7482 478748 7488
rect 478144 2984 478196 2990
rect 478144 2926 478196 2932
rect 478708 480 478736 7482
rect 479892 5772 479944 5778
rect 479892 5714 479944 5720
rect 479904 480 479932 5714
rect 480916 2854 480944 117778
rect 493324 117700 493376 117706
rect 493324 117642 493376 117648
rect 482284 117632 482336 117638
rect 482284 117574 482336 117580
rect 481088 10328 481140 10334
rect 481088 10270 481140 10276
rect 480904 2848 480956 2854
rect 480904 2790 480956 2796
rect 481100 480 481128 10270
rect 482296 7698 482324 117574
rect 486424 117428 486476 117434
rect 486424 117370 486476 117376
rect 482204 7670 482324 7698
rect 482204 2990 482232 7670
rect 483480 7404 483532 7410
rect 483480 7346 483532 7352
rect 482284 3324 482336 3330
rect 482284 3266 482336 3272
rect 482192 2984 482244 2990
rect 482192 2926 482244 2932
rect 482296 480 482324 3266
rect 483492 480 483520 7346
rect 484584 5976 484636 5982
rect 484584 5918 484636 5924
rect 484596 480 484624 5918
rect 486436 3330 486464 117370
rect 489184 117360 489236 117366
rect 489184 117302 489236 117308
rect 486976 8288 487028 8294
rect 486976 8230 487028 8236
rect 486424 3324 486476 3330
rect 486424 3266 486476 3272
rect 485780 2916 485832 2922
rect 485780 2858 485832 2864
rect 485792 480 485820 2858
rect 486988 480 487016 8230
rect 488172 5908 488224 5914
rect 488172 5850 488224 5856
rect 488184 480 488212 5850
rect 489196 3058 489224 117302
rect 490564 8220 490616 8226
rect 490564 8162 490616 8168
rect 489368 3120 489420 3126
rect 489368 3062 489420 3068
rect 489184 3052 489236 3058
rect 489184 2994 489236 3000
rect 489380 480 489408 3062
rect 490576 480 490604 8162
rect 491760 6044 491812 6050
rect 491760 5986 491812 5992
rect 491772 480 491800 5986
rect 492956 3392 493008 3398
rect 492956 3334 493008 3340
rect 492968 480 492996 3334
rect 493336 3330 493364 117642
rect 496084 117564 496136 117570
rect 496084 117506 496136 117512
rect 494152 8152 494204 8158
rect 494152 8094 494204 8100
rect 493324 3324 493376 3330
rect 493324 3266 493376 3272
rect 494164 480 494192 8094
rect 495348 6112 495400 6118
rect 495348 6054 495400 6060
rect 495360 480 495388 6054
rect 496096 3398 496124 117506
rect 497740 8084 497792 8090
rect 497740 8026 497792 8032
rect 496084 3392 496136 3398
rect 496084 3334 496136 3340
rect 496544 3188 496596 3194
rect 496544 3130 496596 3136
rect 496556 480 496584 3130
rect 497752 480 497780 8026
rect 498936 6860 498988 6866
rect 498936 6802 498988 6808
rect 498948 480 498976 6802
rect 500236 4146 500264 117846
rect 502984 117768 503036 117774
rect 502984 117710 503036 117716
rect 501236 8016 501288 8022
rect 501236 7958 501288 7964
rect 500132 4140 500184 4146
rect 500132 4082 500184 4088
rect 500224 4140 500276 4146
rect 500224 4082 500276 4088
rect 500144 480 500172 4082
rect 501248 480 501276 7958
rect 502432 6792 502484 6798
rect 502432 6734 502484 6740
rect 502444 480 502472 6734
rect 502996 3330 503024 117710
rect 507124 117496 507176 117502
rect 507124 117438 507176 117444
rect 504824 7948 504876 7954
rect 504824 7890 504876 7896
rect 502984 3324 503036 3330
rect 502984 3266 503036 3272
rect 503628 3256 503680 3262
rect 503628 3198 503680 3204
rect 503640 480 503668 3198
rect 504836 480 504864 7890
rect 506020 6724 506072 6730
rect 506020 6666 506072 6672
rect 506032 480 506060 6666
rect 507136 4146 507164 117438
rect 508412 7880 508464 7886
rect 508412 7822 508464 7828
rect 507124 4140 507176 4146
rect 507124 4082 507176 4088
rect 507216 4072 507268 4078
rect 507216 4014 507268 4020
rect 507228 480 507256 4014
rect 508424 480 508452 7822
rect 509608 6656 509660 6662
rect 509608 6598 509660 6604
rect 509620 480 509648 6598
rect 511276 4078 511304 118594
rect 579804 111784 579856 111790
rect 579804 111726 579856 111732
rect 579816 111489 579844 111726
rect 579802 111480 579858 111489
rect 579802 111415 579858 111424
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 580172 77240 580224 77246
rect 580172 77182 580224 77188
rect 580184 76265 580212 77182
rect 580170 76256 580226 76265
rect 580170 76191 580226 76200
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 580172 30320 580224 30326
rect 580172 30262 580224 30268
rect 580184 29345 580212 30262
rect 580170 29336 580226 29345
rect 580170 29271 580226 29280
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 552388 9444 552440 9450
rect 552388 9386 552440 9392
rect 541716 7812 541768 7818
rect 541716 7754 541768 7760
rect 513196 6588 513248 6594
rect 513196 6530 513248 6536
rect 512000 4208 512052 4214
rect 512000 4150 512052 4156
rect 511264 4072 511316 4078
rect 511264 4014 511316 4020
rect 510804 2984 510856 2990
rect 510804 2926 510856 2932
rect 510816 480 510844 2926
rect 512012 480 512040 4150
rect 513208 480 513236 6530
rect 516784 6520 516836 6526
rect 516784 6462 516836 6468
rect 515588 4276 515640 4282
rect 515588 4218 515640 4224
rect 514392 4004 514444 4010
rect 514392 3946 514444 3952
rect 514404 480 514432 3946
rect 515600 480 515628 4218
rect 516796 480 516824 6462
rect 520280 6452 520332 6458
rect 520280 6394 520332 6400
rect 519084 4412 519136 4418
rect 519084 4354 519136 4360
rect 517888 2848 517940 2854
rect 517888 2790 517940 2796
rect 517900 480 517928 2790
rect 519096 480 519124 4354
rect 520292 480 520320 6394
rect 523868 6384 523920 6390
rect 523868 6326 523920 6332
rect 522672 4344 522724 4350
rect 522672 4286 522724 4292
rect 521476 3936 521528 3942
rect 521476 3878 521528 3884
rect 521488 480 521516 3878
rect 522684 480 522712 4286
rect 523880 480 523908 6326
rect 531044 6316 531096 6322
rect 531044 6258 531096 6264
rect 527456 6248 527508 6254
rect 527456 6190 527508 6196
rect 526260 4480 526312 4486
rect 526260 4422 526312 4428
rect 525064 2916 525116 2922
rect 525064 2858 525116 2864
rect 525076 480 525104 2858
rect 526272 480 526300 4422
rect 527468 480 527496 6190
rect 529848 4548 529900 4554
rect 529848 4490 529900 4496
rect 528652 3868 528704 3874
rect 528652 3810 528704 3816
rect 528664 480 528692 3810
rect 529860 480 529888 4490
rect 531056 480 531084 6258
rect 538126 6216 538182 6225
rect 534540 6180 534592 6186
rect 538126 6151 538182 6160
rect 534540 6122 534592 6128
rect 533436 4616 533488 4622
rect 533436 4558 533488 4564
rect 532240 3052 532292 3058
rect 532240 2994 532292 3000
rect 532252 480 532280 2994
rect 533448 480 533476 4558
rect 534552 480 534580 6122
rect 536932 4684 536984 4690
rect 536932 4626 536984 4632
rect 535736 3800 535788 3806
rect 535736 3742 535788 3748
rect 535748 480 535776 3742
rect 536944 480 536972 4626
rect 538140 480 538168 6151
rect 540520 4752 540572 4758
rect 540520 4694 540572 4700
rect 539324 3120 539376 3126
rect 539324 3062 539376 3068
rect 539336 480 539364 3062
rect 540532 480 540560 4694
rect 541728 480 541756 7754
rect 545304 7744 545356 7750
rect 545304 7686 545356 7692
rect 544108 5500 544160 5506
rect 544108 5442 544160 5448
rect 542912 3732 542964 3738
rect 542912 3674 542964 3680
rect 542924 480 542952 3674
rect 544120 480 544148 5442
rect 545316 480 545344 7686
rect 548892 7676 548944 7682
rect 548892 7618 548944 7624
rect 547696 5432 547748 5438
rect 547696 5374 547748 5380
rect 546500 3188 546552 3194
rect 546500 3130 546552 3136
rect 546512 480 546540 3130
rect 547708 480 547736 5374
rect 548904 480 548932 7618
rect 551192 5364 551244 5370
rect 551192 5306 551244 5312
rect 550088 3256 550140 3262
rect 550088 3198 550140 3204
rect 550100 480 550128 3198
rect 551204 480 551232 5306
rect 552400 480 552428 9386
rect 555976 9376 556028 9382
rect 555976 9318 556028 9324
rect 554780 5296 554832 5302
rect 554780 5238 554832 5244
rect 553584 3664 553636 3670
rect 553584 3606 553636 3612
rect 553596 480 553624 3606
rect 554792 480 554820 5238
rect 555988 480 556016 9318
rect 559564 9308 559616 9314
rect 559564 9250 559616 9256
rect 558368 5228 558420 5234
rect 558368 5170 558420 5176
rect 557172 3324 557224 3330
rect 557172 3266 557224 3272
rect 557184 480 557212 3266
rect 558380 480 558408 5170
rect 559576 480 559604 9250
rect 563152 9240 563204 9246
rect 563152 9182 563204 9188
rect 561956 5092 562008 5098
rect 561956 5034 562008 5040
rect 560760 3596 560812 3602
rect 560760 3538 560812 3544
rect 560772 480 560800 3538
rect 561968 480 561996 5034
rect 563164 480 563192 9182
rect 566740 9172 566792 9178
rect 566740 9114 566792 9120
rect 565544 5160 565596 5166
rect 565544 5102 565596 5108
rect 564348 3392 564400 3398
rect 564348 3334 564400 3340
rect 564360 480 564388 3334
rect 565556 480 565584 5102
rect 566752 480 566780 9114
rect 570236 9104 570288 9110
rect 570236 9046 570288 9052
rect 569040 5024 569092 5030
rect 569040 4966 569092 4972
rect 567844 3528 567896 3534
rect 567844 3470 567896 3476
rect 567856 480 567884 3470
rect 569052 480 569080 4966
rect 570248 480 570276 9046
rect 577412 9036 577464 9042
rect 577412 8978 577464 8984
rect 573824 7608 573876 7614
rect 573824 7550 573876 7556
rect 572628 4956 572680 4962
rect 572628 4898 572680 4904
rect 571432 4140 571484 4146
rect 571432 4082 571484 4088
rect 571444 480 571472 4082
rect 572640 480 572668 4898
rect 573836 480 573864 7550
rect 576216 4888 576268 4894
rect 576216 4830 576268 4836
rect 575018 3360 575074 3369
rect 575018 3295 575074 3304
rect 575032 480 575060 3295
rect 576228 480 576256 4830
rect 577424 480 577452 8978
rect 581000 8968 581052 8974
rect 581000 8910 581052 8916
rect 579804 4820 579856 4826
rect 579804 4762 579856 4768
rect 578608 4072 578660 4078
rect 578608 4014 578660 4020
rect 578620 480 578648 4014
rect 579816 480 579844 4762
rect 581012 480 581040 8910
rect 582196 3460 582248 3466
rect 582196 3402 582248 3408
rect 582208 480 582236 3402
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3514 682216 3570 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 4802 653520 4858 653576
rect 3422 624824 3478 624880
rect 3422 610408 3478 610464
rect 4066 595992 4122 596048
rect 3422 567296 3478 567352
rect 3146 553016 3202 553072
rect 3330 495508 3386 495544
rect 3330 495488 3332 495508
rect 3332 495488 3384 495508
rect 3384 495488 3386 495508
rect 3054 452376 3110 452432
rect 2778 366152 2834 366208
rect 2962 337456 3018 337512
rect 3330 294344 3386 294400
rect 2778 265648 2834 265704
rect 3330 251252 3386 251288
rect 3330 251232 3332 251252
rect 3332 251232 3384 251252
rect 3384 251232 3386 251252
rect 3330 236952 3386 237008
rect 2962 222536 3018 222592
rect 2962 208120 3018 208176
rect 2870 179424 2926 179480
rect 3238 165008 3294 165064
rect 3514 538600 3570 538656
rect 3238 150728 3294 150784
rect 3330 136312 3386 136368
rect 3330 122032 3386 122088
rect 2778 93200 2834 93256
rect 3238 78920 3294 78976
rect 3330 64504 3386 64560
rect 3606 509904 3662 509960
rect 4066 481072 4122 481128
rect 3698 437960 3754 438016
rect 3606 193840 3662 193896
rect 4066 423700 4122 423736
rect 4066 423680 4068 423700
rect 4068 423680 4120 423700
rect 4120 423680 4122 423700
rect 3882 394984 3938 395040
rect 3790 380568 3846 380624
rect 3974 323040 4030 323096
rect 4066 308760 4122 308816
rect 4066 280064 4122 280120
rect 3514 107616 3570 107672
rect 3422 50088 3478 50144
rect 3422 35844 3424 35864
rect 3424 35844 3476 35864
rect 3476 35844 3478 35864
rect 3422 35808 3478 35844
rect 3146 21392 3202 21448
rect 3422 7112 3478 7168
rect 30286 4800 30342 4856
rect 69938 385192 69994 385248
rect 70214 377848 70270 377904
rect 70122 370232 70178 370288
rect 70030 362888 70086 362944
rect 70214 355544 70270 355600
rect 71594 392536 71650 392592
rect 71042 377848 71098 377904
rect 70306 348200 70362 348256
rect 70214 341944 70270 342000
rect 69662 118496 69718 118552
rect 71594 370232 71650 370288
rect 71502 348200 71558 348256
rect 84106 545808 84162 545864
rect 84014 541456 84070 541512
rect 83922 528672 83978 528728
rect 82818 524864 82874 524920
rect 85302 533024 85358 533080
rect 85394 525544 85450 525600
rect 86406 549908 86462 549944
rect 86406 549888 86408 549908
rect 86408 549888 86460 549908
rect 86460 549888 86462 549908
rect 85578 537716 85634 537772
rect 118054 546488 118110 546544
rect 117318 537376 117374 537432
rect 117318 533296 117374 533352
rect 117962 529488 118018 529544
rect 117318 525136 117374 525192
rect 117318 521056 117374 521112
rect 118238 542408 118294 542464
rect 118238 521600 118294 521656
rect 118422 521600 118478 521656
rect 118422 498072 118478 498128
rect 118330 482976 118386 483032
rect 118606 482976 118662 483032
rect 118054 454008 118110 454064
rect 118238 454008 118294 454064
rect 118054 434696 118110 434752
rect 118238 434696 118294 434752
rect 99286 118632 99342 118688
rect 71594 117816 71650 117872
rect 79966 117816 80022 117872
rect 80150 117680 80206 117736
rect 89810 117816 89866 117872
rect 89626 117680 89682 117736
rect 99194 117852 99196 117872
rect 99196 117852 99248 117872
rect 99248 117852 99250 117872
rect 99194 117816 99250 117852
rect 110326 118360 110382 118416
rect 101218 117852 101220 117872
rect 101220 117852 101272 117872
rect 101272 117852 101274 117872
rect 101218 117816 101274 117852
rect 103518 117816 103574 117872
rect 97998 117272 98054 117328
rect 99286 117272 99342 117328
rect 104990 117700 105046 117736
rect 104990 117680 104992 117700
rect 104992 117680 105044 117700
rect 105044 117680 105046 117700
rect 115202 117816 115258 117872
rect 124218 153992 124274 154048
rect 122838 117816 122894 117872
rect 102782 6160 102838 6216
rect 128542 511944 128598 512000
rect 128726 511944 128782 512000
rect 129646 582392 129702 582448
rect 128542 482976 128598 483032
rect 128818 482976 128874 483032
rect 128542 463664 128598 463720
rect 128818 463664 128874 463720
rect 128542 444352 128598 444408
rect 128818 444352 128874 444408
rect 128542 425040 128598 425096
rect 128818 425040 128874 425096
rect 128726 388476 128782 388512
rect 128726 388456 128728 388476
rect 128728 388456 128780 388476
rect 128780 388456 128782 388476
rect 129094 380568 129150 380624
rect 128450 373224 128506 373280
rect 128358 358264 128414 358320
rect 129002 350920 129058 350976
rect 129002 343576 129058 343632
rect 126518 182144 126574 182200
rect 126794 182144 126850 182200
rect 126426 153176 126482 153232
rect 126702 153040 126758 153096
rect 128174 144472 128230 144528
rect 126518 143520 126574 143576
rect 126702 143520 126758 143576
rect 128910 299376 128966 299432
rect 128818 289856 128874 289912
rect 128910 280064 128966 280120
rect 129002 279928 129058 279984
rect 128542 190440 128598 190496
rect 128726 190440 128782 190496
rect 128266 118224 128322 118280
rect 126058 117544 126114 117600
rect 129186 373224 129242 373280
rect 129370 365880 129426 365936
rect 129278 358264 129334 358320
rect 127622 117272 127678 117328
rect 128266 117272 128322 117328
rect 128634 67632 128690 67688
rect 128818 67632 128874 67688
rect 131026 500248 131082 500304
rect 130934 500112 130990 500168
rect 130290 341944 130346 342000
rect 130474 196152 130530 196208
rect 130474 194656 130530 194712
rect 130474 194420 130476 194440
rect 130476 194420 130528 194440
rect 130528 194420 130530 194440
rect 130474 194384 130530 194420
rect 130474 193060 130476 193080
rect 130476 193060 130528 193080
rect 130528 193060 130530 193080
rect 130474 193024 130530 193060
rect 130382 192480 130438 192536
rect 130474 191392 130530 191448
rect 130474 190304 130530 190360
rect 130474 188808 130530 188864
rect 130382 188264 130438 188320
rect 130474 187176 130530 187232
rect 129462 117680 129518 117736
rect 131210 185544 131266 185600
rect 131210 184456 131266 184512
rect 131210 183524 131266 183560
rect 131210 183504 131212 183524
rect 131212 183504 131264 183524
rect 131264 183504 131266 183524
rect 131210 178200 131266 178256
rect 131394 198192 131450 198248
rect 131394 197104 131450 197160
rect 131302 164464 131358 164520
rect 131210 161336 131266 161392
rect 131302 157120 131358 157176
rect 131118 156168 131174 156224
rect 131118 155080 131174 155136
rect 131118 152904 131174 152960
rect 131210 151952 131266 152008
rect 131118 150864 131174 150920
rect 131118 149776 131174 149832
rect 131118 148688 131174 148744
rect 131118 147736 131174 147792
rect 131118 146648 131174 146704
rect 131118 145560 131174 145616
rect 131118 143520 131174 143576
rect 131302 139304 131358 139360
rect 131394 131960 131450 132016
rect 131762 199280 131818 199336
rect 131670 167728 131726 167784
rect 131670 158208 131726 158264
rect 131578 125568 131634 125624
rect 131486 124480 131542 124536
rect 131118 124208 131174 124264
rect 131302 124208 131358 124264
rect 131210 96600 131266 96656
rect 131394 96600 131450 96656
rect 131946 128696 132002 128752
rect 132222 170856 132278 170912
rect 132222 159296 132278 159352
rect 132130 130872 132186 130928
rect 132038 127744 132094 127800
rect 131854 126656 131910 126712
rect 132130 121352 132186 121408
rect 132498 179288 132554 179344
rect 132590 177112 132646 177168
rect 132406 171944 132462 172000
rect 132958 168680 133014 168736
rect 132774 166640 132830 166696
rect 132682 165552 132738 165608
rect 132406 162424 132462 162480
rect 132314 138216 132370 138272
rect 132406 120400 132462 120456
rect 132866 118088 132922 118144
rect 133142 169768 133198 169824
rect 133326 182416 133382 182472
rect 133418 181328 133474 181384
rect 133602 163512 133658 163568
rect 133602 160384 133658 160440
rect 133510 142432 133566 142488
rect 133234 129784 133290 129840
rect 133326 118088 133382 118144
rect 133050 117952 133106 118008
rect 133694 141344 133750 141400
rect 147586 697076 147588 697096
rect 147588 697076 147640 697096
rect 147640 697076 147642 697096
rect 147586 697040 147642 697076
rect 154486 697176 154542 697232
rect 173806 697176 173862 697232
rect 193126 697176 193182 697232
rect 212446 697176 212502 697232
rect 231766 697176 231822 697232
rect 251086 697176 251142 697232
rect 270406 697176 270462 697232
rect 289726 697176 289782 697232
rect 309046 697176 309102 697232
rect 328366 697176 328422 697232
rect 166906 697076 166908 697096
rect 166908 697076 166960 697096
rect 166960 697076 166962 697096
rect 166906 697040 166962 697076
rect 186226 697076 186228 697096
rect 186228 697076 186280 697096
rect 186280 697076 186282 697096
rect 186226 697040 186282 697076
rect 205546 697076 205548 697096
rect 205548 697076 205600 697096
rect 205600 697076 205602 697096
rect 205546 697040 205602 697076
rect 224866 697076 224868 697096
rect 224868 697076 224920 697096
rect 224920 697076 224922 697096
rect 224866 697040 224922 697076
rect 244186 697076 244188 697096
rect 244188 697076 244240 697096
rect 244240 697076 244242 697096
rect 244186 697040 244242 697076
rect 263506 697076 263508 697096
rect 263508 697076 263560 697096
rect 263560 697076 263562 697096
rect 263506 697040 263562 697076
rect 282826 697076 282828 697096
rect 282828 697076 282880 697096
rect 282880 697076 282882 697096
rect 282826 697040 282882 697076
rect 302146 697076 302148 697096
rect 302148 697076 302200 697096
rect 302200 697076 302202 697096
rect 302146 697040 302202 697076
rect 321466 697076 321468 697096
rect 321468 697076 321520 697096
rect 321520 697076 321522 697096
rect 321466 697040 321522 697076
rect 135258 686180 135314 686216
rect 135258 686160 135260 686180
rect 135260 686160 135312 686180
rect 135312 686160 135314 686180
rect 147770 686296 147826 686352
rect 147586 686024 147642 686080
rect 169022 686432 169078 686488
rect 154578 686316 154634 686352
rect 154578 686296 154580 686316
rect 154580 686296 154632 686316
rect 154632 686296 154634 686316
rect 159454 686160 159510 686216
rect 169022 686160 169078 686216
rect 142894 685888 142950 685944
rect 169022 650528 169078 650584
rect 135258 650276 135314 650312
rect 135258 650256 135260 650276
rect 135260 650256 135312 650276
rect 135312 650256 135314 650276
rect 147770 650392 147826 650448
rect 154578 650412 154634 650448
rect 154578 650392 154580 650412
rect 154580 650392 154632 650412
rect 154632 650392 154634 650412
rect 159454 650256 159510 650312
rect 169022 650256 169078 650312
rect 147586 650120 147642 650176
rect 142894 649984 142950 650040
rect 157062 639240 157118 639296
rect 157246 639240 157302 639296
rect 171046 639240 171102 639296
rect 171046 638832 171102 638888
rect 157062 603336 157118 603392
rect 157246 603336 157302 603392
rect 171046 603336 171102 603392
rect 171046 602928 171102 602984
rect 153382 598848 153438 598904
rect 153566 598848 153622 598904
rect 157062 592320 157118 592376
rect 157246 592320 157302 592376
rect 171046 592320 171102 592376
rect 171046 591912 171102 591968
rect 133970 180648 134026 180704
rect 133786 140392 133842 140448
rect 133970 122984 134026 123040
rect 153474 531256 153530 531312
rect 153750 531256 153806 531312
rect 153290 482976 153346 483032
rect 153474 482976 153530 483032
rect 153474 425176 153530 425232
rect 153198 425040 153254 425096
rect 197082 202816 197138 202872
rect 196990 202680 197046 202736
rect 211618 561720 211674 561776
rect 222198 556144 222254 556200
rect 198646 534112 198702 534168
rect 198554 524592 198610 524648
rect 198002 378664 198058 378720
rect 197910 374312 197966 374368
rect 197818 370232 197874 370288
rect 197726 361800 197782 361856
rect 197542 357448 197598 357504
rect 197450 353368 197506 353424
rect 197358 349016 197414 349072
rect 197634 344936 197690 344992
rect 197266 202408 197322 202464
rect 197174 202136 197230 202192
rect 198462 399608 198518 399664
rect 198370 387096 198426 387152
rect 198738 529216 198794 529272
rect 198830 403688 198886 403744
rect 198922 395256 198978 395312
rect 199014 391176 199070 391232
rect 199106 382744 199162 382800
rect 199198 365880 199254 365936
rect 203338 410352 203394 410408
rect 222290 552064 222346 552120
rect 222566 546896 222622 546952
rect 222474 542544 222530 542600
rect 222382 538328 222438 538384
rect 222658 533296 222714 533352
rect 222750 528944 222806 529000
rect 222842 524456 222898 524512
rect 226154 410080 226210 410136
rect 231858 410216 231914 410272
rect 263138 409944 263194 410000
rect 209778 241440 209834 241496
rect 209962 241440 210018 241496
rect 209778 222128 209834 222184
rect 209962 222128 210018 222184
rect 211158 201592 211214 201648
rect 212538 201864 212594 201920
rect 213458 201728 213514 201784
rect 218058 202000 218114 202056
rect 220358 202816 220414 202872
rect 237194 338680 237250 338736
rect 223854 202680 223910 202736
rect 225142 202544 225198 202600
rect 226338 202408 226394 202464
rect 232134 202272 232190 202328
rect 232410 201864 232466 201920
rect 233422 202136 233478 202192
rect 238666 201864 238722 201920
rect 257710 317328 257766 317384
rect 257802 311752 257858 311808
rect 257802 220768 257858 220824
rect 257986 220768 258042 220824
rect 257066 202136 257122 202192
rect 262678 201592 262734 201648
rect 266174 201456 266230 201512
rect 267186 399608 267242 399664
rect 267278 357448 267334 357504
rect 267370 353368 267426 353424
rect 267462 349016 267518 349072
rect 267830 403688 267886 403744
rect 267922 395256 267978 395312
rect 268014 391176 268070 391232
rect 268106 386824 268162 386880
rect 268198 382744 268254 382800
rect 268290 378392 268346 378448
rect 268382 374312 268438 374368
rect 268474 369960 268530 370016
rect 268566 365880 268622 365936
rect 268658 361528 268714 361584
rect 269026 344936 269082 344992
rect 274546 582528 274602 582584
rect 288346 392128 288402 392184
rect 288162 391992 288218 392048
rect 288346 382200 288402 382256
rect 288530 382200 288586 382256
rect 288254 231784 288310 231840
rect 288530 231784 288586 231840
rect 296718 575728 296774 575784
rect 297454 572872 297510 572928
rect 296442 565800 296498 565856
rect 296902 563352 296958 563408
rect 297086 556824 297142 556880
rect 297362 541048 297418 541104
rect 296534 531392 296590 531448
rect 297086 522144 297142 522200
rect 298006 570016 298062 570072
rect 298006 560360 298062 560416
rect 297914 553560 297970 553616
rect 297822 544040 297878 544096
rect 297730 538328 297786 538384
rect 297454 528808 297510 528864
rect 297730 519152 297786 519208
rect 297730 516180 297786 516216
rect 297730 516160 297732 516180
rect 297732 516160 297784 516180
rect 297784 516160 297786 516180
rect 297730 513440 297786 513496
rect 297638 509632 297694 509688
rect 297638 506640 297694 506696
rect 299294 550704 299350 550760
rect 299202 547848 299258 547904
rect 299110 525816 299166 525872
rect 299570 535404 299626 535460
rect 299662 503852 299718 503908
rect 349526 582392 349582 582448
rect 368662 582528 368718 582584
rect 304170 492632 304226 492688
rect 304538 492632 304594 492688
rect 304262 473340 304318 473376
rect 304262 473320 304264 473340
rect 304264 473320 304316 473340
rect 304316 473320 304318 473340
rect 304446 473320 304502 473376
rect 304170 338034 304226 338090
rect 304446 337864 304502 337920
rect 304078 260888 304134 260944
rect 304446 260888 304502 260944
rect 304262 231784 304318 231840
rect 304538 231784 304594 231840
rect 319718 498072 319774 498128
rect 377310 565800 377366 565856
rect 377402 563080 377458 563136
rect 378138 560156 378194 560212
rect 377494 556552 377550 556608
rect 378230 550636 378286 550692
rect 378322 547644 378378 547700
rect 380622 575456 380678 575512
rect 379518 569064 379574 569120
rect 378966 515480 379022 515536
rect 379610 553424 379666 553480
rect 379702 543768 379758 543824
rect 379794 537512 379850 537568
rect 379886 534520 379942 534576
rect 379978 531392 380034 531448
rect 380530 528672 380586 528728
rect 380070 525000 380126 525056
rect 380162 521736 380218 521792
rect 380254 512488 380310 512544
rect 380346 509360 380402 509416
rect 380438 506504 380494 506560
rect 380714 519152 380770 519208
rect 380714 502968 380770 503024
rect 380898 381384 380954 381440
rect 380898 377168 380954 377224
rect 380898 374060 380954 374096
rect 380898 374040 380900 374060
rect 380900 374040 380952 374060
rect 380952 374040 380954 374060
rect 380898 370368 380954 370424
rect 381634 367376 381690 367432
rect 380898 363568 380954 363624
rect 380898 353504 380954 353560
rect 381726 360304 381782 360360
rect 381818 356768 381874 356824
rect 415398 363908 415454 363964
rect 416870 380840 416926 380896
rect 416778 376896 416834 376952
rect 416962 374584 417018 374640
rect 416870 370096 416926 370152
rect 416962 367104 417018 367160
rect 417054 360168 417110 360224
rect 417146 356496 417202 356552
rect 417238 353368 417294 353424
rect 434258 169632 434314 169688
rect 434534 186224 434590 186280
rect 434994 196152 435050 196208
rect 434902 184592 434958 184648
rect 434810 173848 434866 173904
rect 434718 171944 434774 172000
rect 434442 167728 434498 167784
rect 434350 165552 434406 165608
rect 434166 163512 434222 163568
rect 434074 161200 434130 161256
rect 433982 159296 434038 159352
rect 433890 157256 433946 157312
rect 134062 121896 134118 121952
rect 133786 117816 133842 117872
rect 133786 106256 133842 106312
rect 133970 117680 134026 117736
rect 134154 117680 134210 117736
rect 133970 106276 134026 106312
rect 133970 106256 133972 106276
rect 133972 106256 134024 106276
rect 134024 106256 134026 106276
rect 138524 119720 138580 119776
rect 140870 38528 140926 38584
rect 140962 29008 141018 29064
rect 145562 118360 145618 118416
rect 151910 117680 151966 117736
rect 149058 4800 149114 4856
rect 153474 118496 153530 118552
rect 157522 115912 157578 115968
rect 157890 115912 157946 115968
rect 157338 70352 157394 70408
rect 157338 66272 157394 66328
rect 161754 115912 161810 115968
rect 162122 115912 162178 115968
rect 175278 117952 175334 118008
rect 179694 37440 179750 37496
rect 179418 37304 179474 37360
rect 184938 118632 184994 118688
rect 183834 115912 183890 115968
rect 184110 115912 184166 115968
rect 186410 6160 186466 6216
rect 188434 118088 188490 118144
rect 190918 96736 190974 96792
rect 190642 96600 190698 96656
rect 193954 118224 194010 118280
rect 197634 117544 197690 117600
rect 214102 86944 214158 87000
rect 214286 86944 214342 87000
rect 216954 115912 217010 115968
rect 217322 115912 217378 115968
rect 220726 53896 220782 53952
rect 221002 115912 221058 115968
rect 221462 115912 221518 115968
rect 221002 53896 221058 53952
rect 221002 53760 221058 53816
rect 221186 53760 221242 53816
rect 221002 34448 221058 34504
rect 221186 34448 221242 34504
rect 227902 34584 227958 34640
rect 228178 34584 228234 34640
rect 230386 35808 230442 35864
rect 230478 26288 230534 26344
rect 230662 35672 230718 35728
rect 230662 26288 230718 26344
rect 243634 117272 243690 117328
rect 245750 117272 245806 117328
rect 248418 96600 248474 96656
rect 248602 96600 248658 96656
rect 276018 106392 276074 106448
rect 275006 106256 275062 106312
rect 275374 106256 275430 106312
rect 276110 106256 276166 106312
rect 274730 96600 274786 96656
rect 275006 96600 275062 96656
rect 276110 48320 276166 48376
rect 276294 48320 276350 48376
rect 290646 99456 290702 99512
rect 290554 96620 290610 96656
rect 290554 96600 290556 96620
rect 290556 96600 290608 96620
rect 290608 96600 290610 96620
rect 290554 67632 290610 67688
rect 290462 66272 290518 66328
rect 301410 116048 301466 116104
rect 301778 115912 301834 115968
rect 301870 26288 301926 26344
rect 302054 26288 302110 26344
rect 325514 48320 325570 48376
rect 325698 48320 325754 48376
rect 341430 99456 341486 99512
rect 341338 96620 341394 96656
rect 341338 96600 341340 96620
rect 341340 96600 341392 96620
rect 341392 96600 341394 96620
rect 341062 86944 341118 87000
rect 341246 86944 341302 87000
rect 357346 4800 357402 4856
rect 388350 116048 388406 116104
rect 388718 115932 388774 115968
rect 388718 115912 388720 115932
rect 388720 115912 388772 115932
rect 388772 115912 388774 115932
rect 388718 106276 388774 106312
rect 388718 106256 388720 106276
rect 388720 106256 388772 106276
rect 388772 106256 388774 106276
rect 388902 106256 388958 106312
rect 408314 3712 408370 3768
rect 408498 3712 408554 3768
rect 411074 6160 411130 6216
rect 415030 48320 415086 48376
rect 415214 48320 415270 48376
rect 417882 3576 417938 3632
rect 418158 117716 418160 117736
rect 418160 117716 418212 117736
rect 418212 117716 418214 117736
rect 418158 117680 418214 117716
rect 418342 3576 418398 3632
rect 420274 77288 420330 77344
rect 420458 77288 420514 77344
rect 420642 61376 420698 61432
rect 420550 48320 420606 48376
rect 420642 42064 420698 42120
rect 420550 29008 420606 29064
rect 426070 48320 426126 48376
rect 426254 48320 426310 48376
rect 427726 117700 427782 117736
rect 427726 117680 427728 117700
rect 427728 117680 427780 117700
rect 427780 117680 427782 117700
rect 427634 3596 427690 3632
rect 427634 3576 427636 3596
rect 427636 3576 427688 3596
rect 427688 3576 427690 3596
rect 427818 3576 427874 3632
rect 431590 46960 431646 47016
rect 431774 46960 431830 47016
rect 433982 117952 434038 118008
rect 435178 190168 435234 190224
rect 435086 188808 435142 188864
rect 436190 198872 436246 198928
rect 436098 180240 436154 180296
rect 436098 155080 436154 155136
rect 436098 148688 436154 148744
rect 436098 142060 436100 142080
rect 436100 142060 436152 142080
rect 436152 142060 436154 142080
rect 436098 142024 436154 142060
rect 436282 193976 436338 194032
rect 436650 193024 436706 193080
rect 436558 182008 436614 182064
rect 436466 177928 436522 177984
rect 436374 176160 436430 176216
rect 436742 140392 436798 140448
rect 478510 700440 478566 700496
rect 437386 152768 437442 152824
rect 437386 150184 437442 150240
rect 437386 146240 437442 146296
rect 437018 144472 437074 144528
rect 456798 375128 456854 375184
rect 504730 378392 504786 378448
rect 457442 357992 457498 358048
rect 504730 360440 504786 360496
rect 503718 340856 503774 340912
rect 504730 343576 504786 343632
rect 503902 340856 503958 340912
rect 504822 328616 504878 328672
rect 504362 328480 504418 328536
rect 504270 260888 504326 260944
rect 504638 260888 504694 260944
rect 504362 183504 504418 183560
rect 504638 183504 504694 183560
rect 504178 154536 504234 154592
rect 504454 154536 504510 154592
rect 437386 137808 437442 137864
rect 543462 700304 543518 700360
rect 580170 674600 580226 674656
rect 580170 627680 580226 627736
rect 580170 580760 580226 580816
rect 580262 557232 580318 557288
rect 580170 533840 580226 533896
rect 580170 498616 580226 498672
rect 580170 486784 580226 486840
rect 579802 463392 579858 463448
rect 580170 451696 580226 451752
rect 580170 439864 580226 439920
rect 579802 416472 579858 416528
rect 579986 346024 580042 346080
rect 579618 322632 579674 322688
rect 579710 310800 579766 310856
rect 579618 275712 579674 275768
rect 580170 263880 580226 263936
rect 580170 228792 580226 228848
rect 579618 216960 579674 217016
rect 580354 545536 580410 545592
rect 580446 510312 580502 510368
rect 580630 404776 580686 404832
rect 580538 392944 580594 393000
rect 527178 200640 527234 200696
rect 580262 181872 580318 181928
rect 580262 170040 580318 170096
rect 580170 158344 580226 158400
rect 437018 136040 437074 136096
rect 437386 133592 437442 133648
rect 437386 131960 437442 132016
rect 437386 129512 437442 129568
rect 436834 127744 436890 127800
rect 436926 124480 436982 124536
rect 436834 122848 436890 122904
rect 436742 120400 436798 120456
rect 580722 369552 580778 369608
rect 580814 357856 580870 357912
rect 580630 299104 580686 299160
rect 580354 134816 580410 134872
rect 580722 252184 580778 252240
rect 580814 205264 580870 205320
rect 580906 123120 580962 123176
rect 442262 117952 442318 118008
rect 433522 4800 433578 4856
rect 431222 3304 431278 3360
rect 579802 111424 579858 111480
rect 580170 87896 580226 87952
rect 580170 76200 580226 76256
rect 579802 64504 579858 64560
rect 580170 40976 580226 41032
rect 580170 29280 580226 29336
rect 579802 17584 579858 17640
rect 538126 6160 538182 6216
rect 575018 3304 575074 3360
<< metal3 >>
rect 132166 700436 132172 700500
rect 132236 700498 132242 700500
rect 478505 700498 478571 700501
rect 132236 700496 478571 700498
rect 132236 700440 478510 700496
rect 478566 700440 478571 700496
rect 132236 700438 478571 700440
rect 132236 700436 132242 700438
rect 478505 700435 478571 700438
rect 132350 700300 132356 700364
rect 132420 700362 132426 700364
rect 543457 700362 543523 700365
rect 132420 700360 543523 700362
rect 132420 700304 543462 700360
rect 543518 700304 543523 700360
rect 132420 700302 543523 700304
rect 132420 700300 132426 700302
rect 543457 700299 543523 700302
rect 583520 698050 584960 698140
rect 583342 697990 584960 698050
rect 133638 697172 133644 697236
rect 133708 697234 133714 697236
rect 154481 697234 154547 697237
rect 173801 697234 173867 697237
rect 193121 697234 193187 697237
rect 212441 697234 212507 697237
rect 231761 697234 231827 697237
rect 251081 697234 251147 697237
rect 270401 697234 270467 697237
rect 289721 697234 289787 697237
rect 309041 697234 309107 697237
rect 328361 697234 328427 697237
rect 133708 697174 138122 697234
rect 133708 697172 133714 697174
rect 138062 697098 138122 697174
rect 154481 697232 157442 697234
rect 154481 697176 154486 697232
rect 154542 697176 157442 697232
rect 154481 697174 157442 697176
rect 154481 697171 154547 697174
rect 147581 697098 147647 697101
rect 138062 697096 147647 697098
rect 138062 697040 147586 697096
rect 147642 697040 147647 697096
rect 138062 697038 147647 697040
rect 157382 697098 157442 697174
rect 173801 697232 176762 697234
rect 173801 697176 173806 697232
rect 173862 697176 176762 697232
rect 173801 697174 176762 697176
rect 173801 697171 173867 697174
rect 166901 697098 166967 697101
rect 157382 697096 166967 697098
rect 157382 697040 166906 697096
rect 166962 697040 166967 697096
rect 157382 697038 166967 697040
rect 176702 697098 176762 697174
rect 193121 697232 196082 697234
rect 193121 697176 193126 697232
rect 193182 697176 196082 697232
rect 193121 697174 196082 697176
rect 193121 697171 193187 697174
rect 186221 697098 186287 697101
rect 176702 697096 186287 697098
rect 176702 697040 186226 697096
rect 186282 697040 186287 697096
rect 176702 697038 186287 697040
rect 196022 697098 196082 697174
rect 212441 697232 215402 697234
rect 212441 697176 212446 697232
rect 212502 697176 215402 697232
rect 212441 697174 215402 697176
rect 212441 697171 212507 697174
rect 205541 697098 205607 697101
rect 196022 697096 205607 697098
rect 196022 697040 205546 697096
rect 205602 697040 205607 697096
rect 196022 697038 205607 697040
rect 215342 697098 215402 697174
rect 231761 697232 234722 697234
rect 231761 697176 231766 697232
rect 231822 697176 234722 697232
rect 231761 697174 234722 697176
rect 231761 697171 231827 697174
rect 224861 697098 224927 697101
rect 215342 697096 224927 697098
rect 215342 697040 224866 697096
rect 224922 697040 224927 697096
rect 215342 697038 224927 697040
rect 234662 697098 234722 697174
rect 251081 697232 254042 697234
rect 251081 697176 251086 697232
rect 251142 697176 254042 697232
rect 251081 697174 254042 697176
rect 251081 697171 251147 697174
rect 244181 697098 244247 697101
rect 234662 697096 244247 697098
rect 234662 697040 244186 697096
rect 244242 697040 244247 697096
rect 234662 697038 244247 697040
rect 253982 697098 254042 697174
rect 270401 697232 273362 697234
rect 270401 697176 270406 697232
rect 270462 697176 273362 697232
rect 270401 697174 273362 697176
rect 270401 697171 270467 697174
rect 263501 697098 263567 697101
rect 253982 697096 263567 697098
rect 253982 697040 263506 697096
rect 263562 697040 263567 697096
rect 253982 697038 263567 697040
rect 273302 697098 273362 697174
rect 289721 697232 292682 697234
rect 289721 697176 289726 697232
rect 289782 697176 292682 697232
rect 289721 697174 292682 697176
rect 289721 697171 289787 697174
rect 282821 697098 282887 697101
rect 273302 697096 282887 697098
rect 273302 697040 282826 697096
rect 282882 697040 282887 697096
rect 273302 697038 282887 697040
rect 292622 697098 292682 697174
rect 309041 697232 312002 697234
rect 309041 697176 309046 697232
rect 309102 697176 312002 697232
rect 309041 697174 312002 697176
rect 309041 697171 309107 697174
rect 302141 697098 302207 697101
rect 292622 697096 302207 697098
rect 292622 697040 302146 697096
rect 302202 697040 302207 697096
rect 292622 697038 302207 697040
rect 311942 697098 312002 697174
rect 328361 697232 340890 697234
rect 328361 697176 328366 697232
rect 328422 697176 340890 697232
rect 328361 697174 340890 697176
rect 328361 697171 328427 697174
rect 321461 697098 321527 697101
rect 311942 697096 321527 697098
rect 311942 697040 321466 697096
rect 321522 697040 321527 697096
rect 311942 697038 321527 697040
rect 340830 697098 340890 697174
rect 354630 697174 360210 697234
rect 340830 697038 350458 697098
rect 147581 697035 147647 697038
rect 166901 697035 166967 697038
rect 186221 697035 186287 697038
rect 205541 697035 205607 697038
rect 224861 697035 224927 697038
rect 244181 697035 244247 697038
rect 263501 697035 263567 697038
rect 282821 697035 282887 697038
rect 302141 697035 302207 697038
rect 321461 697035 321527 697038
rect 350398 696962 350458 697038
rect 354630 696962 354690 697174
rect 360150 697098 360210 697174
rect 373950 697174 383578 697234
rect 360150 697038 369778 697098
rect 350398 696902 354690 696962
rect 369718 696962 369778 697038
rect 373950 696962 374010 697174
rect 369718 696902 374010 696962
rect 383518 696962 383578 697174
rect 383702 697174 393330 697234
rect 383702 696962 383762 697174
rect 393270 697098 393330 697174
rect 403022 697174 412650 697234
rect 393270 697038 402898 697098
rect 383518 696902 383762 696962
rect 402838 696962 402898 697038
rect 403022 696962 403082 697174
rect 412590 697098 412650 697174
rect 422342 697174 431970 697234
rect 412590 697038 422218 697098
rect 402838 696902 403082 696962
rect 422158 696962 422218 697038
rect 422342 696962 422402 697174
rect 431910 697098 431970 697174
rect 441662 697174 451290 697234
rect 431910 697038 432154 697098
rect 422158 696902 422402 696962
rect 432094 696962 432154 697038
rect 441662 696962 441722 697174
rect 451230 697098 451290 697174
rect 460982 697174 470610 697234
rect 451230 697038 460858 697098
rect 432094 696902 441722 696962
rect 460798 696962 460858 697038
rect 460982 696962 461042 697174
rect 470550 697098 470610 697174
rect 480302 697174 489930 697234
rect 470550 697038 480178 697098
rect 460798 696902 461042 696962
rect 480118 696962 480178 697038
rect 480302 696962 480362 697174
rect 489870 697098 489930 697174
rect 499622 697174 509250 697234
rect 489870 697038 499498 697098
rect 480118 696902 480362 696962
rect 499438 696962 499498 697038
rect 499622 696962 499682 697174
rect 509190 697098 509250 697174
rect 518942 697174 528570 697234
rect 509190 697038 518818 697098
rect 499438 696902 499682 696962
rect 518758 696962 518818 697038
rect 518942 696962 519002 697174
rect 528510 697098 528570 697174
rect 538262 697174 547890 697234
rect 528510 697038 538138 697098
rect 518758 696902 519002 696962
rect 538078 696962 538138 697038
rect 538262 696962 538322 697174
rect 547830 697098 547890 697174
rect 557582 697174 567210 697234
rect 547830 697038 557458 697098
rect 538078 696902 538322 696962
rect 557398 696962 557458 697038
rect 557582 696962 557642 697174
rect 567150 697098 567210 697174
rect 583342 697098 583402 697990
rect 583520 697900 584960 697990
rect 567150 697038 576778 697098
rect 557398 696902 557642 696962
rect 576718 696962 576778 697038
rect 576902 697038 583402 697098
rect 576902 696962 576962 697038
rect 576718 696902 576962 696962
rect -960 696540 480 696780
rect 164182 686428 164188 686492
rect 164252 686490 164258 686492
rect 169017 686490 169083 686493
rect 164252 686488 169083 686490
rect 164252 686432 169022 686488
rect 169078 686432 169083 686488
rect 164252 686430 169083 686432
rect 164252 686428 164258 686430
rect 169017 686427 169083 686430
rect 147765 686354 147831 686357
rect 154573 686354 154639 686357
rect 583520 686354 584960 686444
rect 147765 686352 154639 686354
rect 147765 686296 147770 686352
rect 147826 686296 154578 686352
rect 154634 686296 154639 686352
rect 147765 686294 154639 686296
rect 147765 686291 147831 686294
rect 154573 686291 154639 686294
rect 583342 686294 584960 686354
rect 135253 686218 135319 686221
rect 132542 686216 135319 686218
rect 132542 686160 135258 686216
rect 135314 686160 135319 686216
rect 132542 686158 135319 686160
rect 131982 685884 131988 685948
rect 132052 685946 132058 685948
rect 132542 685946 132602 686158
rect 135253 686155 135319 686158
rect 159449 686218 159515 686221
rect 164182 686218 164188 686220
rect 159449 686216 164188 686218
rect 159449 686160 159454 686216
rect 159510 686160 164188 686216
rect 159449 686158 164188 686160
rect 159449 686155 159515 686158
rect 164182 686156 164188 686158
rect 164252 686156 164258 686220
rect 169017 686218 169083 686221
rect 169017 686216 180810 686218
rect 169017 686160 169022 686216
rect 169078 686160 180810 686216
rect 169017 686158 180810 686160
rect 169017 686155 169083 686158
rect 147581 686082 147647 686085
rect 144870 686080 147647 686082
rect 144870 686024 147586 686080
rect 147642 686024 147647 686080
rect 144870 686022 147647 686024
rect 180750 686082 180810 686158
rect 190502 686158 200130 686218
rect 180750 686022 190378 686082
rect 132052 685886 132602 685946
rect 142889 685946 142955 685949
rect 144870 685946 144930 686022
rect 147581 686019 147647 686022
rect 142889 685944 144930 685946
rect 142889 685888 142894 685944
rect 142950 685888 144930 685944
rect 142889 685886 144930 685888
rect 190318 685946 190378 686022
rect 190502 685946 190562 686158
rect 200070 686082 200130 686158
rect 209822 686158 219450 686218
rect 200070 686022 209698 686082
rect 190318 685886 190562 685946
rect 209638 685946 209698 686022
rect 209822 685946 209882 686158
rect 219390 686082 219450 686158
rect 229142 686158 238770 686218
rect 219390 686022 229018 686082
rect 209638 685886 209882 685946
rect 228958 685946 229018 686022
rect 229142 685946 229202 686158
rect 238710 686082 238770 686158
rect 248462 686158 258090 686218
rect 238710 686022 248338 686082
rect 228958 685886 229202 685946
rect 248278 685946 248338 686022
rect 248462 685946 248522 686158
rect 258030 686082 258090 686158
rect 267782 686158 277410 686218
rect 258030 686022 267658 686082
rect 248278 685886 248522 685946
rect 267598 685946 267658 686022
rect 267782 685946 267842 686158
rect 277350 686082 277410 686158
rect 287102 686158 296730 686218
rect 277350 686022 286978 686082
rect 267598 685886 267842 685946
rect 286918 685946 286978 686022
rect 287102 685946 287162 686158
rect 296670 686082 296730 686158
rect 306422 686158 316050 686218
rect 296670 686022 306298 686082
rect 286918 685886 287162 685946
rect 306238 685946 306298 686022
rect 306422 685946 306482 686158
rect 315990 686082 316050 686158
rect 325742 686158 335370 686218
rect 315990 686022 325618 686082
rect 306238 685886 306482 685946
rect 325558 685946 325618 686022
rect 325742 685946 325802 686158
rect 335310 686082 335370 686158
rect 345062 686158 354690 686218
rect 335310 686022 344938 686082
rect 325558 685886 325802 685946
rect 344878 685946 344938 686022
rect 345062 685946 345122 686158
rect 354630 686082 354690 686158
rect 364382 686158 374010 686218
rect 354630 686022 364258 686082
rect 344878 685886 345122 685946
rect 364198 685946 364258 686022
rect 364382 685946 364442 686158
rect 373950 686082 374010 686158
rect 383702 686158 393330 686218
rect 373950 686022 383578 686082
rect 364198 685886 364442 685946
rect 383518 685946 383578 686022
rect 383702 685946 383762 686158
rect 393270 686082 393330 686158
rect 403022 686158 412650 686218
rect 393270 686022 402898 686082
rect 383518 685886 383762 685946
rect 402838 685946 402898 686022
rect 403022 685946 403082 686158
rect 412590 686082 412650 686158
rect 422342 686158 431970 686218
rect 412590 686022 422218 686082
rect 402838 685886 403082 685946
rect 422158 685946 422218 686022
rect 422342 685946 422402 686158
rect 431910 686082 431970 686158
rect 441662 686158 451290 686218
rect 431910 686022 441538 686082
rect 422158 685886 422402 685946
rect 441478 685946 441538 686022
rect 441662 685946 441722 686158
rect 451230 686082 451290 686158
rect 460982 686158 470610 686218
rect 451230 686022 460858 686082
rect 441478 685886 441722 685946
rect 460798 685946 460858 686022
rect 460982 685946 461042 686158
rect 470550 686082 470610 686158
rect 480302 686158 489930 686218
rect 470550 686022 480178 686082
rect 460798 685886 461042 685946
rect 480118 685946 480178 686022
rect 480302 685946 480362 686158
rect 489870 686082 489930 686158
rect 499622 686158 509250 686218
rect 489870 686022 499498 686082
rect 480118 685886 480362 685946
rect 499438 685946 499498 686022
rect 499622 685946 499682 686158
rect 509190 686082 509250 686158
rect 518942 686158 528570 686218
rect 509190 686022 518818 686082
rect 499438 685886 499682 685946
rect 518758 685946 518818 686022
rect 518942 685946 519002 686158
rect 528510 686082 528570 686158
rect 538262 686158 547890 686218
rect 528510 686022 538138 686082
rect 518758 685886 519002 685946
rect 538078 685946 538138 686022
rect 538262 685946 538322 686158
rect 547830 686082 547890 686158
rect 557582 686158 567210 686218
rect 547830 686022 557458 686082
rect 538078 685886 538322 685946
rect 557398 685946 557458 686022
rect 557582 685946 557642 686158
rect 567150 686082 567210 686158
rect 583342 686082 583402 686294
rect 583520 686204 584960 686294
rect 567150 686022 576778 686082
rect 557398 685886 557642 685946
rect 576718 685946 576778 686022
rect 576902 686022 583402 686082
rect 576902 685946 576962 686022
rect 576718 685886 576962 685946
rect 132052 685884 132058 685886
rect 142889 685883 142955 685886
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 4797 653578 4863 653581
rect -960 653576 4863 653578
rect -960 653520 4802 653576
rect 4858 653520 4863 653576
rect -960 653518 4863 653520
rect -960 653428 480 653518
rect 4797 653515 4863 653518
rect 583520 651130 584960 651220
rect 583342 651070 584960 651130
rect 164182 650524 164188 650588
rect 164252 650586 164258 650588
rect 169017 650586 169083 650589
rect 164252 650584 169083 650586
rect 164252 650528 169022 650584
rect 169078 650528 169083 650584
rect 164252 650526 169083 650528
rect 164252 650524 164258 650526
rect 169017 650523 169083 650526
rect 147765 650450 147831 650453
rect 154573 650450 154639 650453
rect 147765 650448 154639 650450
rect 147765 650392 147770 650448
rect 147826 650392 154578 650448
rect 154634 650392 154639 650448
rect 147765 650390 154639 650392
rect 147765 650387 147831 650390
rect 154573 650387 154639 650390
rect 133454 650252 133460 650316
rect 133524 650314 133530 650316
rect 135253 650314 135319 650317
rect 133524 650312 135319 650314
rect 133524 650256 135258 650312
rect 135314 650256 135319 650312
rect 133524 650254 135319 650256
rect 133524 650252 133530 650254
rect 135253 650251 135319 650254
rect 159449 650314 159515 650317
rect 164182 650314 164188 650316
rect 159449 650312 164188 650314
rect 159449 650256 159454 650312
rect 159510 650256 164188 650312
rect 159449 650254 164188 650256
rect 159449 650251 159515 650254
rect 164182 650252 164188 650254
rect 164252 650252 164258 650316
rect 169017 650314 169083 650317
rect 169017 650312 180810 650314
rect 169017 650256 169022 650312
rect 169078 650256 180810 650312
rect 169017 650254 180810 650256
rect 169017 650251 169083 650254
rect 147581 650178 147647 650181
rect 144870 650176 147647 650178
rect 144870 650120 147586 650176
rect 147642 650120 147647 650176
rect 144870 650118 147647 650120
rect 180750 650178 180810 650254
rect 190502 650254 200130 650314
rect 180750 650118 190378 650178
rect 142889 650042 142955 650045
rect 144870 650042 144930 650118
rect 147581 650115 147647 650118
rect 142889 650040 144930 650042
rect 142889 649984 142894 650040
rect 142950 649984 144930 650040
rect 142889 649982 144930 649984
rect 190318 650042 190378 650118
rect 190502 650042 190562 650254
rect 200070 650178 200130 650254
rect 209822 650254 219450 650314
rect 200070 650118 209698 650178
rect 190318 649982 190562 650042
rect 209638 650042 209698 650118
rect 209822 650042 209882 650254
rect 219390 650178 219450 650254
rect 229142 650254 238770 650314
rect 219390 650118 229018 650178
rect 209638 649982 209882 650042
rect 228958 650042 229018 650118
rect 229142 650042 229202 650254
rect 238710 650178 238770 650254
rect 248462 650254 258090 650314
rect 238710 650118 248338 650178
rect 228958 649982 229202 650042
rect 248278 650042 248338 650118
rect 248462 650042 248522 650254
rect 258030 650178 258090 650254
rect 267782 650254 277410 650314
rect 258030 650118 267658 650178
rect 248278 649982 248522 650042
rect 267598 650042 267658 650118
rect 267782 650042 267842 650254
rect 277350 650178 277410 650254
rect 287102 650254 296730 650314
rect 277350 650118 286978 650178
rect 267598 649982 267842 650042
rect 286918 650042 286978 650118
rect 287102 650042 287162 650254
rect 296670 650178 296730 650254
rect 306422 650254 316050 650314
rect 296670 650118 306298 650178
rect 286918 649982 287162 650042
rect 306238 650042 306298 650118
rect 306422 650042 306482 650254
rect 315990 650178 316050 650254
rect 325742 650254 335370 650314
rect 315990 650118 325618 650178
rect 306238 649982 306482 650042
rect 325558 650042 325618 650118
rect 325742 650042 325802 650254
rect 335310 650178 335370 650254
rect 345062 650254 354690 650314
rect 335310 650118 344938 650178
rect 325558 649982 325802 650042
rect 344878 650042 344938 650118
rect 345062 650042 345122 650254
rect 354630 650178 354690 650254
rect 364382 650254 374010 650314
rect 354630 650118 364258 650178
rect 344878 649982 345122 650042
rect 364198 650042 364258 650118
rect 364382 650042 364442 650254
rect 373950 650178 374010 650254
rect 383702 650254 393330 650314
rect 373950 650118 383578 650178
rect 364198 649982 364442 650042
rect 383518 650042 383578 650118
rect 383702 650042 383762 650254
rect 393270 650178 393330 650254
rect 403022 650254 412650 650314
rect 393270 650118 402898 650178
rect 383518 649982 383762 650042
rect 402838 650042 402898 650118
rect 403022 650042 403082 650254
rect 412590 650178 412650 650254
rect 422342 650254 431970 650314
rect 412590 650118 422218 650178
rect 402838 649982 403082 650042
rect 422158 650042 422218 650118
rect 422342 650042 422402 650254
rect 431910 650178 431970 650254
rect 441662 650254 451290 650314
rect 431910 650118 441538 650178
rect 422158 649982 422402 650042
rect 441478 650042 441538 650118
rect 441662 650042 441722 650254
rect 451230 650178 451290 650254
rect 460982 650254 470610 650314
rect 451230 650118 460858 650178
rect 441478 649982 441722 650042
rect 460798 650042 460858 650118
rect 460982 650042 461042 650254
rect 470550 650178 470610 650254
rect 480302 650254 489930 650314
rect 470550 650118 480178 650178
rect 460798 649982 461042 650042
rect 480118 650042 480178 650118
rect 480302 650042 480362 650254
rect 489870 650178 489930 650254
rect 499622 650254 509250 650314
rect 489870 650118 499498 650178
rect 480118 649982 480362 650042
rect 499438 650042 499498 650118
rect 499622 650042 499682 650254
rect 509190 650178 509250 650254
rect 518942 650254 528570 650314
rect 509190 650118 518818 650178
rect 499438 649982 499682 650042
rect 518758 650042 518818 650118
rect 518942 650042 519002 650254
rect 528510 650178 528570 650254
rect 538262 650254 547890 650314
rect 528510 650118 538138 650178
rect 518758 649982 519002 650042
rect 538078 650042 538138 650118
rect 538262 650042 538322 650254
rect 547830 650178 547890 650254
rect 557582 650254 567210 650314
rect 547830 650118 557458 650178
rect 538078 649982 538322 650042
rect 557398 650042 557458 650118
rect 557582 650042 557642 650254
rect 567150 650178 567210 650254
rect 583342 650178 583402 651070
rect 583520 650980 584960 651070
rect 567150 650118 576778 650178
rect 557398 649982 557642 650042
rect 576718 650042 576778 650118
rect 576902 650118 583402 650178
rect 576902 650042 576962 650118
rect 576718 649982 576962 650042
rect 142889 649979 142955 649982
rect 583520 639434 584960 639524
rect 583342 639374 584960 639434
rect 157057 639298 157123 639301
rect 132542 639296 157123 639298
rect -960 639012 480 639252
rect 132542 639240 157062 639296
rect 157118 639240 157123 639296
rect 132542 639238 157123 639240
rect 131798 638964 131804 639028
rect 131868 639026 131874 639028
rect 132542 639026 132602 639238
rect 157057 639235 157123 639238
rect 157241 639298 157307 639301
rect 171041 639298 171107 639301
rect 157241 639296 159282 639298
rect 157241 639240 157246 639296
rect 157302 639240 159282 639296
rect 157241 639238 159282 639240
rect 157241 639235 157307 639238
rect 159222 639162 159282 639238
rect 171041 639296 180810 639298
rect 171041 639240 171046 639296
rect 171102 639240 180810 639296
rect 171041 639238 180810 639240
rect 171041 639235 171107 639238
rect 164182 639162 164188 639164
rect 159222 639102 164188 639162
rect 164182 639100 164188 639102
rect 164252 639100 164258 639164
rect 180750 639162 180810 639238
rect 190502 639238 200130 639298
rect 180750 639102 190378 639162
rect 131868 638966 132602 639026
rect 190318 639026 190378 639102
rect 190502 639026 190562 639238
rect 200070 639162 200130 639238
rect 209822 639238 219450 639298
rect 200070 639102 209698 639162
rect 190318 638966 190562 639026
rect 209638 639026 209698 639102
rect 209822 639026 209882 639238
rect 219390 639162 219450 639238
rect 229142 639238 238770 639298
rect 219390 639102 229018 639162
rect 209638 638966 209882 639026
rect 228958 639026 229018 639102
rect 229142 639026 229202 639238
rect 238710 639162 238770 639238
rect 248462 639238 258090 639298
rect 238710 639102 248338 639162
rect 228958 638966 229202 639026
rect 248278 639026 248338 639102
rect 248462 639026 248522 639238
rect 258030 639162 258090 639238
rect 267782 639238 277410 639298
rect 258030 639102 267658 639162
rect 248278 638966 248522 639026
rect 267598 639026 267658 639102
rect 267782 639026 267842 639238
rect 277350 639162 277410 639238
rect 287102 639238 296730 639298
rect 277350 639102 286978 639162
rect 267598 638966 267842 639026
rect 286918 639026 286978 639102
rect 287102 639026 287162 639238
rect 296670 639162 296730 639238
rect 306422 639238 316050 639298
rect 296670 639102 306298 639162
rect 286918 638966 287162 639026
rect 306238 639026 306298 639102
rect 306422 639026 306482 639238
rect 315990 639162 316050 639238
rect 325742 639238 335370 639298
rect 315990 639102 325618 639162
rect 306238 638966 306482 639026
rect 325558 639026 325618 639102
rect 325742 639026 325802 639238
rect 335310 639162 335370 639238
rect 345062 639238 354690 639298
rect 335310 639102 344938 639162
rect 325558 638966 325802 639026
rect 344878 639026 344938 639102
rect 345062 639026 345122 639238
rect 354630 639162 354690 639238
rect 364382 639238 374010 639298
rect 354630 639102 364258 639162
rect 344878 638966 345122 639026
rect 364198 639026 364258 639102
rect 364382 639026 364442 639238
rect 373950 639162 374010 639238
rect 383702 639238 393330 639298
rect 373950 639102 383578 639162
rect 364198 638966 364442 639026
rect 383518 639026 383578 639102
rect 383702 639026 383762 639238
rect 393270 639162 393330 639238
rect 403022 639238 412650 639298
rect 393270 639102 402898 639162
rect 383518 638966 383762 639026
rect 402838 639026 402898 639102
rect 403022 639026 403082 639238
rect 412590 639162 412650 639238
rect 422342 639238 431970 639298
rect 412590 639102 422218 639162
rect 402838 638966 403082 639026
rect 422158 639026 422218 639102
rect 422342 639026 422402 639238
rect 431910 639162 431970 639238
rect 441662 639238 451290 639298
rect 431910 639102 441538 639162
rect 422158 638966 422402 639026
rect 441478 639026 441538 639102
rect 441662 639026 441722 639238
rect 451230 639162 451290 639238
rect 460982 639238 470610 639298
rect 451230 639102 460858 639162
rect 441478 638966 441722 639026
rect 460798 639026 460858 639102
rect 460982 639026 461042 639238
rect 470550 639162 470610 639238
rect 480302 639238 489930 639298
rect 470550 639102 480178 639162
rect 460798 638966 461042 639026
rect 480118 639026 480178 639102
rect 480302 639026 480362 639238
rect 489870 639162 489930 639238
rect 499622 639238 509250 639298
rect 489870 639102 499498 639162
rect 480118 638966 480362 639026
rect 499438 639026 499498 639102
rect 499622 639026 499682 639238
rect 509190 639162 509250 639238
rect 518942 639238 528570 639298
rect 509190 639102 518818 639162
rect 499438 638966 499682 639026
rect 518758 639026 518818 639102
rect 518942 639026 519002 639238
rect 528510 639162 528570 639238
rect 538262 639238 547890 639298
rect 528510 639102 538138 639162
rect 518758 638966 519002 639026
rect 538078 639026 538138 639102
rect 538262 639026 538322 639238
rect 547830 639162 547890 639238
rect 557582 639238 567210 639298
rect 547830 639102 557458 639162
rect 538078 638966 538322 639026
rect 557398 639026 557458 639102
rect 557582 639026 557642 639238
rect 567150 639162 567210 639238
rect 583342 639162 583402 639374
rect 583520 639284 584960 639374
rect 567150 639102 576778 639162
rect 557398 638966 557642 639026
rect 576718 639026 576778 639102
rect 576902 639102 583402 639162
rect 576902 639026 576962 639102
rect 576718 638966 576962 639026
rect 131868 638964 131874 638966
rect 164182 638828 164188 638892
rect 164252 638890 164258 638892
rect 171041 638890 171107 638893
rect 164252 638888 171107 638890
rect 164252 638832 171046 638888
rect 171102 638832 171107 638888
rect 164252 638830 171107 638832
rect 164252 638828 164258 638830
rect 171041 638827 171107 638830
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3417 624882 3483 624885
rect -960 624880 3483 624882
rect -960 624824 3422 624880
rect 3478 624824 3483 624880
rect -960 624822 3483 624824
rect -960 624732 480 624822
rect 3417 624819 3483 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 583520 604210 584960 604300
rect 583342 604150 584960 604210
rect 133086 603332 133092 603396
rect 133156 603394 133162 603396
rect 157057 603394 157123 603397
rect 133156 603392 157123 603394
rect 133156 603336 157062 603392
rect 157118 603336 157123 603392
rect 133156 603334 157123 603336
rect 133156 603332 133162 603334
rect 157057 603331 157123 603334
rect 157241 603394 157307 603397
rect 171041 603394 171107 603397
rect 157241 603392 159466 603394
rect 157241 603336 157246 603392
rect 157302 603336 159466 603392
rect 157241 603334 159466 603336
rect 157241 603331 157307 603334
rect 159406 603258 159466 603334
rect 171041 603392 180810 603394
rect 171041 603336 171046 603392
rect 171102 603336 180810 603392
rect 171041 603334 180810 603336
rect 171041 603331 171107 603334
rect 164182 603258 164188 603260
rect 159406 603198 164188 603258
rect 164182 603196 164188 603198
rect 164252 603196 164258 603260
rect 180750 603258 180810 603334
rect 190502 603334 200130 603394
rect 180750 603198 190378 603258
rect 190318 603122 190378 603198
rect 190502 603122 190562 603334
rect 200070 603258 200130 603334
rect 209822 603334 219450 603394
rect 200070 603198 209698 603258
rect 190318 603062 190562 603122
rect 209638 603122 209698 603198
rect 209822 603122 209882 603334
rect 219390 603258 219450 603334
rect 229142 603334 238770 603394
rect 219390 603198 229018 603258
rect 209638 603062 209882 603122
rect 228958 603122 229018 603198
rect 229142 603122 229202 603334
rect 238710 603258 238770 603334
rect 248462 603334 258090 603394
rect 238710 603198 248338 603258
rect 228958 603062 229202 603122
rect 248278 603122 248338 603198
rect 248462 603122 248522 603334
rect 258030 603258 258090 603334
rect 267782 603334 277410 603394
rect 258030 603198 267658 603258
rect 248278 603062 248522 603122
rect 267598 603122 267658 603198
rect 267782 603122 267842 603334
rect 277350 603258 277410 603334
rect 287102 603334 296730 603394
rect 277350 603198 286978 603258
rect 267598 603062 267842 603122
rect 286918 603122 286978 603198
rect 287102 603122 287162 603334
rect 296670 603258 296730 603334
rect 306422 603334 316050 603394
rect 296670 603198 306298 603258
rect 286918 603062 287162 603122
rect 306238 603122 306298 603198
rect 306422 603122 306482 603334
rect 315990 603258 316050 603334
rect 325742 603334 335370 603394
rect 315990 603198 325618 603258
rect 306238 603062 306482 603122
rect 325558 603122 325618 603198
rect 325742 603122 325802 603334
rect 335310 603258 335370 603334
rect 345062 603334 354690 603394
rect 335310 603198 344938 603258
rect 325558 603062 325802 603122
rect 344878 603122 344938 603198
rect 345062 603122 345122 603334
rect 354630 603258 354690 603334
rect 364382 603334 374010 603394
rect 354630 603198 364258 603258
rect 344878 603062 345122 603122
rect 364198 603122 364258 603198
rect 364382 603122 364442 603334
rect 373950 603258 374010 603334
rect 383702 603334 393330 603394
rect 373950 603198 383578 603258
rect 364198 603062 364442 603122
rect 383518 603122 383578 603198
rect 383702 603122 383762 603334
rect 393270 603258 393330 603334
rect 403022 603334 412650 603394
rect 393270 603198 402898 603258
rect 383518 603062 383762 603122
rect 402838 603122 402898 603198
rect 403022 603122 403082 603334
rect 412590 603258 412650 603334
rect 422342 603334 431970 603394
rect 412590 603198 422218 603258
rect 402838 603062 403082 603122
rect 422158 603122 422218 603198
rect 422342 603122 422402 603334
rect 431910 603258 431970 603334
rect 441662 603334 451290 603394
rect 431910 603198 441538 603258
rect 422158 603062 422402 603122
rect 441478 603122 441538 603198
rect 441662 603122 441722 603334
rect 451230 603258 451290 603334
rect 460982 603334 470610 603394
rect 451230 603198 460858 603258
rect 441478 603062 441722 603122
rect 460798 603122 460858 603198
rect 460982 603122 461042 603334
rect 470550 603258 470610 603334
rect 480302 603334 489930 603394
rect 470550 603198 480178 603258
rect 460798 603062 461042 603122
rect 480118 603122 480178 603198
rect 480302 603122 480362 603334
rect 489870 603258 489930 603334
rect 499622 603334 509250 603394
rect 489870 603198 499498 603258
rect 480118 603062 480362 603122
rect 499438 603122 499498 603198
rect 499622 603122 499682 603334
rect 509190 603258 509250 603334
rect 518942 603334 528570 603394
rect 509190 603198 518818 603258
rect 499438 603062 499682 603122
rect 518758 603122 518818 603198
rect 518942 603122 519002 603334
rect 528510 603258 528570 603334
rect 538262 603334 547890 603394
rect 528510 603198 538138 603258
rect 518758 603062 519002 603122
rect 538078 603122 538138 603198
rect 538262 603122 538322 603334
rect 547830 603258 547890 603334
rect 557582 603334 567210 603394
rect 547830 603198 557458 603258
rect 538078 603062 538322 603122
rect 557398 603122 557458 603198
rect 557582 603122 557642 603334
rect 567150 603258 567210 603334
rect 583342 603258 583402 604150
rect 583520 604060 584960 604150
rect 567150 603198 576778 603258
rect 557398 603062 557642 603122
rect 576718 603122 576778 603198
rect 576902 603198 583402 603258
rect 576902 603122 576962 603198
rect 576718 603062 576962 603122
rect 164182 602924 164188 602988
rect 164252 602986 164258 602988
rect 171041 602986 171107 602989
rect 164252 602984 171107 602986
rect 164252 602928 171046 602984
rect 171102 602928 171107 602984
rect 164252 602926 171107 602928
rect 164252 602924 164258 602926
rect 171041 602923 171107 602926
rect 153377 598906 153443 598909
rect 153561 598906 153627 598909
rect 153377 598904 153627 598906
rect 153377 598848 153382 598904
rect 153438 598848 153566 598904
rect 153622 598848 153627 598904
rect 153377 598846 153627 598848
rect 153377 598843 153443 598846
rect 153561 598843 153627 598846
rect -960 596050 480 596140
rect 4061 596050 4127 596053
rect -960 596048 4127 596050
rect -960 595992 4066 596048
rect 4122 595992 4127 596048
rect -960 595990 4127 595992
rect -960 595900 480 595990
rect 4061 595987 4127 595990
rect 583520 592514 584960 592604
rect 583342 592454 584960 592514
rect 133270 592316 133276 592380
rect 133340 592378 133346 592380
rect 157057 592378 157123 592381
rect 133340 592376 157123 592378
rect 133340 592320 157062 592376
rect 157118 592320 157123 592376
rect 133340 592318 157123 592320
rect 133340 592316 133346 592318
rect 157057 592315 157123 592318
rect 157241 592378 157307 592381
rect 171041 592378 171107 592381
rect 157241 592376 159282 592378
rect 157241 592320 157246 592376
rect 157302 592320 159282 592376
rect 157241 592318 159282 592320
rect 157241 592315 157307 592318
rect 159222 592242 159282 592318
rect 171041 592376 180810 592378
rect 171041 592320 171046 592376
rect 171102 592320 180810 592376
rect 171041 592318 180810 592320
rect 171041 592315 171107 592318
rect 164182 592242 164188 592244
rect 159222 592182 164188 592242
rect 164182 592180 164188 592182
rect 164252 592180 164258 592244
rect 180750 592242 180810 592318
rect 190502 592318 200130 592378
rect 180750 592182 190378 592242
rect 190318 592106 190378 592182
rect 190502 592106 190562 592318
rect 200070 592242 200130 592318
rect 209822 592318 219450 592378
rect 200070 592182 209698 592242
rect 190318 592046 190562 592106
rect 209638 592106 209698 592182
rect 209822 592106 209882 592318
rect 219390 592242 219450 592318
rect 229142 592318 238770 592378
rect 219390 592182 229018 592242
rect 209638 592046 209882 592106
rect 228958 592106 229018 592182
rect 229142 592106 229202 592318
rect 238710 592242 238770 592318
rect 248462 592318 258090 592378
rect 238710 592182 248338 592242
rect 228958 592046 229202 592106
rect 248278 592106 248338 592182
rect 248462 592106 248522 592318
rect 258030 592242 258090 592318
rect 267782 592318 277410 592378
rect 258030 592182 267658 592242
rect 248278 592046 248522 592106
rect 267598 592106 267658 592182
rect 267782 592106 267842 592318
rect 277350 592242 277410 592318
rect 287102 592318 296730 592378
rect 277350 592182 286978 592242
rect 267598 592046 267842 592106
rect 286918 592106 286978 592182
rect 287102 592106 287162 592318
rect 296670 592242 296730 592318
rect 306422 592318 316050 592378
rect 296670 592182 306298 592242
rect 286918 592046 287162 592106
rect 306238 592106 306298 592182
rect 306422 592106 306482 592318
rect 315990 592242 316050 592318
rect 325742 592318 335370 592378
rect 315990 592182 325618 592242
rect 306238 592046 306482 592106
rect 325558 592106 325618 592182
rect 325742 592106 325802 592318
rect 335310 592242 335370 592318
rect 345062 592318 354690 592378
rect 335310 592182 344938 592242
rect 325558 592046 325802 592106
rect 344878 592106 344938 592182
rect 345062 592106 345122 592318
rect 354630 592242 354690 592318
rect 364382 592318 374010 592378
rect 354630 592182 364258 592242
rect 344878 592046 345122 592106
rect 364198 592106 364258 592182
rect 364382 592106 364442 592318
rect 373950 592242 374010 592318
rect 383702 592318 393330 592378
rect 373950 592182 383578 592242
rect 364198 592046 364442 592106
rect 383518 592106 383578 592182
rect 383702 592106 383762 592318
rect 393270 592242 393330 592318
rect 403022 592318 412650 592378
rect 393270 592182 402898 592242
rect 383518 592046 383762 592106
rect 402838 592106 402898 592182
rect 403022 592106 403082 592318
rect 412590 592242 412650 592318
rect 422342 592318 431970 592378
rect 412590 592182 422218 592242
rect 402838 592046 403082 592106
rect 422158 592106 422218 592182
rect 422342 592106 422402 592318
rect 431910 592242 431970 592318
rect 441662 592318 451290 592378
rect 431910 592182 441538 592242
rect 422158 592046 422402 592106
rect 441478 592106 441538 592182
rect 441662 592106 441722 592318
rect 451230 592242 451290 592318
rect 460982 592318 470610 592378
rect 451230 592182 460858 592242
rect 441478 592046 441722 592106
rect 460798 592106 460858 592182
rect 460982 592106 461042 592318
rect 470550 592242 470610 592318
rect 480302 592318 489930 592378
rect 470550 592182 480178 592242
rect 460798 592046 461042 592106
rect 480118 592106 480178 592182
rect 480302 592106 480362 592318
rect 489870 592242 489930 592318
rect 499622 592318 509250 592378
rect 489870 592182 499498 592242
rect 480118 592046 480362 592106
rect 499438 592106 499498 592182
rect 499622 592106 499682 592318
rect 509190 592242 509250 592318
rect 518942 592318 528570 592378
rect 509190 592182 518818 592242
rect 499438 592046 499682 592106
rect 518758 592106 518818 592182
rect 518942 592106 519002 592318
rect 528510 592242 528570 592318
rect 538262 592318 547890 592378
rect 528510 592182 538138 592242
rect 518758 592046 519002 592106
rect 538078 592106 538138 592182
rect 538262 592106 538322 592318
rect 547830 592242 547890 592318
rect 557582 592318 567210 592378
rect 547830 592182 557458 592242
rect 538078 592046 538322 592106
rect 557398 592106 557458 592182
rect 557582 592106 557642 592318
rect 567150 592242 567210 592318
rect 583342 592242 583402 592454
rect 583520 592364 584960 592454
rect 567150 592182 576778 592242
rect 557398 592046 557642 592106
rect 576718 592106 576778 592182
rect 576902 592182 583402 592242
rect 576902 592106 576962 592182
rect 576718 592046 576962 592106
rect 164182 591908 164188 591972
rect 164252 591970 164258 591972
rect 171041 591970 171107 591973
rect 164252 591968 171107 591970
rect 164252 591912 171046 591968
rect 171102 591912 171107 591968
rect 164252 591910 171107 591912
rect 164252 591908 164258 591910
rect 171041 591907 171107 591910
rect 274541 582586 274607 582589
rect 368657 582586 368723 582589
rect 274541 582584 368723 582586
rect 274541 582528 274546 582584
rect 274602 582528 368662 582584
rect 368718 582528 368723 582584
rect 274541 582526 368723 582528
rect 274541 582523 274607 582526
rect 368657 582523 368723 582526
rect 129641 582450 129707 582453
rect 349521 582450 349587 582453
rect 129641 582448 349587 582450
rect 129641 582392 129646 582448
rect 129702 582392 349526 582448
rect 349582 582392 349587 582448
rect 129641 582390 349587 582392
rect 129641 582387 129707 582390
rect 349521 582387 349587 582390
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 296713 575786 296779 575789
rect 299982 575786 300042 576232
rect 296713 575784 300042 575786
rect 296713 575728 296718 575784
rect 296774 575728 300042 575784
rect 296713 575726 300042 575728
rect 296713 575723 296779 575726
rect 377814 575514 377874 575960
rect 380617 575514 380683 575517
rect 377814 575512 380683 575514
rect 377814 575456 380622 575512
rect 380678 575456 380683 575512
rect 377814 575454 380683 575456
rect 380617 575451 380683 575454
rect 297449 572930 297515 572933
rect 299982 572930 300042 572968
rect 297449 572928 300042 572930
rect 297449 572872 297454 572928
rect 297510 572872 300042 572928
rect 297449 572870 300042 572872
rect 297449 572867 297515 572870
rect 377814 572114 377874 572696
rect 379462 572114 379468 572116
rect 377814 572054 379468 572114
rect 379462 572052 379468 572054
rect 379532 572052 379538 572116
rect 298001 570074 298067 570077
rect 298001 570072 300042 570074
rect 298001 570016 298006 570072
rect 298062 570016 300042 570072
rect 298001 570014 300042 570016
rect 298001 570011 298067 570014
rect 299982 569976 300042 570014
rect 377814 569122 377874 569704
rect 379513 569122 379579 569125
rect 377814 569120 379579 569122
rect 377814 569064 379518 569120
rect 379574 569064 379579 569120
rect 377814 569062 379579 569064
rect 379513 569059 379579 569062
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3417 567354 3483 567357
rect -960 567352 3483 567354
rect -960 567296 3422 567352
rect 3478 567296 3483 567352
rect -960 567294 3483 567296
rect -960 567204 480 567294
rect 3417 567291 3483 567294
rect 296437 565858 296503 565861
rect 299982 565858 300042 566712
rect 296437 565856 300042 565858
rect 296437 565800 296442 565856
rect 296498 565800 300042 565856
rect 296437 565798 300042 565800
rect 377262 565861 377322 566440
rect 377262 565856 377371 565861
rect 377262 565800 377310 565856
rect 377366 565800 377371 565856
rect 377262 565798 377371 565800
rect 296437 565795 296503 565798
rect 377305 565795 377371 565798
rect 296897 563410 296963 563413
rect 299982 563410 300042 563720
rect 296897 563408 300042 563410
rect 296897 563352 296902 563408
rect 296958 563352 300042 563408
rect 296897 563350 300042 563352
rect 296897 563347 296963 563350
rect 377446 563141 377506 563448
rect 377397 563136 377506 563141
rect 377397 563080 377402 563136
rect 377458 563080 377506 563136
rect 377397 563078 377506 563080
rect 377397 563075 377463 563078
rect 199694 561716 199700 561780
rect 199764 561778 199770 561780
rect 211613 561778 211679 561781
rect 199764 561776 211679 561778
rect 199764 561720 211618 561776
rect 211674 561720 211679 561776
rect 199764 561718 211679 561720
rect 199764 561716 199770 561718
rect 211613 561715 211679 561718
rect 298001 560418 298067 560421
rect 299982 560418 300042 560456
rect 298001 560416 300042 560418
rect 298001 560360 298006 560416
rect 298062 560360 300042 560416
rect 298001 560358 300042 560360
rect 298001 560355 298067 560358
rect 378133 560214 378199 560217
rect 377844 560212 378199 560214
rect 377844 560156 378138 560212
rect 378194 560156 378199 560212
rect 377844 560154 378199 560156
rect 378133 560151 378199 560154
rect 198590 556684 198596 556748
rect 198660 556746 198666 556748
rect 200070 556746 200130 557328
rect 297081 556882 297147 556885
rect 299982 556882 300042 557464
rect 580257 557290 580323 557293
rect 583520 557290 584960 557380
rect 580257 557288 584960 557290
rect 580257 557232 580262 557288
rect 580318 557232 584960 557288
rect 580257 557230 584960 557232
rect 580257 557227 580323 557230
rect 297081 556880 300042 556882
rect 297081 556824 297086 556880
rect 297142 556824 300042 556880
rect 297081 556822 300042 556824
rect 297081 556819 297147 556822
rect 198660 556686 200130 556746
rect 198660 556684 198666 556686
rect 219942 556202 220002 556784
rect 377446 556613 377506 557192
rect 583520 557140 584960 557230
rect 377446 556608 377555 556613
rect 377446 556552 377494 556608
rect 377550 556552 377555 556608
rect 377446 556550 377555 556552
rect 377489 556547 377555 556550
rect 222193 556202 222259 556205
rect 219942 556200 222259 556202
rect 219942 556144 222198 556200
rect 222254 556144 222259 556200
rect 219942 556142 222259 556144
rect 222193 556139 222259 556142
rect 297909 553618 297975 553621
rect 299982 553618 300042 554200
rect 297909 553616 300042 553618
rect 297909 553560 297914 553616
rect 297970 553560 300042 553616
rect 297909 553558 300042 553560
rect 297909 553555 297975 553558
rect 377814 553482 377874 553928
rect 379605 553482 379671 553485
rect 377814 553480 379671 553482
rect 377814 553424 379610 553480
rect 379666 553424 379671 553480
rect 377814 553422 379671 553424
rect 379605 553419 379671 553422
rect -960 553074 480 553164
rect 3141 553074 3207 553077
rect -960 553072 3207 553074
rect -960 553016 3146 553072
rect 3202 553016 3207 553072
rect -960 553014 3207 553016
rect -960 552924 480 553014
rect 3141 553011 3207 553014
rect 198406 552060 198412 552124
rect 198476 552122 198482 552124
rect 200070 552122 200130 552704
rect 198476 552062 200130 552122
rect 219942 552122 220002 552160
rect 222285 552122 222351 552125
rect 219942 552120 222351 552122
rect 219942 552064 222290 552120
rect 222346 552064 222351 552120
rect 219942 552062 222351 552064
rect 198476 552060 198482 552062
rect 222285 552059 222351 552062
rect 299289 550762 299355 550765
rect 299982 550762 300042 550936
rect 299289 550760 300042 550762
rect 299289 550704 299294 550760
rect 299350 550704 300042 550760
rect 299289 550702 300042 550704
rect 299289 550699 299355 550702
rect 378225 550694 378291 550697
rect 377844 550692 378291 550694
rect 377844 550636 378230 550692
rect 378286 550636 378291 550692
rect 377844 550634 378291 550636
rect 378225 550631 378291 550634
rect 86358 549949 86418 550528
rect 86358 549944 86467 549949
rect 86358 549888 86406 549944
rect 86462 549888 86467 549944
rect 86358 549886 86467 549888
rect 86401 549883 86467 549886
rect 198222 547844 198228 547908
rect 198292 547906 198298 547908
rect 200070 547906 200130 548080
rect 198292 547846 200130 547906
rect 299197 547906 299263 547909
rect 299982 547906 300042 547944
rect 299197 547904 300042 547906
rect 299197 547848 299202 547904
rect 299258 547848 300042 547904
rect 299197 547846 300042 547848
rect 198292 547844 198298 547846
rect 299197 547843 299263 547846
rect 378317 547702 378383 547705
rect 377844 547700 378383 547702
rect 377844 547644 378322 547700
rect 378378 547644 378383 547700
rect 377844 547642 378383 547644
rect 378317 547639 378383 547642
rect 219942 546954 220002 547536
rect 222561 546954 222627 546957
rect 219942 546952 222627 546954
rect 219942 546896 222566 546952
rect 222622 546896 222627 546952
rect 219942 546894 222627 546896
rect 222561 546891 222627 546894
rect 115614 546546 115674 546720
rect 118049 546546 118115 546549
rect 115614 546544 118115 546546
rect 115614 546488 118054 546544
rect 118110 546488 118115 546544
rect 115614 546486 118115 546488
rect 118049 546483 118115 546486
rect 84101 545866 84167 545869
rect 85990 545866 86050 546448
rect 84101 545864 86050 545866
rect 84101 545808 84106 545864
rect 84162 545808 86050 545864
rect 84101 545806 86050 545808
rect 84101 545803 84167 545806
rect 580349 545594 580415 545597
rect 583520 545594 584960 545684
rect 580349 545592 584960 545594
rect 580349 545536 580354 545592
rect 580410 545536 584960 545592
rect 580349 545534 584960 545536
rect 580349 545531 580415 545534
rect 583520 545444 584960 545534
rect 297817 544098 297883 544101
rect 299982 544098 300042 544680
rect 297817 544096 300042 544098
rect 297817 544040 297822 544096
rect 297878 544040 300042 544096
rect 297817 544038 300042 544040
rect 297817 544035 297883 544038
rect 198038 543764 198044 543828
rect 198108 543826 198114 543828
rect 377814 543826 377874 544408
rect 379697 543826 379763 543829
rect 198108 543766 200130 543826
rect 377814 543824 379763 543826
rect 377814 543768 379702 543824
rect 379758 543768 379763 543824
rect 377814 543766 379763 543768
rect 198108 543764 198114 543766
rect 200070 543728 200130 543766
rect 379697 543763 379763 543766
rect 219942 542602 220002 543184
rect 222469 542602 222535 542605
rect 219942 542600 222535 542602
rect 219942 542544 222474 542600
rect 222530 542544 222535 542600
rect 219942 542542 222535 542544
rect 222469 542539 222535 542542
rect 118233 542466 118299 542469
rect 115614 542464 118299 542466
rect 115614 542408 118238 542464
rect 118294 542408 118299 542464
rect 115614 542406 118299 542408
rect 115614 542368 115674 542406
rect 118233 542403 118299 542406
rect 84009 541514 84075 541517
rect 85990 541514 86050 542096
rect 84009 541512 86050 541514
rect 84009 541456 84014 541512
rect 84070 541456 86050 541512
rect 84009 541454 86050 541456
rect 84009 541451 84075 541454
rect 297357 541106 297423 541109
rect 299982 541106 300042 541688
rect 297357 541104 300042 541106
rect 297357 541048 297362 541104
rect 297418 541048 300042 541104
rect 297357 541046 300042 541048
rect 377814 541106 377874 541416
rect 379646 541106 379652 541108
rect 377814 541046 379652 541106
rect 297357 541043 297423 541046
rect 379646 541044 379652 541046
rect 379716 541044 379722 541108
rect -960 538658 480 538748
rect 3509 538658 3575 538661
rect -960 538656 3575 538658
rect -960 538600 3514 538656
rect 3570 538600 3575 538656
rect -960 538598 3575 538600
rect -960 538508 480 538598
rect 3509 538595 3575 538598
rect 197854 538460 197860 538524
rect 197924 538522 197930 538524
rect 200070 538522 200130 539104
rect 197924 538462 200130 538522
rect 197924 538460 197930 538462
rect 219942 538386 220002 538560
rect 222377 538386 222443 538389
rect 219942 538384 222443 538386
rect 219942 538328 222382 538384
rect 222438 538328 222443 538384
rect 219942 538326 222443 538328
rect 222377 538323 222443 538326
rect 297725 538386 297791 538389
rect 299982 538386 300042 538424
rect 297725 538384 300042 538386
rect 297725 538328 297730 538384
rect 297786 538328 300042 538384
rect 297725 538326 300042 538328
rect 297725 538323 297791 538326
rect 85573 537774 85639 537777
rect 85573 537772 86020 537774
rect 85573 537716 85578 537772
rect 85634 537716 86020 537772
rect 85573 537714 86020 537716
rect 85573 537711 85639 537714
rect 115614 537434 115674 538016
rect 377814 537570 377874 538152
rect 379789 537570 379855 537573
rect 377814 537568 379855 537570
rect 377814 537512 379794 537568
rect 379850 537512 379855 537568
rect 377814 537510 379855 537512
rect 379789 537507 379855 537510
rect 117313 537434 117379 537437
rect 115614 537432 117379 537434
rect 115614 537376 117318 537432
rect 117374 537376 117379 537432
rect 115614 537374 117379 537376
rect 117313 537371 117379 537374
rect 299565 535462 299631 535465
rect 299565 535460 300012 535462
rect 299565 535404 299570 535460
rect 299626 535404 300012 535460
rect 299565 535402 300012 535404
rect 299565 535399 299631 535402
rect 377814 534578 377874 535160
rect 379881 534578 379947 534581
rect 377814 534576 379947 534578
rect 377814 534520 379886 534576
rect 379942 534520 379947 534576
rect 377814 534518 379947 534520
rect 379881 534515 379947 534518
rect 198641 534170 198707 534173
rect 200070 534170 200130 534480
rect 198641 534168 200130 534170
rect 198641 534112 198646 534168
rect 198702 534112 200130 534168
rect 198641 534110 200130 534112
rect 198641 534107 198707 534110
rect 85297 533082 85363 533085
rect 85990 533082 86050 533664
rect 115614 533354 115674 533936
rect 117313 533354 117379 533357
rect 115614 533352 117379 533354
rect 115614 533296 117318 533352
rect 117374 533296 117379 533352
rect 115614 533294 117379 533296
rect 219942 533354 220002 533936
rect 580165 533898 580231 533901
rect 583520 533898 584960 533988
rect 580165 533896 584960 533898
rect 580165 533840 580170 533896
rect 580226 533840 584960 533896
rect 580165 533838 584960 533840
rect 580165 533835 580231 533838
rect 583520 533748 584960 533838
rect 222653 533354 222719 533357
rect 219942 533352 222719 533354
rect 219942 533296 222658 533352
rect 222714 533296 222719 533352
rect 219942 533294 222719 533296
rect 117313 533291 117379 533294
rect 222653 533291 222719 533294
rect 85297 533080 86050 533082
rect 85297 533024 85302 533080
rect 85358 533024 86050 533080
rect 85297 533022 86050 533024
rect 85297 533019 85363 533022
rect 296529 531450 296595 531453
rect 299982 531450 300042 532168
rect 296529 531448 300042 531450
rect 296529 531392 296534 531448
rect 296590 531392 300042 531448
rect 296529 531390 300042 531392
rect 377814 531450 377874 531896
rect 379973 531450 380039 531453
rect 377814 531448 380039 531450
rect 377814 531392 379978 531448
rect 380034 531392 380039 531448
rect 377814 531390 380039 531392
rect 296529 531387 296595 531390
rect 379973 531387 380039 531390
rect 153469 531314 153535 531317
rect 153745 531314 153811 531317
rect 153469 531312 153811 531314
rect 153469 531256 153474 531312
rect 153530 531256 153750 531312
rect 153806 531256 153811 531312
rect 153469 531254 153811 531256
rect 153469 531251 153535 531254
rect 153745 531251 153811 531254
rect 115614 529546 115674 529584
rect 117957 529546 118023 529549
rect 115614 529544 118023 529546
rect 115614 529488 117962 529544
rect 118018 529488 118023 529544
rect 115614 529486 118023 529488
rect 117957 529483 118023 529486
rect 83917 528730 83983 528733
rect 85990 528730 86050 529312
rect 198733 529274 198799 529277
rect 200070 529274 200130 529856
rect 198733 529272 200130 529274
rect 198733 529216 198738 529272
rect 198794 529216 200130 529272
rect 198733 529214 200130 529216
rect 198733 529211 198799 529214
rect 219942 529002 220002 529312
rect 222745 529002 222811 529005
rect 219942 529000 222811 529002
rect 219942 528944 222750 529000
rect 222806 528944 222811 529000
rect 219942 528942 222811 528944
rect 222745 528939 222811 528942
rect 297449 528866 297515 528869
rect 299982 528866 300042 529176
rect 297449 528864 300042 528866
rect 297449 528808 297454 528864
rect 297510 528808 300042 528864
rect 297449 528806 300042 528808
rect 297449 528803 297515 528806
rect 83917 528728 86050 528730
rect 83917 528672 83922 528728
rect 83978 528672 86050 528728
rect 83917 528670 86050 528672
rect 377814 528730 377874 528904
rect 380525 528730 380591 528733
rect 377814 528728 380591 528730
rect 377814 528672 380530 528728
rect 380586 528672 380591 528728
rect 377814 528670 380591 528672
rect 83917 528667 83983 528670
rect 380525 528667 380591 528670
rect 299105 525874 299171 525877
rect 299982 525874 300042 525912
rect 299105 525872 300042 525874
rect 299105 525816 299110 525872
rect 299166 525816 300042 525872
rect 299105 525814 300042 525816
rect 299105 525811 299171 525814
rect 85389 525602 85455 525605
rect 85389 525600 86050 525602
rect 85389 525544 85394 525600
rect 85450 525544 86050 525600
rect 85389 525542 86050 525544
rect 85389 525539 85455 525542
rect 82813 524922 82879 524925
rect 85990 524922 86050 525542
rect 115614 525194 115674 525232
rect 117313 525194 117379 525197
rect 115614 525192 117379 525194
rect 115614 525136 117318 525192
rect 117374 525136 117379 525192
rect 115614 525134 117379 525136
rect 117313 525131 117379 525134
rect 82813 524920 86050 524922
rect 82813 524864 82818 524920
rect 82874 524864 86050 524920
rect 82813 524862 86050 524864
rect 82813 524859 82879 524862
rect 198549 524650 198615 524653
rect 200070 524650 200130 525232
rect 377814 525058 377874 525640
rect 380065 525058 380131 525061
rect 377814 525056 380131 525058
rect 377814 525000 380070 525056
rect 380126 525000 380131 525056
rect 377814 524998 380131 525000
rect 380065 524995 380131 524998
rect 198549 524648 200130 524650
rect 198549 524592 198554 524648
rect 198610 524592 200130 524648
rect 198549 524590 200130 524592
rect 198549 524587 198615 524590
rect 219942 524514 220002 524688
rect 222837 524514 222903 524517
rect 219942 524512 222903 524514
rect 219942 524456 222842 524512
rect 222898 524456 222903 524512
rect 219942 524454 222903 524456
rect 222837 524451 222903 524454
rect -960 524092 480 524332
rect 297081 522202 297147 522205
rect 299982 522202 300042 522648
rect 297081 522200 300042 522202
rect 297081 522144 297086 522200
rect 297142 522144 300042 522200
rect 297081 522142 300042 522144
rect 297081 522139 297147 522142
rect 377814 521794 377874 522376
rect 583520 521916 584960 522156
rect 380157 521794 380223 521797
rect 377814 521792 380223 521794
rect 377814 521736 380162 521792
rect 380218 521736 380223 521792
rect 377814 521734 380223 521736
rect 380157 521731 380223 521734
rect 118233 521658 118299 521661
rect 118417 521658 118483 521661
rect 118233 521656 118483 521658
rect 118233 521600 118238 521656
rect 118294 521600 118422 521656
rect 118478 521600 118483 521656
rect 118233 521598 118483 521600
rect 118233 521595 118299 521598
rect 118417 521595 118483 521598
rect 115614 521114 115674 521152
rect 117313 521114 117379 521117
rect 115614 521112 117379 521114
rect 115614 521056 117318 521112
rect 117374 521056 117379 521112
rect 115614 521054 117379 521056
rect 117313 521051 117379 521054
rect 297725 519210 297791 519213
rect 299982 519210 300042 519656
rect 297725 519208 300042 519210
rect 297725 519152 297730 519208
rect 297786 519152 300042 519208
rect 297725 519150 300042 519152
rect 377814 519210 377874 519384
rect 380709 519210 380775 519213
rect 377814 519208 380775 519210
rect 377814 519152 380714 519208
rect 380770 519152 380775 519208
rect 377814 519150 380775 519152
rect 297725 519147 297791 519150
rect 380709 519147 380775 519150
rect 297725 516218 297791 516221
rect 299982 516218 300042 516392
rect 297725 516216 300042 516218
rect 297725 516160 297730 516216
rect 297786 516160 300042 516216
rect 297725 516158 300042 516160
rect 297725 516155 297791 516158
rect 377814 515538 377874 516120
rect 378961 515538 379027 515541
rect 377814 515536 379027 515538
rect 377814 515480 378966 515536
rect 379022 515480 379027 515536
rect 377814 515478 379027 515480
rect 378961 515475 379027 515478
rect 297725 513498 297791 513501
rect 297725 513496 300042 513498
rect 297725 513440 297730 513496
rect 297786 513440 300042 513496
rect 297725 513438 300042 513440
rect 297725 513435 297791 513438
rect 299982 513400 300042 513438
rect 377814 512546 377874 513128
rect 380249 512546 380315 512549
rect 377814 512544 380315 512546
rect 377814 512488 380254 512544
rect 380310 512488 380315 512544
rect 377814 512486 380315 512488
rect 380249 512483 380315 512486
rect 128537 512002 128603 512005
rect 128721 512002 128787 512005
rect 128537 512000 128787 512002
rect 128537 511944 128542 512000
rect 128598 511944 128726 512000
rect 128782 511944 128787 512000
rect 128537 511942 128787 511944
rect 128537 511939 128603 511942
rect 128721 511939 128787 511942
rect 580441 510370 580507 510373
rect 583520 510370 584960 510460
rect 580441 510368 584960 510370
rect 580441 510312 580446 510368
rect 580502 510312 584960 510368
rect 580441 510310 584960 510312
rect 580441 510307 580507 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3601 509962 3667 509965
rect -960 509960 3667 509962
rect -960 509904 3606 509960
rect 3662 509904 3667 509960
rect -960 509902 3667 509904
rect -960 509812 480 509902
rect 3601 509899 3667 509902
rect 297633 509690 297699 509693
rect 299982 509690 300042 510136
rect 297633 509688 300042 509690
rect 297633 509632 297638 509688
rect 297694 509632 300042 509688
rect 297633 509630 300042 509632
rect 297633 509627 297699 509630
rect 377814 509418 377874 509864
rect 380341 509418 380407 509421
rect 377814 509416 380407 509418
rect 377814 509360 380346 509416
rect 380402 509360 380407 509416
rect 377814 509358 380407 509360
rect 380341 509355 380407 509358
rect 297633 506698 297699 506701
rect 299982 506698 300042 507144
rect 297633 506696 300042 506698
rect 297633 506640 297638 506696
rect 297694 506640 300042 506696
rect 297633 506638 300042 506640
rect 297633 506635 297699 506638
rect 377814 506562 377874 506872
rect 380433 506562 380499 506565
rect 377814 506560 380499 506562
rect 377814 506504 380438 506560
rect 380494 506504 380499 506560
rect 377814 506502 380499 506504
rect 380433 506499 380499 506502
rect 299657 503910 299723 503913
rect 299657 503908 300012 503910
rect 299657 503852 299662 503908
rect 299718 503852 300012 503908
rect 299657 503850 300012 503852
rect 299657 503847 299723 503850
rect 377814 503026 377874 503608
rect 380709 503026 380775 503029
rect 377814 503024 380775 503026
rect 377814 502968 380714 503024
rect 380770 502968 380775 503024
rect 377814 502966 380775 502968
rect 380709 502963 380775 502966
rect 131021 500306 131087 500309
rect 379462 500306 379468 500308
rect 131021 500304 379468 500306
rect 131021 500248 131026 500304
rect 131082 500248 379468 500304
rect 131021 500246 379468 500248
rect 131021 500243 131087 500246
rect 379462 500244 379468 500246
rect 379532 500244 379538 500308
rect 130929 500170 130995 500173
rect 379646 500170 379652 500172
rect 130929 500168 379652 500170
rect 130929 500112 130934 500168
rect 130990 500112 379652 500168
rect 130929 500110 379652 500112
rect 130929 500107 130995 500110
rect 379646 500108 379652 500110
rect 379716 500108 379722 500172
rect 580165 498674 580231 498677
rect 583520 498674 584960 498764
rect 580165 498672 584960 498674
rect 580165 498616 580170 498672
rect 580226 498616 584960 498672
rect 580165 498614 584960 498616
rect 580165 498611 580231 498614
rect 583520 498524 584960 498614
rect 118417 498130 118483 498133
rect 319713 498130 319779 498133
rect 118417 498128 319779 498130
rect 118417 498072 118422 498128
rect 118478 498072 319718 498128
rect 319774 498072 319779 498128
rect 118417 498070 319779 498072
rect 118417 498067 118483 498070
rect 319713 498067 319779 498070
rect -960 495546 480 495636
rect 3325 495546 3391 495549
rect -960 495544 3391 495546
rect -960 495488 3330 495544
rect 3386 495488 3391 495544
rect -960 495486 3391 495488
rect -960 495396 480 495486
rect 3325 495483 3391 495486
rect 304165 492690 304231 492693
rect 304533 492690 304599 492693
rect 304165 492688 304599 492690
rect 304165 492632 304170 492688
rect 304226 492632 304538 492688
rect 304594 492632 304599 492688
rect 304165 492630 304599 492632
rect 304165 492627 304231 492630
rect 304533 492627 304599 492630
rect 580165 486842 580231 486845
rect 583520 486842 584960 486932
rect 580165 486840 584960 486842
rect 580165 486784 580170 486840
rect 580226 486784 584960 486840
rect 580165 486782 584960 486784
rect 580165 486779 580231 486782
rect 583520 486692 584960 486782
rect 118325 483034 118391 483037
rect 118601 483034 118667 483037
rect 118325 483032 118667 483034
rect 118325 482976 118330 483032
rect 118386 482976 118606 483032
rect 118662 482976 118667 483032
rect 118325 482974 118667 482976
rect 118325 482971 118391 482974
rect 118601 482971 118667 482974
rect 128537 483034 128603 483037
rect 128813 483034 128879 483037
rect 128537 483032 128879 483034
rect 128537 482976 128542 483032
rect 128598 482976 128818 483032
rect 128874 482976 128879 483032
rect 128537 482974 128879 482976
rect 128537 482971 128603 482974
rect 128813 482971 128879 482974
rect 153285 483034 153351 483037
rect 153469 483034 153535 483037
rect 153285 483032 153535 483034
rect 153285 482976 153290 483032
rect 153346 482976 153474 483032
rect 153530 482976 153535 483032
rect 153285 482974 153535 482976
rect 153285 482971 153351 482974
rect 153469 482971 153535 482974
rect -960 481130 480 481220
rect 4061 481130 4127 481133
rect -960 481128 4127 481130
rect -960 481072 4066 481128
rect 4122 481072 4127 481128
rect -960 481070 4127 481072
rect -960 480980 480 481070
rect 4061 481067 4127 481070
rect 583520 474996 584960 475236
rect 304257 473378 304323 473381
rect 304441 473378 304507 473381
rect 304257 473376 304507 473378
rect 304257 473320 304262 473376
rect 304318 473320 304446 473376
rect 304502 473320 304507 473376
rect 304257 473318 304507 473320
rect 304257 473315 304323 473318
rect 304441 473315 304507 473318
rect -960 466700 480 466940
rect 128537 463722 128603 463725
rect 128813 463722 128879 463725
rect 128537 463720 128879 463722
rect 128537 463664 128542 463720
rect 128598 463664 128818 463720
rect 128874 463664 128879 463720
rect 128537 463662 128879 463664
rect 128537 463659 128603 463662
rect 128813 463659 128879 463662
rect 579797 463450 579863 463453
rect 583520 463450 584960 463540
rect 579797 463448 584960 463450
rect 579797 463392 579802 463448
rect 579858 463392 584960 463448
rect 579797 463390 584960 463392
rect 579797 463387 579863 463390
rect 583520 463300 584960 463390
rect 118049 454066 118115 454069
rect 118233 454066 118299 454069
rect 118049 454064 118299 454066
rect 118049 454008 118054 454064
rect 118110 454008 118238 454064
rect 118294 454008 118299 454064
rect 118049 454006 118299 454008
rect 118049 454003 118115 454006
rect 118233 454003 118299 454006
rect -960 452434 480 452524
rect 3049 452434 3115 452437
rect -960 452432 3115 452434
rect -960 452376 3054 452432
rect 3110 452376 3115 452432
rect -960 452374 3115 452376
rect -960 452284 480 452374
rect 3049 452371 3115 452374
rect 580165 451754 580231 451757
rect 583520 451754 584960 451844
rect 580165 451752 584960 451754
rect 580165 451696 580170 451752
rect 580226 451696 584960 451752
rect 580165 451694 584960 451696
rect 580165 451691 580231 451694
rect 583520 451604 584960 451694
rect 128537 444410 128603 444413
rect 128813 444410 128879 444413
rect 128537 444408 128879 444410
rect 128537 444352 128542 444408
rect 128598 444352 128818 444408
rect 128874 444352 128879 444408
rect 128537 444350 128879 444352
rect 128537 444347 128603 444350
rect 128813 444347 128879 444350
rect 580165 439922 580231 439925
rect 583520 439922 584960 440012
rect 580165 439920 584960 439922
rect 580165 439864 580170 439920
rect 580226 439864 584960 439920
rect 580165 439862 584960 439864
rect 580165 439859 580231 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3693 438018 3759 438021
rect -960 438016 3759 438018
rect -960 437960 3698 438016
rect 3754 437960 3759 438016
rect -960 437958 3759 437960
rect -960 437868 480 437958
rect 3693 437955 3759 437958
rect 118049 434754 118115 434757
rect 118233 434754 118299 434757
rect 118049 434752 118299 434754
rect 118049 434696 118054 434752
rect 118110 434696 118238 434752
rect 118294 434696 118299 434752
rect 118049 434694 118299 434696
rect 118049 434691 118115 434694
rect 118233 434691 118299 434694
rect 583520 428076 584960 428316
rect 153469 425234 153535 425237
rect 153150 425232 153535 425234
rect 153150 425176 153474 425232
rect 153530 425176 153535 425232
rect 153150 425174 153535 425176
rect 153150 425101 153210 425174
rect 153469 425171 153535 425174
rect 128537 425098 128603 425101
rect 128813 425098 128879 425101
rect 128537 425096 128879 425098
rect 128537 425040 128542 425096
rect 128598 425040 128818 425096
rect 128874 425040 128879 425096
rect 128537 425038 128879 425040
rect 153150 425096 153259 425101
rect 153150 425040 153198 425096
rect 153254 425040 153259 425096
rect 153150 425038 153259 425040
rect 128537 425035 128603 425038
rect 128813 425035 128879 425038
rect 153193 425035 153259 425038
rect -960 423738 480 423828
rect 4061 423738 4127 423741
rect -960 423736 4127 423738
rect -960 423680 4066 423736
rect 4122 423680 4127 423736
rect -960 423678 4127 423680
rect -960 423588 480 423678
rect 4061 423675 4127 423678
rect 579797 416530 579863 416533
rect 583520 416530 584960 416620
rect 579797 416528 584960 416530
rect 579797 416472 579802 416528
rect 579858 416472 584960 416528
rect 579797 416470 584960 416472
rect 579797 416467 579863 416470
rect 583520 416380 584960 416470
rect 203333 410410 203399 410413
rect 266854 410410 266860 410412
rect 203333 410408 266860 410410
rect 203333 410352 203338 410408
rect 203394 410352 266860 410408
rect 203333 410350 266860 410352
rect 203333 410347 203399 410350
rect 266854 410348 266860 410350
rect 266924 410348 266930 410412
rect 231853 410274 231919 410277
rect 267958 410274 267964 410276
rect 231853 410272 267964 410274
rect 231853 410216 231858 410272
rect 231914 410216 267964 410272
rect 231853 410214 267964 410216
rect 231853 410211 231919 410214
rect 267958 410212 267964 410214
rect 268028 410212 268034 410276
rect 226149 410138 226215 410141
rect 267774 410138 267780 410140
rect 226149 410136 267780 410138
rect 226149 410080 226154 410136
rect 226210 410080 267780 410136
rect 226149 410078 267780 410080
rect 226149 410075 226215 410078
rect 267774 410076 267780 410078
rect 267844 410076 267850 410140
rect 263133 410002 263199 410005
rect 268142 410002 268148 410004
rect 263133 410000 268148 410002
rect 263133 409944 263138 410000
rect 263194 409944 268148 410000
rect 263133 409942 268148 409944
rect 263133 409939 263199 409942
rect 268142 409940 268148 409942
rect 268212 409940 268218 410004
rect -960 409172 480 409412
rect 580625 404834 580691 404837
rect 583520 404834 584960 404924
rect 580625 404832 584960 404834
rect 580625 404776 580630 404832
rect 580686 404776 584960 404832
rect 580625 404774 584960 404776
rect 580625 404771 580691 404774
rect 583520 404684 584960 404774
rect 198825 403746 198891 403749
rect 267825 403746 267891 403749
rect 198825 403744 200100 403746
rect 198825 403688 198830 403744
rect 198886 403688 200100 403744
rect 198825 403686 200100 403688
rect 266524 403744 267891 403746
rect 266524 403688 267830 403744
rect 267886 403688 267891 403744
rect 266524 403686 267891 403688
rect 198825 403683 198891 403686
rect 267825 403683 267891 403686
rect 198457 399666 198523 399669
rect 267181 399666 267247 399669
rect 198457 399664 200100 399666
rect 198457 399608 198462 399664
rect 198518 399608 200100 399664
rect 198457 399606 200100 399608
rect 266524 399664 267247 399666
rect 266524 399608 267186 399664
rect 267242 399608 267247 399664
rect 266524 399606 267247 399608
rect 198457 399603 198523 399606
rect 267181 399603 267247 399606
rect 198917 395314 198983 395317
rect 267917 395314 267983 395317
rect 198917 395312 200100 395314
rect 198917 395256 198922 395312
rect 198978 395256 200100 395312
rect 198917 395254 200100 395256
rect 266524 395312 267983 395314
rect 266524 395256 267922 395312
rect 267978 395256 267983 395312
rect 266524 395254 267983 395256
rect 198917 395251 198983 395254
rect 267917 395251 267983 395254
rect -960 395042 480 395132
rect 3877 395042 3943 395045
rect -960 395040 3943 395042
rect -960 394984 3882 395040
rect 3938 394984 3943 395040
rect -960 394982 3943 394984
rect -960 394892 480 394982
rect 3877 394979 3943 394982
rect 580533 393002 580599 393005
rect 583520 393002 584960 393092
rect 580533 393000 584960 393002
rect 580533 392944 580538 393000
rect 580594 392944 584960 393000
rect 580533 392942 584960 392944
rect 580533 392939 580599 392942
rect 583520 392852 584960 392942
rect 71589 392594 71655 392597
rect 71589 392592 72036 392594
rect 71589 392536 71594 392592
rect 71650 392536 72036 392592
rect 71589 392534 72036 392536
rect 71589 392531 71655 392534
rect 288341 392186 288407 392189
rect 288022 392184 288407 392186
rect 288022 392128 288346 392184
rect 288402 392128 288407 392184
rect 288022 392126 288407 392128
rect 288022 392050 288082 392126
rect 288341 392123 288407 392126
rect 288157 392050 288223 392053
rect 288022 392048 288223 392050
rect 288022 391992 288162 392048
rect 288218 391992 288223 392048
rect 288022 391990 288223 391992
rect 288157 391987 288223 391990
rect 199009 391234 199075 391237
rect 268009 391234 268075 391237
rect 199009 391232 200100 391234
rect 199009 391176 199014 391232
rect 199070 391176 200100 391232
rect 199009 391174 200100 391176
rect 266524 391232 268075 391234
rect 266524 391176 268014 391232
rect 268070 391176 268075 391232
rect 266524 391174 268075 391176
rect 199009 391171 199075 391174
rect 268009 391171 268075 391174
rect 128721 388514 128787 388517
rect 126102 388512 128787 388514
rect 126102 388456 128726 388512
rect 128782 388456 128787 388512
rect 126102 388454 128787 388456
rect 126102 387940 126162 388454
rect 128721 388451 128787 388454
rect 198365 387154 198431 387157
rect 198365 387152 200100 387154
rect 198365 387096 198370 387152
rect 198426 387096 200100 387152
rect 198365 387094 200100 387096
rect 198365 387091 198431 387094
rect 268101 386882 268167 386885
rect 266524 386880 268167 386882
rect 266524 386824 268106 386880
rect 268162 386824 268167 386880
rect 266524 386822 268167 386824
rect 268101 386819 268167 386822
rect 69933 385250 69999 385253
rect 69933 385248 72036 385250
rect 69933 385192 69938 385248
rect 69994 385192 72036 385248
rect 69933 385190 72036 385192
rect 69933 385187 69999 385190
rect 199101 382802 199167 382805
rect 268193 382802 268259 382805
rect 199101 382800 200100 382802
rect 199101 382744 199106 382800
rect 199162 382744 200100 382800
rect 199101 382742 200100 382744
rect 266524 382800 268259 382802
rect 266524 382744 268198 382800
rect 268254 382744 268259 382800
rect 266524 382742 268259 382744
rect 199101 382739 199167 382742
rect 268193 382739 268259 382742
rect 288341 382258 288407 382261
rect 288525 382258 288591 382261
rect 288341 382256 288591 382258
rect 288341 382200 288346 382256
rect 288402 382200 288530 382256
rect 288586 382200 288591 382256
rect 288341 382198 288591 382200
rect 288341 382195 288407 382198
rect 288525 382195 288591 382198
rect 380893 381442 380959 381445
rect 380893 381440 384130 381442
rect 380893 381384 380898 381440
rect 380954 381384 384130 381440
rect 380893 381382 384130 381384
rect 380893 381379 380959 381382
rect 384070 381344 384130 381382
rect 583520 381156 584960 381396
rect 416865 380898 416931 380901
rect 415166 380896 416931 380898
rect 415166 380840 416870 380896
rect 416926 380840 416931 380896
rect 415166 380838 416931 380840
rect 415166 380800 415226 380838
rect 416865 380835 416931 380838
rect -960 380626 480 380716
rect 3785 380626 3851 380629
rect 129089 380626 129155 380629
rect -960 380624 3851 380626
rect -960 380568 3790 380624
rect 3846 380568 3851 380624
rect -960 380566 3851 380568
rect 126132 380624 129155 380626
rect 126132 380568 129094 380624
rect 129150 380568 129155 380624
rect 126132 380566 129155 380568
rect -960 380476 480 380566
rect 3785 380563 3851 380566
rect 129089 380563 129155 380566
rect 197997 378722 198063 378725
rect 197997 378720 200100 378722
rect 197997 378664 198002 378720
rect 198058 378664 200100 378720
rect 197997 378662 200100 378664
rect 197997 378659 198063 378662
rect 268285 378450 268351 378453
rect 266524 378448 268351 378450
rect 266524 378392 268290 378448
rect 268346 378392 268351 378448
rect 266524 378390 268351 378392
rect 268285 378387 268351 378390
rect 504725 378450 504791 378453
rect 504725 378448 504834 378450
rect 504725 378392 504730 378448
rect 504786 378392 504834 378448
rect 504725 378387 504834 378392
rect 504774 378148 504834 378387
rect 70209 377906 70275 377909
rect 71037 377906 71103 377909
rect 70209 377904 72036 377906
rect 70209 377848 70214 377904
rect 70270 377848 71042 377904
rect 71098 377848 72036 377904
rect 70209 377846 72036 377848
rect 70209 377843 70275 377846
rect 71037 377843 71103 377846
rect 380893 377226 380959 377229
rect 384070 377226 384130 377808
rect 380893 377224 384130 377226
rect 380893 377168 380898 377224
rect 380954 377168 384130 377224
rect 380893 377166 384130 377168
rect 380893 377163 380959 377166
rect 415166 376954 415226 377536
rect 416773 376954 416839 376957
rect 415166 376952 416839 376954
rect 415166 376896 416778 376952
rect 416834 376896 416839 376952
rect 415166 376894 416839 376896
rect 416773 376891 416839 376894
rect 456793 375186 456859 375189
rect 456793 375184 460092 375186
rect 456793 375128 456798 375184
rect 456854 375128 460092 375184
rect 456793 375126 460092 375128
rect 456793 375123 456859 375126
rect 416957 374642 417023 374645
rect 415166 374640 417023 374642
rect 415166 374584 416962 374640
rect 417018 374584 417023 374640
rect 415166 374582 417023 374584
rect 197905 374370 197971 374373
rect 268377 374370 268443 374373
rect 197905 374368 200100 374370
rect 197905 374312 197910 374368
rect 197966 374312 200100 374368
rect 197905 374310 200100 374312
rect 266524 374368 268443 374370
rect 266524 374312 268382 374368
rect 268438 374312 268443 374368
rect 266524 374310 268443 374312
rect 197905 374307 197971 374310
rect 268377 374307 268443 374310
rect 380893 374098 380959 374101
rect 384070 374098 384130 374544
rect 380893 374096 384130 374098
rect 380893 374040 380898 374096
rect 380954 374040 384130 374096
rect 380893 374038 384130 374040
rect 380893 374035 380959 374038
rect 415166 374000 415226 374582
rect 416957 374579 417023 374582
rect 128445 373282 128511 373285
rect 129181 373282 129247 373285
rect 126132 373280 129247 373282
rect 126132 373224 128450 373280
rect 128506 373224 129186 373280
rect 129242 373224 129247 373280
rect 126132 373222 129247 373224
rect 128445 373219 128511 373222
rect 129181 373219 129247 373222
rect 380893 370426 380959 370429
rect 384070 370426 384130 371008
rect 380893 370424 384130 370426
rect 380893 370368 380898 370424
rect 380954 370368 384130 370424
rect 380893 370366 384130 370368
rect 380893 370363 380959 370366
rect 70117 370290 70183 370293
rect 71589 370290 71655 370293
rect 197813 370290 197879 370293
rect 70117 370288 72036 370290
rect 70117 370232 70122 370288
rect 70178 370232 71594 370288
rect 71650 370232 72036 370288
rect 70117 370230 72036 370232
rect 197813 370288 200100 370290
rect 197813 370232 197818 370288
rect 197874 370232 200100 370288
rect 197813 370230 200100 370232
rect 70117 370227 70183 370230
rect 71589 370227 71655 370230
rect 197813 370227 197879 370230
rect 415166 370154 415226 370736
rect 416865 370154 416931 370157
rect 415166 370152 416931 370154
rect 415166 370096 416870 370152
rect 416926 370096 416931 370152
rect 415166 370094 416931 370096
rect 416865 370091 416931 370094
rect 268469 370018 268535 370021
rect 266524 370016 268535 370018
rect 266524 369960 268474 370016
rect 268530 369960 268535 370016
rect 266524 369958 268535 369960
rect 268469 369955 268535 369958
rect 580717 369610 580783 369613
rect 583520 369610 584960 369700
rect 580717 369608 584960 369610
rect 580717 369552 580722 369608
rect 580778 369552 584960 369608
rect 580717 369550 584960 369552
rect 580717 369547 580783 369550
rect 583520 369460 584960 369550
rect 381629 367434 381695 367437
rect 384070 367434 384130 367744
rect 381629 367432 384130 367434
rect 381629 367376 381634 367432
rect 381690 367376 384130 367432
rect 381629 367374 384130 367376
rect 381629 367371 381695 367374
rect 415166 367162 415226 367200
rect 416957 367162 417023 367165
rect 415166 367160 417023 367162
rect 415166 367104 416962 367160
rect 417018 367104 417023 367160
rect 415166 367102 417023 367104
rect 416957 367099 417023 367102
rect -960 366210 480 366300
rect 2773 366210 2839 366213
rect -960 366208 2839 366210
rect -960 366152 2778 366208
rect 2834 366152 2839 366208
rect -960 366150 2839 366152
rect -960 366060 480 366150
rect 2773 366147 2839 366150
rect 129365 365938 129431 365941
rect 126132 365936 129431 365938
rect 126132 365880 129370 365936
rect 129426 365880 129431 365936
rect 126132 365878 129431 365880
rect 129365 365875 129431 365878
rect 199193 365938 199259 365941
rect 268561 365938 268627 365941
rect 199193 365936 200100 365938
rect 199193 365880 199198 365936
rect 199254 365880 200100 365936
rect 199193 365878 200100 365880
rect 266524 365936 268627 365938
rect 266524 365880 268566 365936
rect 268622 365880 268627 365936
rect 266524 365878 268627 365880
rect 199193 365875 199259 365878
rect 268561 365875 268627 365878
rect 380893 363626 380959 363629
rect 384070 363626 384130 364208
rect 415393 363966 415459 363969
rect 415196 363964 415459 363966
rect 415196 363908 415398 363964
rect 415454 363908 415459 363964
rect 415196 363906 415459 363908
rect 415393 363903 415459 363906
rect 380893 363624 384130 363626
rect 380893 363568 380898 363624
rect 380954 363568 384130 363624
rect 380893 363566 384130 363568
rect 380893 363563 380959 363566
rect 70025 362946 70091 362949
rect 70025 362944 72036 362946
rect 70025 362888 70030 362944
rect 70086 362888 72036 362944
rect 70025 362886 72036 362888
rect 70025 362883 70091 362886
rect 197721 361858 197787 361861
rect 197721 361856 200100 361858
rect 197721 361800 197726 361856
rect 197782 361800 200100 361856
rect 197721 361798 200100 361800
rect 197721 361795 197787 361798
rect 268653 361586 268719 361589
rect 266524 361584 268719 361586
rect 266524 361528 268658 361584
rect 268714 361528 268719 361584
rect 266524 361526 268719 361528
rect 268653 361523 268719 361526
rect 381721 360362 381787 360365
rect 384070 360362 384130 360944
rect 504774 360501 504834 361012
rect 504725 360496 504834 360501
rect 504725 360440 504730 360496
rect 504786 360440 504834 360496
rect 504725 360438 504834 360440
rect 504725 360435 504791 360438
rect 381721 360360 384130 360362
rect 381721 360304 381726 360360
rect 381782 360304 384130 360360
rect 381721 360302 384130 360304
rect 381721 360299 381787 360302
rect 415166 360226 415226 360400
rect 417049 360226 417115 360229
rect 415166 360224 417115 360226
rect 415166 360168 417054 360224
rect 417110 360168 417115 360224
rect 415166 360166 417115 360168
rect 417049 360163 417115 360166
rect 128353 358322 128419 358325
rect 129273 358322 129339 358325
rect 126132 358320 129339 358322
rect 126132 358264 128358 358320
rect 128414 358264 129278 358320
rect 129334 358264 129339 358320
rect 126132 358262 129339 358264
rect 128353 358259 128419 358262
rect 129273 358259 129339 358262
rect 457437 358050 457503 358053
rect 457437 358048 460092 358050
rect 457437 357992 457442 358048
rect 457498 357992 460092 358048
rect 457437 357990 460092 357992
rect 457437 357987 457503 357990
rect 580809 357914 580875 357917
rect 583520 357914 584960 358004
rect 580809 357912 584960 357914
rect 580809 357856 580814 357912
rect 580870 357856 584960 357912
rect 580809 357854 584960 357856
rect 580809 357851 580875 357854
rect 583520 357764 584960 357854
rect 197537 357506 197603 357509
rect 267273 357506 267339 357509
rect 197537 357504 200100 357506
rect 197537 357448 197542 357504
rect 197598 357448 200100 357504
rect 197537 357446 200100 357448
rect 266524 357504 267339 357506
rect 266524 357448 267278 357504
rect 267334 357448 267339 357504
rect 266524 357446 267339 357448
rect 197537 357443 197603 357446
rect 267273 357443 267339 357446
rect 381813 356826 381879 356829
rect 384070 356826 384130 357408
rect 381813 356824 384130 356826
rect 381813 356768 381818 356824
rect 381874 356768 384130 356824
rect 381813 356766 384130 356768
rect 381813 356763 381879 356766
rect 415166 356554 415226 357136
rect 417141 356554 417207 356557
rect 415166 356552 417207 356554
rect 415166 356496 417146 356552
rect 417202 356496 417207 356552
rect 415166 356494 417207 356496
rect 417141 356491 417207 356494
rect 70209 355602 70275 355605
rect 70209 355600 72036 355602
rect 70209 355544 70214 355600
rect 70270 355544 72036 355600
rect 70209 355542 72036 355544
rect 70209 355539 70275 355542
rect 380893 353562 380959 353565
rect 384070 353562 384130 354144
rect 380893 353560 384130 353562
rect 380893 353504 380898 353560
rect 380954 353504 384130 353560
rect 380893 353502 384130 353504
rect 380893 353499 380959 353502
rect 197445 353426 197511 353429
rect 267365 353426 267431 353429
rect 197445 353424 200100 353426
rect 197445 353368 197450 353424
rect 197506 353368 200100 353424
rect 197445 353366 200100 353368
rect 266524 353424 267431 353426
rect 266524 353368 267370 353424
rect 267426 353368 267431 353424
rect 266524 353366 267431 353368
rect 415166 353426 415226 353600
rect 417233 353426 417299 353429
rect 415166 353424 417299 353426
rect 415166 353368 417238 353424
rect 417294 353368 417299 353424
rect 415166 353366 417299 353368
rect 197445 353363 197511 353366
rect 267365 353363 267431 353366
rect 417233 353363 417299 353366
rect -960 351780 480 352020
rect 128997 350978 129063 350981
rect 126132 350976 129063 350978
rect 126132 350920 129002 350976
rect 129058 350920 129063 350976
rect 126132 350918 129063 350920
rect 128997 350915 129063 350918
rect 197353 349074 197419 349077
rect 267457 349074 267523 349077
rect 197353 349072 200100 349074
rect 197353 349016 197358 349072
rect 197414 349016 200100 349072
rect 197353 349014 200100 349016
rect 266524 349072 267523 349074
rect 266524 349016 267462 349072
rect 267518 349016 267523 349072
rect 266524 349014 267523 349016
rect 197353 349011 197419 349014
rect 267457 349011 267523 349014
rect 70301 348258 70367 348261
rect 71497 348258 71563 348261
rect 70301 348256 72036 348258
rect 70301 348200 70306 348256
rect 70362 348200 71502 348256
rect 71558 348200 72036 348256
rect 70301 348198 72036 348200
rect 70301 348195 70367 348198
rect 71497 348195 71563 348198
rect 579981 346082 580047 346085
rect 583520 346082 584960 346172
rect 579981 346080 584960 346082
rect 579981 346024 579986 346080
rect 580042 346024 584960 346080
rect 579981 346022 584960 346024
rect 579981 346019 580047 346022
rect 583520 345932 584960 346022
rect 197629 344994 197695 344997
rect 269021 344994 269087 344997
rect 197629 344992 200100 344994
rect 197629 344936 197634 344992
rect 197690 344936 200100 344992
rect 197629 344934 200100 344936
rect 266524 344992 269087 344994
rect 266524 344936 269026 344992
rect 269082 344936 269087 344992
rect 266524 344934 269087 344936
rect 197629 344931 197695 344934
rect 269021 344931 269087 344934
rect 504774 343637 504834 343876
rect 128997 343634 129063 343637
rect 126132 343632 129063 343634
rect 126132 343576 129002 343632
rect 129058 343576 129063 343632
rect 126132 343574 129063 343576
rect 128997 343571 129063 343574
rect 504725 343632 504834 343637
rect 504725 343576 504730 343632
rect 504786 343576 504834 343632
rect 504725 343574 504834 343576
rect 504725 343571 504791 343574
rect 70209 342002 70275 342005
rect 130285 342002 130351 342005
rect 70209 342000 130351 342002
rect 70209 341944 70214 342000
rect 70270 341944 130290 342000
rect 130346 341944 130351 342000
rect 70209 341942 130351 341944
rect 70209 341939 70275 341942
rect 130285 341939 130351 341942
rect 503713 340914 503779 340917
rect 503897 340914 503963 340917
rect 503713 340912 503963 340914
rect 503713 340856 503718 340912
rect 503774 340856 503902 340912
rect 503958 340856 503963 340912
rect 503713 340854 503963 340856
rect 503713 340851 503779 340854
rect 503897 340851 503963 340854
rect 237189 338738 237255 338741
rect 268142 338738 268148 338740
rect 237189 338736 268148 338738
rect 237189 338680 237194 338736
rect 237250 338680 268148 338736
rect 237189 338678 268148 338680
rect 237189 338675 237255 338678
rect 268142 338676 268148 338678
rect 268212 338676 268218 338740
rect 304165 338092 304231 338095
rect 304030 338090 304231 338092
rect 304030 338034 304170 338090
rect 304226 338034 304231 338090
rect 304030 338032 304231 338034
rect 304030 337922 304090 338032
rect 304165 338029 304231 338032
rect 304441 337922 304507 337925
rect 304030 337920 304507 337922
rect 304030 337864 304446 337920
rect 304502 337864 304507 337920
rect 304030 337862 304507 337864
rect 304441 337859 304507 337862
rect -960 337514 480 337604
rect 2957 337514 3023 337517
rect -960 337512 3023 337514
rect -960 337456 2962 337512
rect 3018 337456 3023 337512
rect -960 337454 3023 337456
rect -960 337364 480 337454
rect 2957 337451 3023 337454
rect 583520 334236 584960 334476
rect 504817 328674 504883 328677
rect 504222 328672 504883 328674
rect 504222 328616 504822 328672
rect 504878 328616 504883 328672
rect 504222 328614 504883 328616
rect 504222 328538 504282 328614
rect 504817 328611 504883 328614
rect 504357 328538 504423 328541
rect 504222 328536 504423 328538
rect 504222 328480 504362 328536
rect 504418 328480 504423 328536
rect 504222 328478 504423 328480
rect 504357 328475 504423 328478
rect -960 323098 480 323188
rect 3969 323098 4035 323101
rect -960 323096 4035 323098
rect -960 323040 3974 323096
rect 4030 323040 4035 323096
rect -960 323038 4035 323040
rect -960 322948 480 323038
rect 3969 323035 4035 323038
rect 579613 322690 579679 322693
rect 583520 322690 584960 322780
rect 579613 322688 584960 322690
rect 579613 322632 579618 322688
rect 579674 322632 584960 322688
rect 579613 322630 584960 322632
rect 579613 322627 579679 322630
rect 583520 322540 584960 322630
rect 257705 317388 257771 317389
rect 257654 317324 257660 317388
rect 257724 317386 257771 317388
rect 257724 317384 257816 317386
rect 257766 317328 257816 317384
rect 257724 317326 257816 317328
rect 257724 317324 257771 317326
rect 257705 317323 257771 317324
rect 257654 311748 257660 311812
rect 257724 311810 257730 311812
rect 257797 311810 257863 311813
rect 257724 311808 257863 311810
rect 257724 311752 257802 311808
rect 257858 311752 257863 311808
rect 257724 311750 257863 311752
rect 257724 311748 257730 311750
rect 257797 311747 257863 311750
rect 579705 310858 579771 310861
rect 583520 310858 584960 310948
rect 579705 310856 584960 310858
rect 579705 310800 579710 310856
rect 579766 310800 584960 310856
rect 579705 310798 584960 310800
rect 579705 310795 579771 310798
rect 583520 310708 584960 310798
rect -960 308818 480 308908
rect 4061 308818 4127 308821
rect -960 308816 4127 308818
rect -960 308760 4066 308816
rect 4122 308760 4127 308816
rect -960 308758 4127 308760
rect -960 308668 480 308758
rect 4061 308755 4127 308758
rect 128905 299434 128971 299437
rect 128905 299432 129106 299434
rect 128905 299376 128910 299432
rect 128966 299376 129106 299432
rect 128905 299374 129106 299376
rect 128905 299371 128971 299374
rect 128854 299236 128860 299300
rect 128924 299298 128930 299300
rect 129046 299298 129106 299374
rect 128924 299238 129106 299298
rect 128924 299236 128930 299238
rect 580625 299162 580691 299165
rect 583520 299162 584960 299252
rect 580625 299160 584960 299162
rect 580625 299104 580630 299160
rect 580686 299104 584960 299160
rect 580625 299102 584960 299104
rect 580625 299099 580691 299102
rect 583520 299012 584960 299102
rect -960 294402 480 294492
rect 3325 294402 3391 294405
rect -960 294400 3391 294402
rect -960 294344 3330 294400
rect 3386 294344 3391 294400
rect -960 294342 3391 294344
rect -960 294252 480 294342
rect 3325 294339 3391 294342
rect 128813 289916 128879 289917
rect 128813 289912 128860 289916
rect 128924 289914 128930 289916
rect 128813 289856 128818 289912
rect 128813 289852 128860 289856
rect 128924 289854 128970 289914
rect 128924 289852 128930 289854
rect 128813 289851 128879 289852
rect 583520 287316 584960 287556
rect -960 280122 480 280212
rect 4061 280122 4127 280125
rect -960 280120 4127 280122
rect -960 280064 4066 280120
rect 4122 280064 4127 280120
rect -960 280062 4127 280064
rect -960 279972 480 280062
rect 4061 280059 4127 280062
rect 128905 280122 128971 280125
rect 128905 280120 129106 280122
rect 128905 280064 128910 280120
rect 128966 280064 129106 280120
rect 128905 280062 129106 280064
rect 128905 280059 128971 280062
rect 129046 279989 129106 280062
rect 128997 279984 129106 279989
rect 128997 279928 129002 279984
rect 129058 279928 129106 279984
rect 128997 279926 129106 279928
rect 128997 279923 129063 279926
rect 579613 275770 579679 275773
rect 583520 275770 584960 275860
rect 579613 275768 584960 275770
rect 579613 275712 579618 275768
rect 579674 275712 584960 275768
rect 579613 275710 584960 275712
rect 579613 275707 579679 275710
rect 583520 275620 584960 275710
rect -960 265706 480 265796
rect 2773 265706 2839 265709
rect -960 265704 2839 265706
rect -960 265648 2778 265704
rect 2834 265648 2839 265704
rect -960 265646 2839 265648
rect -960 265556 480 265646
rect 2773 265643 2839 265646
rect 580165 263938 580231 263941
rect 583520 263938 584960 264028
rect 580165 263936 584960 263938
rect 580165 263880 580170 263936
rect 580226 263880 584960 263936
rect 580165 263878 584960 263880
rect 580165 263875 580231 263878
rect 583520 263788 584960 263878
rect 304073 260946 304139 260949
rect 304441 260946 304507 260949
rect 304073 260944 304507 260946
rect 304073 260888 304078 260944
rect 304134 260888 304446 260944
rect 304502 260888 304507 260944
rect 304073 260886 304507 260888
rect 304073 260883 304139 260886
rect 304441 260883 304507 260886
rect 504265 260946 504331 260949
rect 504633 260946 504699 260949
rect 504265 260944 504699 260946
rect 504265 260888 504270 260944
rect 504326 260888 504638 260944
rect 504694 260888 504699 260944
rect 504265 260886 504699 260888
rect 504265 260883 504331 260886
rect 504633 260883 504699 260886
rect 580717 252242 580783 252245
rect 583520 252242 584960 252332
rect 580717 252240 584960 252242
rect 580717 252184 580722 252240
rect 580778 252184 584960 252240
rect 580717 252182 584960 252184
rect 580717 252179 580783 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3325 251290 3391 251293
rect -960 251288 3391 251290
rect -960 251232 3330 251288
rect 3386 251232 3391 251288
rect -960 251230 3391 251232
rect -960 251140 480 251230
rect 3325 251227 3391 251230
rect 209773 241498 209839 241501
rect 209957 241498 210023 241501
rect 209773 241496 210023 241498
rect 209773 241440 209778 241496
rect 209834 241440 209962 241496
rect 210018 241440 210023 241496
rect 209773 241438 210023 241440
rect 209773 241435 209839 241438
rect 209957 241435 210023 241438
rect 583520 240396 584960 240636
rect -960 237010 480 237100
rect 3325 237010 3391 237013
rect -960 237008 3391 237010
rect -960 236952 3330 237008
rect 3386 236952 3391 237008
rect -960 236950 3391 236952
rect -960 236860 480 236950
rect 3325 236947 3391 236950
rect 288249 231842 288315 231845
rect 288525 231842 288591 231845
rect 288249 231840 288591 231842
rect 288249 231784 288254 231840
rect 288310 231784 288530 231840
rect 288586 231784 288591 231840
rect 288249 231782 288591 231784
rect 288249 231779 288315 231782
rect 288525 231779 288591 231782
rect 304257 231842 304323 231845
rect 304533 231842 304599 231845
rect 304257 231840 304599 231842
rect 304257 231784 304262 231840
rect 304318 231784 304538 231840
rect 304594 231784 304599 231840
rect 304257 231782 304599 231784
rect 304257 231779 304323 231782
rect 304533 231779 304599 231782
rect 580165 228850 580231 228853
rect 583520 228850 584960 228940
rect 580165 228848 584960 228850
rect 580165 228792 580170 228848
rect 580226 228792 584960 228848
rect 580165 228790 584960 228792
rect 580165 228787 580231 228790
rect 583520 228700 584960 228790
rect -960 222594 480 222684
rect 2957 222594 3023 222597
rect -960 222592 3023 222594
rect -960 222536 2962 222592
rect 3018 222536 3023 222592
rect -960 222534 3023 222536
rect -960 222444 480 222534
rect 2957 222531 3023 222534
rect 209773 222186 209839 222189
rect 209957 222186 210023 222189
rect 209773 222184 210023 222186
rect 209773 222128 209778 222184
rect 209834 222128 209962 222184
rect 210018 222128 210023 222184
rect 209773 222126 210023 222128
rect 209773 222123 209839 222126
rect 209957 222123 210023 222126
rect 257797 220826 257863 220829
rect 257981 220826 258047 220829
rect 257797 220824 258047 220826
rect 257797 220768 257802 220824
rect 257858 220768 257986 220824
rect 258042 220768 258047 220824
rect 257797 220766 258047 220768
rect 257797 220763 257863 220766
rect 257981 220763 258047 220766
rect 579613 217018 579679 217021
rect 583520 217018 584960 217108
rect 579613 217016 584960 217018
rect 579613 216960 579618 217016
rect 579674 216960 584960 217016
rect 579613 216958 584960 216960
rect 579613 216955 579679 216958
rect 583520 216868 584960 216958
rect -960 208178 480 208268
rect 2957 208178 3023 208181
rect -960 208176 3023 208178
rect -960 208120 2962 208176
rect 3018 208120 3023 208176
rect -960 208118 3023 208120
rect -960 208028 480 208118
rect 2957 208115 3023 208118
rect 580809 205322 580875 205325
rect 583520 205322 584960 205412
rect 580809 205320 584960 205322
rect 580809 205264 580814 205320
rect 580870 205264 584960 205320
rect 580809 205262 584960 205264
rect 580809 205259 580875 205262
rect 583520 205172 584960 205262
rect 197077 202874 197143 202877
rect 220353 202874 220419 202877
rect 197077 202872 220419 202874
rect 197077 202816 197082 202872
rect 197138 202816 220358 202872
rect 220414 202816 220419 202872
rect 197077 202814 220419 202816
rect 197077 202811 197143 202814
rect 220353 202811 220419 202814
rect 196985 202738 197051 202741
rect 223849 202738 223915 202741
rect 196985 202736 223915 202738
rect 196985 202680 196990 202736
rect 197046 202680 223854 202736
rect 223910 202680 223915 202736
rect 196985 202678 223915 202680
rect 196985 202675 197051 202678
rect 223849 202675 223915 202678
rect 197854 202540 197860 202604
rect 197924 202602 197930 202604
rect 225137 202602 225203 202605
rect 197924 202600 225203 202602
rect 197924 202544 225142 202600
rect 225198 202544 225203 202600
rect 197924 202542 225203 202544
rect 197924 202540 197930 202542
rect 225137 202539 225203 202542
rect 197261 202466 197327 202469
rect 226333 202466 226399 202469
rect 197261 202464 226399 202466
rect 197261 202408 197266 202464
rect 197322 202408 226338 202464
rect 226394 202408 226399 202464
rect 197261 202406 226399 202408
rect 197261 202403 197327 202406
rect 226333 202403 226399 202406
rect 198222 202268 198228 202332
rect 198292 202330 198298 202332
rect 232129 202330 232195 202333
rect 198292 202328 232195 202330
rect 198292 202272 232134 202328
rect 232190 202272 232195 202328
rect 198292 202270 232195 202272
rect 198292 202268 198298 202270
rect 232129 202267 232195 202270
rect 197169 202194 197235 202197
rect 233417 202194 233483 202197
rect 197169 202192 233483 202194
rect 197169 202136 197174 202192
rect 197230 202136 233422 202192
rect 233478 202136 233483 202192
rect 197169 202134 233483 202136
rect 197169 202131 197235 202134
rect 233417 202131 233483 202134
rect 257061 202194 257127 202197
rect 267958 202194 267964 202196
rect 257061 202192 267964 202194
rect 257061 202136 257066 202192
rect 257122 202136 267964 202192
rect 257061 202134 267964 202136
rect 257061 202131 257127 202134
rect 267958 202132 267964 202134
rect 268028 202132 268034 202196
rect 199694 201996 199700 202060
rect 199764 202058 199770 202060
rect 218053 202058 218119 202061
rect 199764 202056 218119 202058
rect 199764 202000 218058 202056
rect 218114 202000 218119 202056
rect 199764 201998 218119 202000
rect 199764 201996 199770 201998
rect 218053 201995 218119 201998
rect 198406 201860 198412 201924
rect 198476 201922 198482 201924
rect 212533 201922 212599 201925
rect 198476 201920 212599 201922
rect 198476 201864 212538 201920
rect 212594 201864 212599 201920
rect 198476 201862 212599 201864
rect 198476 201860 198482 201862
rect 212533 201859 212599 201862
rect 232405 201922 232471 201925
rect 238661 201922 238727 201925
rect 232405 201920 238727 201922
rect 232405 201864 232410 201920
rect 232466 201864 238666 201920
rect 238722 201864 238727 201920
rect 232405 201862 238727 201864
rect 232405 201859 232471 201862
rect 238661 201859 238727 201862
rect 198590 201724 198596 201788
rect 198660 201786 198666 201788
rect 213453 201786 213519 201789
rect 198660 201784 213519 201786
rect 198660 201728 213458 201784
rect 213514 201728 213519 201784
rect 198660 201726 213519 201728
rect 198660 201724 198666 201726
rect 213453 201723 213519 201726
rect 198038 201588 198044 201652
rect 198108 201650 198114 201652
rect 211153 201650 211219 201653
rect 198108 201648 211219 201650
rect 198108 201592 211158 201648
rect 211214 201592 211219 201648
rect 198108 201590 211219 201592
rect 198108 201588 198114 201590
rect 211153 201587 211219 201590
rect 262673 201650 262739 201653
rect 267774 201650 267780 201652
rect 262673 201648 267780 201650
rect 262673 201592 262678 201648
rect 262734 201592 267780 201648
rect 262673 201590 267780 201592
rect 262673 201587 262739 201590
rect 267774 201588 267780 201590
rect 267844 201588 267850 201652
rect 266169 201514 266235 201517
rect 266854 201514 266860 201516
rect 266169 201512 266860 201514
rect 266169 201456 266174 201512
rect 266230 201456 266860 201512
rect 266169 201454 266860 201456
rect 266169 201451 266235 201454
rect 266854 201452 266860 201454
rect 266924 201452 266930 201516
rect 132902 200636 132908 200700
rect 132972 200698 132978 200700
rect 527173 200698 527239 200701
rect 132972 200696 527239 200698
rect 132972 200640 527178 200696
rect 527234 200640 527239 200696
rect 132972 200638 527239 200640
rect 132972 200636 132978 200638
rect 527173 200635 527239 200638
rect 131757 199338 131823 199341
rect 131757 199336 134044 199338
rect 131757 199280 131762 199336
rect 131818 199280 134044 199336
rect 131757 199278 134044 199280
rect 131757 199275 131823 199278
rect 436185 198930 436251 198933
rect 433934 198928 436251 198930
rect 433934 198872 436190 198928
rect 436246 198872 436251 198928
rect 433934 198870 436251 198872
rect 433934 198764 433994 198870
rect 436185 198867 436251 198870
rect 131389 198250 131455 198253
rect 131389 198248 134044 198250
rect 131389 198192 131394 198248
rect 131450 198192 134044 198248
rect 131389 198190 134044 198192
rect 131389 198187 131455 198190
rect 131389 197162 131455 197165
rect 131389 197160 134044 197162
rect 131389 197104 131394 197160
rect 131450 197104 134044 197160
rect 131389 197102 134044 197104
rect 131389 197099 131455 197102
rect 130469 196210 130535 196213
rect 433934 196210 433994 196724
rect 434989 196210 435055 196213
rect 130469 196208 134044 196210
rect 130469 196152 130474 196208
rect 130530 196152 134044 196208
rect 130469 196150 134044 196152
rect 433934 196208 435055 196210
rect 433934 196152 434994 196208
rect 435050 196152 435055 196208
rect 433934 196150 435055 196152
rect 130469 196147 130535 196150
rect 434989 196147 435055 196150
rect 130469 194714 130535 194717
rect 134014 194714 134074 195092
rect 130469 194712 134074 194714
rect 130469 194656 130474 194712
rect 130530 194656 134074 194712
rect 130469 194654 134074 194656
rect 130469 194651 130535 194654
rect 130469 194442 130535 194445
rect 130469 194440 134074 194442
rect 130469 194384 130474 194440
rect 130530 194384 134074 194440
rect 130469 194382 134074 194384
rect 130469 194379 130535 194382
rect 134014 194004 134074 194382
rect 433934 194034 433994 194548
rect 436277 194034 436343 194037
rect 433934 194032 436343 194034
rect -960 193898 480 193988
rect 433934 193976 436282 194032
rect 436338 193976 436343 194032
rect 433934 193974 436343 193976
rect 436277 193971 436343 193974
rect 3601 193898 3667 193901
rect -960 193896 3667 193898
rect -960 193840 3606 193896
rect 3662 193840 3667 193896
rect -960 193838 3667 193840
rect -960 193748 480 193838
rect 3601 193835 3667 193838
rect 583520 193476 584960 193716
rect 130469 193082 130535 193085
rect 436645 193082 436711 193085
rect 130469 193080 134074 193082
rect 130469 193024 130474 193080
rect 130530 193024 134074 193080
rect 130469 193022 134074 193024
rect 130469 193019 130535 193022
rect 134014 192916 134074 193022
rect 433934 193080 436711 193082
rect 433934 193024 436650 193080
rect 436706 193024 436711 193080
rect 433934 193022 436711 193024
rect 130377 192538 130443 192541
rect 130377 192536 134074 192538
rect 130377 192480 130382 192536
rect 130438 192480 134074 192536
rect 433934 192508 433994 193022
rect 436645 193019 436711 193022
rect 130377 192478 134074 192480
rect 130377 192475 130443 192478
rect 134014 191964 134074 192478
rect 130469 191450 130535 191453
rect 130469 191448 134074 191450
rect 130469 191392 130474 191448
rect 130530 191392 134074 191448
rect 130469 191390 134074 191392
rect 130469 191387 130535 191390
rect 134014 190876 134074 191390
rect 128537 190498 128603 190501
rect 128721 190498 128787 190501
rect 128537 190496 128787 190498
rect 128537 190440 128542 190496
rect 128598 190440 128726 190496
rect 128782 190440 128787 190496
rect 128537 190438 128787 190440
rect 128537 190435 128603 190438
rect 128721 190435 128787 190438
rect 130469 190362 130535 190365
rect 130469 190360 134074 190362
rect 130469 190304 130474 190360
rect 130530 190304 134074 190360
rect 130469 190302 134074 190304
rect 130469 190299 130535 190302
rect 134014 189788 134074 190302
rect 433934 190226 433994 190332
rect 435173 190226 435239 190229
rect 433934 190224 435239 190226
rect 433934 190168 435178 190224
rect 435234 190168 435239 190224
rect 433934 190166 435239 190168
rect 435173 190163 435239 190166
rect 130469 188866 130535 188869
rect 435081 188866 435147 188869
rect 130469 188864 134074 188866
rect 130469 188808 130474 188864
rect 130530 188808 134074 188864
rect 130469 188806 134074 188808
rect 130469 188803 130535 188806
rect 134014 188700 134074 188806
rect 433934 188864 435147 188866
rect 433934 188808 435086 188864
rect 435142 188808 435147 188864
rect 433934 188806 435147 188808
rect 130377 188322 130443 188325
rect 130377 188320 134074 188322
rect 130377 188264 130382 188320
rect 130438 188264 134074 188320
rect 433934 188292 433994 188806
rect 435081 188803 435147 188806
rect 130377 188262 134074 188264
rect 130377 188259 130443 188262
rect 134014 187748 134074 188262
rect 130469 187234 130535 187237
rect 130469 187232 134074 187234
rect 130469 187176 130474 187232
rect 130530 187176 134074 187232
rect 130469 187174 134074 187176
rect 130469 187171 130535 187174
rect 134014 186660 134074 187174
rect 434529 186282 434595 186285
rect 433934 186280 434595 186282
rect 433934 186224 434534 186280
rect 434590 186224 434595 186280
rect 433934 186222 434595 186224
rect 433934 186116 433994 186222
rect 434529 186219 434595 186222
rect 131205 185602 131271 185605
rect 131205 185600 134044 185602
rect 131205 185544 131210 185600
rect 131266 185544 134044 185600
rect 131205 185542 134044 185544
rect 131205 185539 131271 185542
rect 434897 184650 434963 184653
rect 433934 184648 434963 184650
rect 433934 184592 434902 184648
rect 434958 184592 434963 184648
rect 433934 184590 434963 184592
rect 131205 184514 131271 184517
rect 131205 184512 134044 184514
rect 131205 184456 131210 184512
rect 131266 184456 134044 184512
rect 131205 184454 134044 184456
rect 131205 184451 131271 184454
rect 433934 184076 433994 184590
rect 434897 184587 434963 184590
rect 131205 183562 131271 183565
rect 504357 183562 504423 183565
rect 504633 183562 504699 183565
rect 131205 183560 134044 183562
rect 131205 183504 131210 183560
rect 131266 183504 134044 183560
rect 131205 183502 134044 183504
rect 504357 183560 504699 183562
rect 504357 183504 504362 183560
rect 504418 183504 504638 183560
rect 504694 183504 504699 183560
rect 504357 183502 504699 183504
rect 131205 183499 131271 183502
rect 504357 183499 504423 183502
rect 504633 183499 504699 183502
rect 133321 182474 133387 182477
rect 133321 182472 134044 182474
rect 133321 182416 133326 182472
rect 133382 182416 134044 182472
rect 133321 182414 134044 182416
rect 133321 182411 133387 182414
rect 126513 182202 126579 182205
rect 126789 182202 126855 182205
rect 126513 182200 126855 182202
rect 126513 182144 126518 182200
rect 126574 182144 126794 182200
rect 126850 182144 126855 182200
rect 126513 182142 126855 182144
rect 126513 182139 126579 182142
rect 126789 182139 126855 182142
rect 436553 182066 436619 182069
rect 433934 182064 436619 182066
rect 433934 182008 436558 182064
rect 436614 182008 436619 182064
rect 433934 182006 436619 182008
rect 433934 181900 433994 182006
rect 436553 182003 436619 182006
rect 580257 181930 580323 181933
rect 583520 181930 584960 182020
rect 580257 181928 584960 181930
rect 580257 181872 580262 181928
rect 580318 181872 584960 181928
rect 580257 181870 584960 181872
rect 580257 181867 580323 181870
rect 583520 181780 584960 181870
rect 133413 181386 133479 181389
rect 133413 181384 134044 181386
rect 133413 181328 133418 181384
rect 133474 181328 134044 181384
rect 133413 181326 134044 181328
rect 133413 181323 133479 181326
rect 133965 180706 134031 180709
rect 133965 180704 134074 180706
rect 133965 180648 133970 180704
rect 134026 180648 134074 180704
rect 133965 180643 134074 180648
rect 134014 180404 134074 180643
rect 436093 180298 436159 180301
rect 433934 180296 436159 180298
rect 433934 180240 436098 180296
rect 436154 180240 436159 180296
rect 433934 180238 436159 180240
rect 433934 179860 433994 180238
rect 436093 180235 436159 180238
rect -960 179482 480 179572
rect 2865 179482 2931 179485
rect -960 179480 2931 179482
rect -960 179424 2870 179480
rect 2926 179424 2931 179480
rect -960 179422 2931 179424
rect -960 179332 480 179422
rect 2865 179419 2931 179422
rect 132493 179346 132559 179349
rect 132493 179344 134044 179346
rect 132493 179288 132498 179344
rect 132554 179288 134044 179344
rect 132493 179286 134044 179288
rect 132493 179283 132559 179286
rect 131205 178258 131271 178261
rect 131205 178256 134044 178258
rect 131205 178200 131210 178256
rect 131266 178200 134044 178256
rect 131205 178198 134044 178200
rect 131205 178195 131271 178198
rect 436461 177986 436527 177989
rect 433934 177984 436527 177986
rect 433934 177928 436466 177984
rect 436522 177928 436527 177984
rect 433934 177926 436527 177928
rect 433934 177684 433994 177926
rect 436461 177923 436527 177926
rect 132585 177170 132651 177173
rect 132585 177168 134044 177170
rect 132585 177112 132590 177168
rect 132646 177112 134044 177168
rect 132585 177110 134044 177112
rect 132585 177107 132651 177110
rect 132902 176156 132908 176220
rect 132972 176218 132978 176220
rect 436369 176218 436435 176221
rect 132972 176158 134044 176218
rect 433934 176216 436435 176218
rect 433934 176160 436374 176216
rect 436430 176160 436435 176216
rect 433934 176158 436435 176160
rect 132972 176156 132978 176158
rect 433934 175644 433994 176158
rect 436369 176155 436435 176158
rect 133638 175068 133644 175132
rect 133708 175130 133714 175132
rect 133708 175070 134044 175130
rect 133708 175068 133714 175070
rect 133454 173980 133460 174044
rect 133524 174042 133530 174044
rect 133524 173982 134044 174042
rect 133524 173980 133530 173982
rect 434805 173906 434871 173909
rect 433934 173904 434871 173906
rect 433934 173848 434810 173904
rect 434866 173848 434871 173904
rect 433934 173846 434871 173848
rect 433934 173468 433994 173846
rect 434805 173843 434871 173846
rect 133086 172892 133092 172956
rect 133156 172954 133162 172956
rect 133156 172894 134044 172954
rect 133156 172892 133162 172894
rect 132401 172002 132467 172005
rect 434713 172002 434779 172005
rect 132401 172000 134044 172002
rect 132401 171944 132406 172000
rect 132462 171944 134044 172000
rect 132401 171942 134044 171944
rect 433934 172000 434779 172002
rect 433934 171944 434718 172000
rect 434774 171944 434779 172000
rect 433934 171942 434779 171944
rect 132401 171939 132467 171942
rect 433934 171428 433994 171942
rect 434713 171939 434779 171942
rect 132217 170914 132283 170917
rect 132217 170912 134044 170914
rect 132217 170856 132222 170912
rect 132278 170856 134044 170912
rect 132217 170854 134044 170856
rect 132217 170851 132283 170854
rect 580257 170098 580323 170101
rect 583520 170098 584960 170188
rect 580257 170096 584960 170098
rect 580257 170040 580262 170096
rect 580318 170040 584960 170096
rect 580257 170038 584960 170040
rect 580257 170035 580323 170038
rect 583520 169948 584960 170038
rect 133137 169826 133203 169829
rect 133137 169824 134044 169826
rect 133137 169768 133142 169824
rect 133198 169768 134044 169824
rect 133137 169766 134044 169768
rect 133137 169763 133203 169766
rect 434253 169690 434319 169693
rect 433934 169688 434319 169690
rect 433934 169632 434258 169688
rect 434314 169632 434319 169688
rect 433934 169630 434319 169632
rect 433934 169252 433994 169630
rect 434253 169627 434319 169630
rect 132953 168738 133019 168741
rect 132953 168736 134044 168738
rect 132953 168680 132958 168736
rect 133014 168680 134044 168736
rect 132953 168678 134044 168680
rect 132953 168675 133019 168678
rect 131665 167786 131731 167789
rect 434437 167786 434503 167789
rect 131665 167784 134044 167786
rect 131665 167728 131670 167784
rect 131726 167728 134044 167784
rect 131665 167726 134044 167728
rect 433934 167784 434503 167786
rect 433934 167728 434442 167784
rect 434498 167728 434503 167784
rect 433934 167726 434503 167728
rect 131665 167723 131731 167726
rect 433934 167212 433994 167726
rect 434437 167723 434503 167726
rect 132769 166698 132835 166701
rect 132769 166696 134044 166698
rect 132769 166640 132774 166696
rect 132830 166640 134044 166696
rect 132769 166638 134044 166640
rect 132769 166635 132835 166638
rect 132677 165610 132743 165613
rect 434345 165610 434411 165613
rect 132677 165608 134044 165610
rect 132677 165552 132682 165608
rect 132738 165552 134044 165608
rect 132677 165550 134044 165552
rect 433934 165608 434411 165610
rect 433934 165552 434350 165608
rect 434406 165552 434411 165608
rect 433934 165550 434411 165552
rect 132677 165547 132743 165550
rect -960 165066 480 165156
rect 3233 165066 3299 165069
rect -960 165064 3299 165066
rect -960 165008 3238 165064
rect 3294 165008 3299 165064
rect 433934 165036 433994 165550
rect 434345 165547 434411 165550
rect -960 165006 3299 165008
rect -960 164916 480 165006
rect 3233 165003 3299 165006
rect 131297 164522 131363 164525
rect 131297 164520 134044 164522
rect 131297 164464 131302 164520
rect 131358 164464 134044 164520
rect 131297 164462 134044 164464
rect 131297 164459 131363 164462
rect 133597 163570 133663 163573
rect 434161 163570 434227 163573
rect 133597 163568 134044 163570
rect 133597 163512 133602 163568
rect 133658 163512 134044 163568
rect 133597 163510 134044 163512
rect 433934 163568 434227 163570
rect 433934 163512 434166 163568
rect 434222 163512 434227 163568
rect 433934 163510 434227 163512
rect 133597 163507 133663 163510
rect 433934 162996 433994 163510
rect 434161 163507 434227 163510
rect 132401 162482 132467 162485
rect 132401 162480 134044 162482
rect 132401 162424 132406 162480
rect 132462 162424 134044 162480
rect 132401 162422 134044 162424
rect 132401 162419 132467 162422
rect 131205 161394 131271 161397
rect 131205 161392 134044 161394
rect 131205 161336 131210 161392
rect 131266 161336 134044 161392
rect 131205 161334 134044 161336
rect 131205 161331 131271 161334
rect 434069 161258 434135 161261
rect 433934 161256 434135 161258
rect 433934 161200 434074 161256
rect 434130 161200 434135 161256
rect 433934 161198 434135 161200
rect 433934 160956 433994 161198
rect 434069 161195 434135 161198
rect 133597 160442 133663 160445
rect 133597 160440 134044 160442
rect 133597 160384 133602 160440
rect 133658 160384 134044 160440
rect 133597 160382 134044 160384
rect 133597 160379 133663 160382
rect 132217 159354 132283 159357
rect 433977 159354 434043 159357
rect 132217 159352 134044 159354
rect 132217 159296 132222 159352
rect 132278 159296 134044 159352
rect 132217 159294 134044 159296
rect 433934 159352 434043 159354
rect 433934 159296 433982 159352
rect 434038 159296 434043 159352
rect 132217 159291 132283 159294
rect 433934 159291 434043 159296
rect 433934 158780 433994 159291
rect 580165 158402 580231 158405
rect 583520 158402 584960 158492
rect 580165 158400 584960 158402
rect 580165 158344 580170 158400
rect 580226 158344 584960 158400
rect 580165 158342 584960 158344
rect 580165 158339 580231 158342
rect 131665 158266 131731 158269
rect 131665 158264 134044 158266
rect 131665 158208 131670 158264
rect 131726 158208 134044 158264
rect 583520 158252 584960 158342
rect 131665 158206 134044 158208
rect 131665 158203 131731 158206
rect 433885 157314 433951 157317
rect 433885 157312 433994 157314
rect 433885 157256 433890 157312
rect 433946 157256 433994 157312
rect 433885 157251 433994 157256
rect 131297 157178 131363 157181
rect 131297 157176 134044 157178
rect 131297 157120 131302 157176
rect 131358 157120 134044 157176
rect 131297 157118 134044 157120
rect 131297 157115 131363 157118
rect 433934 156740 433994 157251
rect 131113 156226 131179 156229
rect 131113 156224 134044 156226
rect 131113 156168 131118 156224
rect 131174 156168 134044 156224
rect 131113 156166 134044 156168
rect 131113 156163 131179 156166
rect 131113 155138 131179 155141
rect 436093 155138 436159 155141
rect 131113 155136 134044 155138
rect 131113 155080 131118 155136
rect 131174 155080 134044 155136
rect 131113 155078 134044 155080
rect 433934 155136 436159 155138
rect 433934 155080 436098 155136
rect 436154 155080 436159 155136
rect 433934 155078 436159 155080
rect 131113 155075 131179 155078
rect 433934 154564 433994 155078
rect 436093 155075 436159 155078
rect 504173 154594 504239 154597
rect 504449 154594 504515 154597
rect 504173 154592 504515 154594
rect 504173 154536 504178 154592
rect 504234 154536 504454 154592
rect 504510 154536 504515 154592
rect 504173 154534 504515 154536
rect 504173 154531 504239 154534
rect 504449 154531 504515 154534
rect 124213 154050 124279 154053
rect 124213 154048 134044 154050
rect 124213 153992 124218 154048
rect 124274 153992 134044 154048
rect 124213 153990 134044 153992
rect 124213 153987 124279 153990
rect 126421 153234 126487 153237
rect 126421 153232 126530 153234
rect 126421 153176 126426 153232
rect 126482 153176 126530 153232
rect 126421 153171 126530 153176
rect 126470 153098 126530 153171
rect 126697 153098 126763 153101
rect 126470 153096 126763 153098
rect 126470 153040 126702 153096
rect 126758 153040 126763 153096
rect 126470 153038 126763 153040
rect 126697 153035 126763 153038
rect 131113 152962 131179 152965
rect 131113 152960 134044 152962
rect 131113 152904 131118 152960
rect 131174 152904 134044 152960
rect 131113 152902 134044 152904
rect 131113 152899 131179 152902
rect 437381 152826 437447 152829
rect 433934 152824 437447 152826
rect 433934 152768 437386 152824
rect 437442 152768 437447 152824
rect 433934 152766 437447 152768
rect 433934 152524 433994 152766
rect 437381 152763 437447 152766
rect 131205 152010 131271 152013
rect 131205 152008 134044 152010
rect 131205 151952 131210 152008
rect 131266 151952 134044 152008
rect 131205 151950 134044 151952
rect 131205 151947 131271 151950
rect 131113 150922 131179 150925
rect 131113 150920 134044 150922
rect -960 150786 480 150876
rect 131113 150864 131118 150920
rect 131174 150864 134044 150920
rect 131113 150862 134044 150864
rect 131113 150859 131179 150862
rect 3233 150786 3299 150789
rect -960 150784 3299 150786
rect -960 150728 3238 150784
rect 3294 150728 3299 150784
rect -960 150726 3299 150728
rect -960 150636 480 150726
rect 3233 150723 3299 150726
rect 433934 150242 433994 150348
rect 437381 150242 437447 150245
rect 433934 150240 437447 150242
rect 433934 150184 437386 150240
rect 437442 150184 437447 150240
rect 433934 150182 437447 150184
rect 437381 150179 437447 150182
rect 131113 149834 131179 149837
rect 131113 149832 134044 149834
rect 131113 149776 131118 149832
rect 131174 149776 134044 149832
rect 131113 149774 134044 149776
rect 131113 149771 131179 149774
rect 131113 148746 131179 148749
rect 436093 148746 436159 148749
rect 131113 148744 134044 148746
rect 131113 148688 131118 148744
rect 131174 148688 134044 148744
rect 131113 148686 134044 148688
rect 433934 148744 436159 148746
rect 433934 148688 436098 148744
rect 436154 148688 436159 148744
rect 433934 148686 436159 148688
rect 131113 148683 131179 148686
rect 433934 148308 433994 148686
rect 436093 148683 436159 148686
rect 131113 147794 131179 147797
rect 131113 147792 134044 147794
rect 131113 147736 131118 147792
rect 131174 147736 134044 147792
rect 131113 147734 134044 147736
rect 131113 147731 131179 147734
rect 131113 146706 131179 146709
rect 131113 146704 134044 146706
rect 131113 146648 131118 146704
rect 131174 146648 134044 146704
rect 131113 146646 134044 146648
rect 131113 146643 131179 146646
rect 583520 146556 584960 146796
rect 437381 146298 437447 146301
rect 433934 146296 437447 146298
rect 433934 146240 437386 146296
rect 437442 146240 437447 146296
rect 433934 146238 437447 146240
rect 433934 146132 433994 146238
rect 437381 146235 437447 146238
rect 131113 145618 131179 145621
rect 131113 145616 134044 145618
rect 131113 145560 131118 145616
rect 131174 145560 134044 145616
rect 131113 145558 134044 145560
rect 131113 145555 131179 145558
rect 128169 144530 128235 144533
rect 437013 144530 437079 144533
rect 128169 144528 134044 144530
rect 128169 144472 128174 144528
rect 128230 144472 134044 144528
rect 128169 144470 134044 144472
rect 433934 144528 437079 144530
rect 433934 144472 437018 144528
rect 437074 144472 437079 144528
rect 433934 144470 437079 144472
rect 128169 144467 128235 144470
rect 433934 144092 433994 144470
rect 437013 144467 437079 144470
rect 126513 143578 126579 143581
rect 126697 143578 126763 143581
rect 126513 143576 126763 143578
rect 126513 143520 126518 143576
rect 126574 143520 126702 143576
rect 126758 143520 126763 143576
rect 126513 143518 126763 143520
rect 126513 143515 126579 143518
rect 126697 143515 126763 143518
rect 131113 143578 131179 143581
rect 131113 143576 134044 143578
rect 131113 143520 131118 143576
rect 131174 143520 134044 143576
rect 131113 143518 134044 143520
rect 131113 143515 131179 143518
rect 133505 142490 133571 142493
rect 133505 142488 134044 142490
rect 133505 142432 133510 142488
rect 133566 142432 134044 142488
rect 133505 142430 134044 142432
rect 133505 142427 133571 142430
rect 436093 142082 436159 142085
rect 433934 142080 436159 142082
rect 433934 142024 436098 142080
rect 436154 142024 436159 142080
rect 433934 142022 436159 142024
rect 433934 141916 433994 142022
rect 436093 142019 436159 142022
rect 133689 141402 133755 141405
rect 133689 141400 134044 141402
rect 133689 141344 133694 141400
rect 133750 141344 134044 141400
rect 133689 141342 134044 141344
rect 133689 141339 133755 141342
rect 133781 140450 133847 140453
rect 436737 140450 436803 140453
rect 133781 140448 134044 140450
rect 133781 140392 133786 140448
rect 133842 140392 134044 140448
rect 133781 140390 134044 140392
rect 433934 140448 436803 140450
rect 433934 140392 436742 140448
rect 436798 140392 436803 140448
rect 433934 140390 436803 140392
rect 133781 140387 133847 140390
rect 433934 139876 433994 140390
rect 436737 140387 436803 140390
rect 131297 139362 131363 139365
rect 131297 139360 134044 139362
rect 131297 139304 131302 139360
rect 131358 139304 134044 139360
rect 131297 139302 134044 139304
rect 131297 139299 131363 139302
rect 132309 138274 132375 138277
rect 132309 138272 134044 138274
rect 132309 138216 132314 138272
rect 132370 138216 134044 138272
rect 132309 138214 134044 138216
rect 132309 138211 132375 138214
rect 437381 137866 437447 137869
rect 433934 137864 437447 137866
rect 433934 137808 437386 137864
rect 437442 137808 437447 137864
rect 433934 137806 437447 137808
rect 433934 137700 433994 137806
rect 437381 137803 437447 137806
rect 132166 137124 132172 137188
rect 132236 137186 132242 137188
rect 132236 137126 134044 137186
rect 132236 137124 132242 137126
rect -960 136370 480 136460
rect 3325 136370 3391 136373
rect -960 136368 3391 136370
rect -960 136312 3330 136368
rect 3386 136312 3391 136368
rect -960 136310 3391 136312
rect -960 136220 480 136310
rect 3325 136307 3391 136310
rect 132350 136172 132356 136236
rect 132420 136234 132426 136236
rect 132420 136174 134044 136234
rect 132420 136172 132426 136174
rect 437013 136098 437079 136101
rect 433934 136096 437079 136098
rect 433934 136040 437018 136096
rect 437074 136040 437079 136096
rect 433934 136038 437079 136040
rect 433934 135660 433994 136038
rect 437013 136035 437079 136038
rect 131982 135084 131988 135148
rect 132052 135146 132058 135148
rect 132052 135086 134044 135146
rect 132052 135084 132058 135086
rect 580349 134874 580415 134877
rect 583520 134874 584960 134964
rect 580349 134872 584960 134874
rect 580349 134816 580354 134872
rect 580410 134816 584960 134872
rect 580349 134814 584960 134816
rect 580349 134811 580415 134814
rect 583520 134724 584960 134814
rect 131798 133996 131804 134060
rect 131868 134058 131874 134060
rect 131868 133998 134044 134058
rect 131868 133996 131874 133998
rect 437381 133650 437447 133653
rect 433934 133648 437447 133650
rect 433934 133592 437386 133648
rect 437442 133592 437447 133648
rect 433934 133590 437447 133592
rect 433934 133484 433994 133590
rect 437381 133587 437447 133590
rect 133270 132908 133276 132972
rect 133340 132970 133346 132972
rect 133340 132910 134044 132970
rect 133340 132908 133346 132910
rect 131389 132018 131455 132021
rect 437381 132018 437447 132021
rect 131389 132016 134044 132018
rect 131389 131960 131394 132016
rect 131450 131960 134044 132016
rect 131389 131958 134044 131960
rect 433934 132016 437447 132018
rect 433934 131960 437386 132016
rect 437442 131960 437447 132016
rect 433934 131958 437447 131960
rect 131389 131955 131455 131958
rect 433934 131444 433994 131958
rect 437381 131955 437447 131958
rect 132125 130930 132191 130933
rect 132125 130928 134044 130930
rect 132125 130872 132130 130928
rect 132186 130872 134044 130928
rect 132125 130870 134044 130872
rect 132125 130867 132191 130870
rect 133229 129842 133295 129845
rect 133229 129840 134044 129842
rect 133229 129784 133234 129840
rect 133290 129784 134044 129840
rect 133229 129782 134044 129784
rect 133229 129779 133295 129782
rect 437381 129570 437447 129573
rect 433934 129568 437447 129570
rect 433934 129512 437386 129568
rect 437442 129512 437447 129568
rect 433934 129510 437447 129512
rect 433934 129268 433994 129510
rect 437381 129507 437447 129510
rect 131941 128754 132007 128757
rect 131941 128752 134044 128754
rect 131941 128696 131946 128752
rect 132002 128696 134044 128752
rect 131941 128694 134044 128696
rect 131941 128691 132007 128694
rect 132033 127802 132099 127805
rect 436829 127802 436895 127805
rect 132033 127800 134044 127802
rect 132033 127744 132038 127800
rect 132094 127744 134044 127800
rect 132033 127742 134044 127744
rect 433934 127800 436895 127802
rect 433934 127744 436834 127800
rect 436890 127744 436895 127800
rect 433934 127742 436895 127744
rect 132033 127739 132099 127742
rect 433934 127228 433994 127742
rect 436829 127739 436895 127742
rect 131849 126714 131915 126717
rect 131849 126712 134044 126714
rect 131849 126656 131854 126712
rect 131910 126656 134044 126712
rect 131849 126654 134044 126656
rect 131849 126651 131915 126654
rect 131573 125626 131639 125629
rect 131573 125624 134044 125626
rect 131573 125568 131578 125624
rect 131634 125568 134044 125624
rect 131573 125566 134044 125568
rect 131573 125563 131639 125566
rect 131481 124538 131547 124541
rect 433934 124538 433994 125052
rect 436921 124538 436987 124541
rect 131481 124536 134044 124538
rect 131481 124480 131486 124536
rect 131542 124480 134044 124536
rect 131481 124478 134044 124480
rect 433934 124536 436987 124538
rect 433934 124480 436926 124536
rect 436982 124480 436987 124536
rect 433934 124478 436987 124480
rect 131481 124475 131547 124478
rect 436921 124475 436987 124478
rect 131113 124266 131179 124269
rect 131297 124266 131363 124269
rect 131113 124264 131363 124266
rect 131113 124208 131118 124264
rect 131174 124208 131302 124264
rect 131358 124208 131363 124264
rect 131113 124206 131363 124208
rect 131113 124203 131179 124206
rect 131297 124203 131363 124206
rect 134014 123045 134074 123556
rect 580901 123178 580967 123181
rect 583520 123178 584960 123268
rect 580901 123176 584960 123178
rect 580901 123120 580906 123176
rect 580962 123120 584960 123176
rect 580901 123118 584960 123120
rect 580901 123115 580967 123118
rect 133965 123040 134074 123045
rect 133965 122984 133970 123040
rect 134026 122984 134074 123040
rect 583520 123028 584960 123118
rect 133965 122982 134074 122984
rect 133965 122979 134031 122982
rect 433934 122906 433994 123012
rect 436829 122906 436895 122909
rect 433934 122904 436895 122906
rect 433934 122848 436834 122904
rect 436890 122848 436895 122904
rect 433934 122846 436895 122848
rect 436829 122843 436895 122846
rect -960 122090 480 122180
rect 3325 122090 3391 122093
rect -960 122088 3391 122090
rect -960 122032 3330 122088
rect 3386 122032 3391 122088
rect -960 122030 3391 122032
rect -960 121940 480 122030
rect 3325 122027 3391 122030
rect 134014 121957 134074 122468
rect 134014 121952 134123 121957
rect 134014 121896 134062 121952
rect 134118 121896 134123 121952
rect 134014 121894 134123 121896
rect 134057 121891 134123 121894
rect 132125 121410 132191 121413
rect 132125 121408 134044 121410
rect 132125 121352 132130 121408
rect 132186 121352 134044 121408
rect 132125 121350 134044 121352
rect 132125 121347 132191 121350
rect 132401 120458 132467 120461
rect 433934 120458 433994 120972
rect 436737 120458 436803 120461
rect 132401 120456 134044 120458
rect 132401 120400 132406 120456
rect 132462 120400 134044 120456
rect 132401 120398 134044 120400
rect 433934 120456 436803 120458
rect 433934 120400 436742 120456
rect 436798 120400 436803 120456
rect 433934 120398 436803 120400
rect 132401 120395 132467 120398
rect 436737 120395 436803 120398
rect 133822 119716 133828 119780
rect 133892 119778 133898 119780
rect 138519 119778 138585 119781
rect 133892 119776 138585 119778
rect 133892 119720 138524 119776
rect 138580 119720 138585 119776
rect 133892 119718 138585 119720
rect 133892 119716 133898 119718
rect 138519 119715 138585 119718
rect 99281 118690 99347 118693
rect 184933 118690 184999 118693
rect 99281 118688 184999 118690
rect 99281 118632 99286 118688
rect 99342 118632 184938 118688
rect 184994 118632 184999 118688
rect 99281 118630 184999 118632
rect 99281 118627 99347 118630
rect 184933 118627 184999 118630
rect 69657 118554 69723 118557
rect 153469 118554 153535 118557
rect 69657 118552 153535 118554
rect 69657 118496 69662 118552
rect 69718 118496 153474 118552
rect 153530 118496 153535 118552
rect 69657 118494 153535 118496
rect 69657 118491 69723 118494
rect 153469 118491 153535 118494
rect 110321 118418 110387 118421
rect 145557 118418 145623 118421
rect 110321 118416 145623 118418
rect 110321 118360 110326 118416
rect 110382 118360 145562 118416
rect 145618 118360 145623 118416
rect 110321 118358 145623 118360
rect 110321 118355 110387 118358
rect 145557 118355 145623 118358
rect 128261 118282 128327 118285
rect 193949 118282 194015 118285
rect 128261 118280 194015 118282
rect 128261 118224 128266 118280
rect 128322 118224 193954 118280
rect 194010 118224 194015 118280
rect 128261 118222 194015 118224
rect 128261 118219 128327 118222
rect 193949 118219 194015 118222
rect 132861 118146 132927 118149
rect 133321 118146 133387 118149
rect 188429 118146 188495 118149
rect 132861 118144 188495 118146
rect 132861 118088 132866 118144
rect 132922 118088 133326 118144
rect 133382 118088 188434 118144
rect 188490 118088 188495 118144
rect 132861 118086 188495 118088
rect 132861 118083 132927 118086
rect 133321 118083 133387 118086
rect 188429 118083 188495 118086
rect 133045 118010 133111 118013
rect 175273 118010 175339 118013
rect 133045 118008 175339 118010
rect 133045 117952 133050 118008
rect 133106 117952 175278 118008
rect 175334 117952 175339 118008
rect 133045 117950 175339 117952
rect 133045 117947 133111 117950
rect 175273 117947 175339 117950
rect 433977 118010 434043 118013
rect 442257 118010 442323 118013
rect 433977 118008 442323 118010
rect 433977 117952 433982 118008
rect 434038 117952 442262 118008
rect 442318 117952 442323 118008
rect 433977 117950 442323 117952
rect 433977 117947 434043 117950
rect 442257 117947 442323 117950
rect 71589 117874 71655 117877
rect 79961 117874 80027 117877
rect 71589 117872 80027 117874
rect 71589 117816 71594 117872
rect 71650 117816 79966 117872
rect 80022 117816 80027 117872
rect 71589 117814 80027 117816
rect 71589 117811 71655 117814
rect 79961 117811 80027 117814
rect 89805 117874 89871 117877
rect 99189 117874 99255 117877
rect 89805 117872 99255 117874
rect 89805 117816 89810 117872
rect 89866 117816 99194 117872
rect 99250 117816 99255 117872
rect 89805 117814 99255 117816
rect 89805 117811 89871 117814
rect 99189 117811 99255 117814
rect 101213 117874 101279 117877
rect 103513 117874 103579 117877
rect 115197 117874 115263 117877
rect 122833 117874 122899 117877
rect 133781 117876 133847 117877
rect 133781 117874 133828 117876
rect 101213 117872 104818 117874
rect 101213 117816 101218 117872
rect 101274 117816 103518 117872
rect 103574 117816 104818 117872
rect 101213 117814 104818 117816
rect 101213 117811 101279 117814
rect 103513 117811 103579 117814
rect 80145 117738 80211 117741
rect 89621 117738 89687 117741
rect 80145 117736 89687 117738
rect 80145 117680 80150 117736
rect 80206 117680 89626 117736
rect 89682 117680 89687 117736
rect 80145 117678 89687 117680
rect 104758 117738 104818 117814
rect 115197 117872 122899 117874
rect 115197 117816 115202 117872
rect 115258 117816 122838 117872
rect 122894 117816 122899 117872
rect 115197 117814 122899 117816
rect 133740 117872 133828 117874
rect 133740 117816 133786 117872
rect 133740 117814 133828 117816
rect 115197 117811 115263 117814
rect 122833 117811 122899 117814
rect 133781 117812 133828 117814
rect 133892 117812 133898 117876
rect 133781 117811 133847 117812
rect 104985 117738 105051 117741
rect 104758 117736 105051 117738
rect 104758 117680 104990 117736
rect 105046 117680 105051 117736
rect 104758 117678 105051 117680
rect 80145 117675 80211 117678
rect 89621 117675 89687 117678
rect 104985 117675 105051 117678
rect 129457 117738 129523 117741
rect 133965 117738 134031 117741
rect 129457 117736 134031 117738
rect 129457 117680 129462 117736
rect 129518 117680 133970 117736
rect 134026 117680 134031 117736
rect 129457 117678 134031 117680
rect 129457 117675 129523 117678
rect 133965 117675 134031 117678
rect 134149 117738 134215 117741
rect 151905 117738 151971 117741
rect 134149 117736 151971 117738
rect 134149 117680 134154 117736
rect 134210 117680 151910 117736
rect 151966 117680 151971 117736
rect 134149 117678 151971 117680
rect 134149 117675 134215 117678
rect 151905 117675 151971 117678
rect 418153 117738 418219 117741
rect 427721 117738 427787 117741
rect 418153 117736 427787 117738
rect 418153 117680 418158 117736
rect 418214 117680 427726 117736
rect 427782 117680 427787 117736
rect 418153 117678 427787 117680
rect 418153 117675 418219 117678
rect 427721 117675 427787 117678
rect 126053 117602 126119 117605
rect 133822 117602 133828 117604
rect 126053 117600 133828 117602
rect 126053 117544 126058 117600
rect 126114 117544 133828 117600
rect 126053 117542 133828 117544
rect 126053 117539 126119 117542
rect 133822 117540 133828 117542
rect 133892 117540 133898 117604
rect 197629 117602 197695 117605
rect 134060 117600 197695 117602
rect 134060 117544 197634 117600
rect 197690 117544 197695 117600
rect 134060 117542 197695 117544
rect 133822 117404 133828 117468
rect 133892 117466 133898 117468
rect 134060 117466 134120 117542
rect 197629 117539 197695 117542
rect 133892 117406 134120 117466
rect 133892 117404 133898 117406
rect 97993 117330 98059 117333
rect 99281 117330 99347 117333
rect 97993 117328 99347 117330
rect 97993 117272 97998 117328
rect 98054 117272 99286 117328
rect 99342 117272 99347 117328
rect 97993 117270 99347 117272
rect 97993 117267 98059 117270
rect 99281 117267 99347 117270
rect 127617 117330 127683 117333
rect 128261 117330 128327 117333
rect 127617 117328 128327 117330
rect 127617 117272 127622 117328
rect 127678 117272 128266 117328
rect 128322 117272 128327 117328
rect 127617 117270 128327 117272
rect 127617 117267 127683 117270
rect 128261 117267 128327 117270
rect 243629 117330 243695 117333
rect 245745 117330 245811 117333
rect 243629 117328 245811 117330
rect 243629 117272 243634 117328
rect 243690 117272 245750 117328
rect 245806 117272 245811 117328
rect 243629 117270 245811 117272
rect 243629 117267 243695 117270
rect 245745 117267 245811 117270
rect 301405 116106 301471 116109
rect 388345 116106 388411 116109
rect 301405 116104 301882 116106
rect 301405 116048 301410 116104
rect 301466 116048 301882 116104
rect 301405 116046 301882 116048
rect 301405 116043 301471 116046
rect 301822 115973 301882 116046
rect 388345 116104 388914 116106
rect 388345 116048 388350 116104
rect 388406 116048 388914 116104
rect 388345 116046 388914 116048
rect 388345 116043 388411 116046
rect 157517 115970 157583 115973
rect 157885 115970 157951 115973
rect 157517 115968 157951 115970
rect 157517 115912 157522 115968
rect 157578 115912 157890 115968
rect 157946 115912 157951 115968
rect 157517 115910 157951 115912
rect 157517 115907 157583 115910
rect 157885 115907 157951 115910
rect 161749 115970 161815 115973
rect 162117 115970 162183 115973
rect 161749 115968 162183 115970
rect 161749 115912 161754 115968
rect 161810 115912 162122 115968
rect 162178 115912 162183 115968
rect 161749 115910 162183 115912
rect 161749 115907 161815 115910
rect 162117 115907 162183 115910
rect 183829 115970 183895 115973
rect 184105 115970 184171 115973
rect 183829 115968 184171 115970
rect 183829 115912 183834 115968
rect 183890 115912 184110 115968
rect 184166 115912 184171 115968
rect 183829 115910 184171 115912
rect 183829 115907 183895 115910
rect 184105 115907 184171 115910
rect 216949 115970 217015 115973
rect 217317 115970 217383 115973
rect 216949 115968 217383 115970
rect 216949 115912 216954 115968
rect 217010 115912 217322 115968
rect 217378 115912 217383 115968
rect 216949 115910 217383 115912
rect 216949 115907 217015 115910
rect 217317 115907 217383 115910
rect 220997 115970 221063 115973
rect 221457 115970 221523 115973
rect 220997 115968 221523 115970
rect 220997 115912 221002 115968
rect 221058 115912 221462 115968
rect 221518 115912 221523 115968
rect 220997 115910 221523 115912
rect 220997 115907 221063 115910
rect 221457 115907 221523 115910
rect 301773 115968 301882 115973
rect 301773 115912 301778 115968
rect 301834 115912 301882 115968
rect 301773 115910 301882 115912
rect 388713 115970 388779 115973
rect 388854 115970 388914 116046
rect 388713 115968 388914 115970
rect 388713 115912 388718 115968
rect 388774 115912 388914 115968
rect 388713 115910 388914 115912
rect 301773 115907 301839 115910
rect 388713 115907 388779 115910
rect 579797 111482 579863 111485
rect 583520 111482 584960 111572
rect 579797 111480 584960 111482
rect 579797 111424 579802 111480
rect 579858 111424 584960 111480
rect 579797 111422 584960 111424
rect 579797 111419 579863 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3509 107674 3575 107677
rect -960 107672 3575 107674
rect -960 107616 3514 107672
rect 3570 107616 3575 107672
rect -960 107614 3575 107616
rect -960 107524 480 107614
rect 3509 107611 3575 107614
rect 276013 106450 276079 106453
rect 276013 106448 276122 106450
rect 276013 106392 276018 106448
rect 276074 106392 276122 106448
rect 276013 106387 276122 106392
rect 276062 106317 276122 106387
rect 133781 106314 133847 106317
rect 133965 106314 134031 106317
rect 133781 106312 134031 106314
rect 133781 106256 133786 106312
rect 133842 106256 133970 106312
rect 134026 106256 134031 106312
rect 133781 106254 134031 106256
rect 133781 106251 133847 106254
rect 133965 106251 134031 106254
rect 275001 106314 275067 106317
rect 275369 106314 275435 106317
rect 275001 106312 275435 106314
rect 275001 106256 275006 106312
rect 275062 106256 275374 106312
rect 275430 106256 275435 106312
rect 275001 106254 275435 106256
rect 276062 106312 276171 106317
rect 276062 106256 276110 106312
rect 276166 106256 276171 106312
rect 276062 106254 276171 106256
rect 275001 106251 275067 106254
rect 275369 106251 275435 106254
rect 276105 106251 276171 106254
rect 388713 106314 388779 106317
rect 388897 106314 388963 106317
rect 388713 106312 388963 106314
rect 388713 106256 388718 106312
rect 388774 106256 388902 106312
rect 388958 106256 388963 106312
rect 388713 106254 388963 106256
rect 388713 106251 388779 106254
rect 388897 106251 388963 106254
rect 583520 99636 584960 99876
rect 290641 99516 290707 99517
rect 341425 99516 341491 99517
rect 290590 99514 290596 99516
rect 290550 99454 290596 99514
rect 290660 99512 290707 99516
rect 341374 99514 341380 99516
rect 290702 99456 290707 99512
rect 290590 99452 290596 99454
rect 290660 99452 290707 99456
rect 341334 99454 341380 99514
rect 341444 99512 341491 99516
rect 341486 99456 341491 99512
rect 341374 99452 341380 99454
rect 341444 99452 341491 99456
rect 290641 99451 290707 99452
rect 341425 99451 341491 99452
rect 190913 96794 190979 96797
rect 190502 96792 190979 96794
rect 190502 96736 190918 96792
rect 190974 96736 190979 96792
rect 190502 96734 190979 96736
rect 131205 96658 131271 96661
rect 131389 96658 131455 96661
rect 131205 96656 131455 96658
rect 131205 96600 131210 96656
rect 131266 96600 131394 96656
rect 131450 96600 131455 96656
rect 131205 96598 131455 96600
rect 190502 96658 190562 96734
rect 190913 96731 190979 96734
rect 190637 96658 190703 96661
rect 190502 96656 190703 96658
rect 190502 96600 190642 96656
rect 190698 96600 190703 96656
rect 190502 96598 190703 96600
rect 131205 96595 131271 96598
rect 131389 96595 131455 96598
rect 190637 96595 190703 96598
rect 248413 96658 248479 96661
rect 248597 96658 248663 96661
rect 248413 96656 248663 96658
rect 248413 96600 248418 96656
rect 248474 96600 248602 96656
rect 248658 96600 248663 96656
rect 248413 96598 248663 96600
rect 248413 96595 248479 96598
rect 248597 96595 248663 96598
rect 274725 96658 274791 96661
rect 275001 96658 275067 96661
rect 274725 96656 275067 96658
rect 274725 96600 274730 96656
rect 274786 96600 275006 96656
rect 275062 96600 275067 96656
rect 274725 96598 275067 96600
rect 274725 96595 274791 96598
rect 275001 96595 275067 96598
rect 290549 96660 290615 96661
rect 341333 96660 341399 96661
rect 290549 96656 290596 96660
rect 290660 96658 290666 96660
rect 290549 96600 290554 96656
rect 290549 96596 290596 96600
rect 290660 96598 290706 96658
rect 341333 96656 341380 96660
rect 341444 96658 341450 96660
rect 341333 96600 341338 96656
rect 290660 96596 290666 96598
rect 341333 96596 341380 96600
rect 341444 96598 341490 96658
rect 341444 96596 341450 96598
rect 290549 96595 290615 96596
rect 341333 96595 341399 96596
rect -960 93258 480 93348
rect 2773 93258 2839 93261
rect -960 93256 2839 93258
rect -960 93200 2778 93256
rect 2834 93200 2839 93256
rect -960 93198 2839 93200
rect -960 93108 480 93198
rect 2773 93195 2839 93198
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect 214097 87002 214163 87005
rect 214281 87002 214347 87005
rect 214097 87000 214347 87002
rect 214097 86944 214102 87000
rect 214158 86944 214286 87000
rect 214342 86944 214347 87000
rect 214097 86942 214347 86944
rect 214097 86939 214163 86942
rect 214281 86939 214347 86942
rect 341057 87002 341123 87005
rect 341241 87002 341307 87005
rect 341057 87000 341307 87002
rect 341057 86944 341062 87000
rect 341118 86944 341246 87000
rect 341302 86944 341307 87000
rect 341057 86942 341307 86944
rect 341057 86939 341123 86942
rect 341241 86939 341307 86942
rect -960 78978 480 79068
rect 3233 78978 3299 78981
rect -960 78976 3299 78978
rect -960 78920 3238 78976
rect 3294 78920 3299 78976
rect -960 78918 3299 78920
rect -960 78828 480 78918
rect 3233 78915 3299 78918
rect 420269 77346 420335 77349
rect 420453 77346 420519 77349
rect 420269 77344 420519 77346
rect 420269 77288 420274 77344
rect 420330 77288 420458 77344
rect 420514 77288 420519 77344
rect 420269 77286 420519 77288
rect 420269 77283 420335 77286
rect 420453 77283 420519 77286
rect 580165 76258 580231 76261
rect 583520 76258 584960 76348
rect 580165 76256 584960 76258
rect 580165 76200 580170 76256
rect 580226 76200 584960 76256
rect 580165 76198 584960 76200
rect 580165 76195 580231 76198
rect 583520 76108 584960 76198
rect 157333 70412 157399 70413
rect 157333 70408 157380 70412
rect 157444 70410 157450 70412
rect 157333 70352 157338 70408
rect 157333 70348 157380 70352
rect 157444 70350 157490 70410
rect 157444 70348 157450 70350
rect 157333 70347 157399 70348
rect 128629 67690 128695 67693
rect 128813 67690 128879 67693
rect 128629 67688 128879 67690
rect 128629 67632 128634 67688
rect 128690 67632 128818 67688
rect 128874 67632 128879 67688
rect 128629 67630 128879 67632
rect 128629 67627 128695 67630
rect 128813 67627 128879 67630
rect 290406 67628 290412 67692
rect 290476 67690 290482 67692
rect 290549 67690 290615 67693
rect 290476 67688 290615 67690
rect 290476 67632 290554 67688
rect 290610 67632 290615 67688
rect 290476 67630 290615 67632
rect 290476 67628 290482 67630
rect 290549 67627 290615 67630
rect 157333 66332 157399 66333
rect 290457 66332 290523 66333
rect 157333 66328 157380 66332
rect 157444 66330 157450 66332
rect 157333 66272 157338 66328
rect 157333 66268 157380 66272
rect 157444 66270 157490 66330
rect 157444 66268 157450 66270
rect 290406 66268 290412 66332
rect 290476 66330 290523 66332
rect 290476 66328 290568 66330
rect 290518 66272 290568 66328
rect 290476 66270 290568 66272
rect 290476 66268 290523 66270
rect 157333 66267 157399 66268
rect 290457 66267 290523 66268
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 420637 61436 420703 61437
rect 420637 61434 420684 61436
rect 420592 61432 420684 61434
rect 420592 61376 420642 61432
rect 420592 61374 420684 61376
rect 420637 61372 420684 61374
rect 420748 61372 420754 61436
rect 420637 61371 420703 61372
rect 220721 53954 220787 53957
rect 220997 53954 221063 53957
rect 220721 53952 221063 53954
rect 220721 53896 220726 53952
rect 220782 53896 221002 53952
rect 221058 53896 221063 53952
rect 220721 53894 221063 53896
rect 220721 53891 220787 53894
rect 220997 53891 221063 53894
rect 220997 53818 221063 53821
rect 221181 53818 221247 53821
rect 220997 53816 221247 53818
rect 220997 53760 221002 53816
rect 221058 53760 221186 53816
rect 221242 53760 221247 53816
rect 220997 53758 221247 53760
rect 220997 53755 221063 53758
rect 221181 53755 221247 53758
rect 583520 52716 584960 52956
rect -960 50146 480 50236
rect 3417 50146 3483 50149
rect -960 50144 3483 50146
rect -960 50088 3422 50144
rect 3478 50088 3483 50144
rect -960 50086 3483 50088
rect -960 49996 480 50086
rect 3417 50083 3483 50086
rect 276105 48378 276171 48381
rect 276289 48378 276355 48381
rect 276105 48376 276355 48378
rect 276105 48320 276110 48376
rect 276166 48320 276294 48376
rect 276350 48320 276355 48376
rect 276105 48318 276355 48320
rect 276105 48315 276171 48318
rect 276289 48315 276355 48318
rect 325509 48378 325575 48381
rect 325693 48378 325759 48381
rect 325509 48376 325759 48378
rect 325509 48320 325514 48376
rect 325570 48320 325698 48376
rect 325754 48320 325759 48376
rect 325509 48318 325759 48320
rect 325509 48315 325575 48318
rect 325693 48315 325759 48318
rect 415025 48378 415091 48381
rect 415209 48378 415275 48381
rect 415025 48376 415275 48378
rect 415025 48320 415030 48376
rect 415086 48320 415214 48376
rect 415270 48320 415275 48376
rect 415025 48318 415275 48320
rect 415025 48315 415091 48318
rect 415209 48315 415275 48318
rect 420545 48378 420611 48381
rect 420678 48378 420684 48380
rect 420545 48376 420684 48378
rect 420545 48320 420550 48376
rect 420606 48320 420684 48376
rect 420545 48318 420684 48320
rect 420545 48315 420611 48318
rect 420678 48316 420684 48318
rect 420748 48316 420754 48380
rect 426065 48378 426131 48381
rect 426249 48378 426315 48381
rect 426065 48376 426315 48378
rect 426065 48320 426070 48376
rect 426126 48320 426254 48376
rect 426310 48320 426315 48376
rect 426065 48318 426315 48320
rect 426065 48315 426131 48318
rect 426249 48315 426315 48318
rect 431585 47018 431651 47021
rect 431769 47018 431835 47021
rect 431585 47016 431835 47018
rect 431585 46960 431590 47016
rect 431646 46960 431774 47016
rect 431830 46960 431835 47016
rect 431585 46958 431835 46960
rect 431585 46955 431651 46958
rect 431769 46955 431835 46958
rect 420637 42124 420703 42125
rect 420637 42122 420684 42124
rect 420592 42120 420684 42122
rect 420592 42064 420642 42120
rect 420592 42062 420684 42064
rect 420637 42060 420684 42062
rect 420748 42060 420754 42124
rect 420637 42059 420703 42060
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect 140865 38588 140931 38589
rect 140814 38524 140820 38588
rect 140884 38586 140931 38588
rect 140884 38584 140976 38586
rect 140926 38528 140976 38584
rect 140884 38526 140976 38528
rect 140884 38524 140931 38526
rect 140865 38523 140931 38524
rect 179689 37498 179755 37501
rect 179278 37496 179755 37498
rect 179278 37440 179694 37496
rect 179750 37440 179755 37496
rect 179278 37438 179755 37440
rect 179278 37362 179338 37438
rect 179689 37435 179755 37438
rect 179413 37362 179479 37365
rect 179278 37360 179479 37362
rect 179278 37304 179418 37360
rect 179474 37304 179479 37360
rect 179278 37302 179479 37304
rect 179413 37299 179479 37302
rect -960 35866 480 35956
rect 3417 35866 3483 35869
rect 230381 35866 230447 35869
rect -960 35864 3483 35866
rect -960 35808 3422 35864
rect 3478 35808 3483 35864
rect -960 35806 3483 35808
rect -960 35716 480 35806
rect 3417 35803 3483 35806
rect 230246 35864 230447 35866
rect 230246 35808 230386 35864
rect 230442 35808 230447 35864
rect 230246 35806 230447 35808
rect 230246 35730 230306 35806
rect 230381 35803 230447 35806
rect 230657 35730 230723 35733
rect 230246 35728 230723 35730
rect 230246 35672 230662 35728
rect 230718 35672 230723 35728
rect 230246 35670 230723 35672
rect 230657 35667 230723 35670
rect 227897 34642 227963 34645
rect 228173 34642 228239 34645
rect 227897 34640 228239 34642
rect 227897 34584 227902 34640
rect 227958 34584 228178 34640
rect 228234 34584 228239 34640
rect 227897 34582 228239 34584
rect 227897 34579 227963 34582
rect 228173 34579 228239 34582
rect 220997 34506 221063 34509
rect 221181 34506 221247 34509
rect 220997 34504 221247 34506
rect 220997 34448 221002 34504
rect 221058 34448 221186 34504
rect 221242 34448 221247 34504
rect 220997 34446 221247 34448
rect 220997 34443 221063 34446
rect 221181 34443 221247 34446
rect 580165 29338 580231 29341
rect 583520 29338 584960 29428
rect 580165 29336 584960 29338
rect 580165 29280 580170 29336
rect 580226 29280 584960 29336
rect 580165 29278 584960 29280
rect 580165 29275 580231 29278
rect 583520 29188 584960 29278
rect 140814 29004 140820 29068
rect 140884 29066 140890 29068
rect 140957 29066 141023 29069
rect 140884 29064 141023 29066
rect 140884 29008 140962 29064
rect 141018 29008 141023 29064
rect 140884 29006 141023 29008
rect 140884 29004 140890 29006
rect 140957 29003 141023 29006
rect 420545 29066 420611 29069
rect 420678 29066 420684 29068
rect 420545 29064 420684 29066
rect 420545 29008 420550 29064
rect 420606 29008 420684 29064
rect 420545 29006 420684 29008
rect 420545 29003 420611 29006
rect 420678 29004 420684 29006
rect 420748 29004 420754 29068
rect 230473 26346 230539 26349
rect 230657 26346 230723 26349
rect 230473 26344 230723 26346
rect 230473 26288 230478 26344
rect 230534 26288 230662 26344
rect 230718 26288 230723 26344
rect 230473 26286 230723 26288
rect 230473 26283 230539 26286
rect 230657 26283 230723 26286
rect 301865 26346 301931 26349
rect 302049 26346 302115 26349
rect 301865 26344 302115 26346
rect 301865 26288 301870 26344
rect 301926 26288 302054 26344
rect 302110 26288 302115 26344
rect 301865 26286 302115 26288
rect 301865 26283 301931 26286
rect 302049 26283 302115 26286
rect -960 21450 480 21540
rect 3141 21450 3207 21453
rect -960 21448 3207 21450
rect -960 21392 3146 21448
rect 3202 21392 3207 21448
rect -960 21390 3207 21392
rect -960 21300 480 21390
rect 3141 21387 3207 21390
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 102777 6218 102843 6221
rect 186405 6218 186471 6221
rect 102777 6216 186471 6218
rect 102777 6160 102782 6216
rect 102838 6160 186410 6216
rect 186466 6160 186471 6216
rect 102777 6158 186471 6160
rect 102777 6155 102843 6158
rect 186405 6155 186471 6158
rect 411069 6218 411135 6221
rect 538121 6218 538187 6221
rect 411069 6216 538187 6218
rect 411069 6160 411074 6216
rect 411130 6160 538126 6216
rect 538182 6160 538187 6216
rect 411069 6158 538187 6160
rect 411069 6155 411135 6158
rect 538121 6155 538187 6158
rect 583520 5796 584960 6036
rect 30281 4858 30347 4861
rect 149053 4858 149119 4861
rect 30281 4856 149119 4858
rect 30281 4800 30286 4856
rect 30342 4800 149058 4856
rect 149114 4800 149119 4856
rect 30281 4798 149119 4800
rect 30281 4795 30347 4798
rect 149053 4795 149119 4798
rect 357341 4858 357407 4861
rect 433517 4858 433583 4861
rect 357341 4856 433583 4858
rect 357341 4800 357346 4856
rect 357402 4800 433522 4856
rect 433578 4800 433583 4856
rect 357341 4798 433583 4800
rect 357341 4795 357407 4798
rect 433517 4795 433583 4798
rect 408309 3770 408375 3773
rect 408493 3770 408559 3773
rect 408309 3768 408559 3770
rect 408309 3712 408314 3768
rect 408370 3712 408498 3768
rect 408554 3712 408559 3768
rect 408309 3710 408559 3712
rect 408309 3707 408375 3710
rect 408493 3707 408559 3710
rect 417877 3634 417943 3637
rect 418337 3634 418403 3637
rect 417877 3632 418403 3634
rect 417877 3576 417882 3632
rect 417938 3576 418342 3632
rect 418398 3576 418403 3632
rect 417877 3574 418403 3576
rect 417877 3571 417943 3574
rect 418337 3571 418403 3574
rect 427629 3634 427695 3637
rect 427813 3634 427879 3637
rect 427629 3632 427879 3634
rect 427629 3576 427634 3632
rect 427690 3576 427818 3632
rect 427874 3576 427879 3632
rect 427629 3574 427879 3576
rect 427629 3571 427695 3574
rect 427813 3571 427879 3574
rect 431217 3362 431283 3365
rect 575013 3362 575079 3365
rect 431217 3360 575079 3362
rect 431217 3304 431222 3360
rect 431278 3304 575018 3360
rect 575074 3304 575079 3360
rect 431217 3302 575079 3304
rect 431217 3299 431283 3302
rect 575013 3299 575079 3302
<< via3 >>
rect 132172 700436 132236 700500
rect 132356 700300 132420 700364
rect 133644 697172 133708 697236
rect 164188 686428 164252 686492
rect 131988 685884 132052 685948
rect 164188 686156 164252 686220
rect 164188 650524 164252 650588
rect 133460 650252 133524 650316
rect 164188 650252 164252 650316
rect 131804 638964 131868 639028
rect 164188 639100 164252 639164
rect 164188 638828 164252 638892
rect 133092 603332 133156 603396
rect 164188 603196 164252 603260
rect 164188 602924 164252 602988
rect 133276 592316 133340 592380
rect 164188 592180 164252 592244
rect 164188 591908 164252 591972
rect 379468 572052 379532 572116
rect 199700 561716 199764 561780
rect 198596 556684 198660 556748
rect 198412 552060 198476 552124
rect 198228 547844 198292 547908
rect 198044 543764 198108 543828
rect 379652 541044 379716 541108
rect 197860 538460 197924 538524
rect 379468 500244 379532 500308
rect 379652 500108 379716 500172
rect 266860 410348 266924 410412
rect 267964 410212 268028 410276
rect 267780 410076 267844 410140
rect 268148 409940 268212 410004
rect 268148 338676 268212 338740
rect 257660 317384 257724 317388
rect 257660 317328 257710 317384
rect 257710 317328 257724 317384
rect 257660 317324 257724 317328
rect 257660 311748 257724 311812
rect 128860 299236 128924 299300
rect 128860 289912 128924 289916
rect 128860 289856 128874 289912
rect 128874 289856 128924 289912
rect 128860 289852 128924 289856
rect 197860 202540 197924 202604
rect 198228 202268 198292 202332
rect 267964 202132 268028 202196
rect 199700 201996 199764 202060
rect 198412 201860 198476 201924
rect 198596 201724 198660 201788
rect 198044 201588 198108 201652
rect 267780 201588 267844 201652
rect 266860 201452 266924 201516
rect 132908 200636 132972 200700
rect 132908 176156 132972 176220
rect 133644 175068 133708 175132
rect 133460 173980 133524 174044
rect 133092 172892 133156 172956
rect 132172 137124 132236 137188
rect 132356 136172 132420 136236
rect 131988 135084 132052 135148
rect 131804 133996 131868 134060
rect 133276 132908 133340 132972
rect 133828 119716 133892 119780
rect 133828 117872 133892 117876
rect 133828 117816 133842 117872
rect 133842 117816 133892 117872
rect 133828 117812 133892 117816
rect 133828 117540 133892 117604
rect 133828 117404 133892 117468
rect 290596 99512 290660 99516
rect 290596 99456 290646 99512
rect 290646 99456 290660 99512
rect 290596 99452 290660 99456
rect 341380 99512 341444 99516
rect 341380 99456 341430 99512
rect 341430 99456 341444 99512
rect 341380 99452 341444 99456
rect 290596 96656 290660 96660
rect 290596 96600 290610 96656
rect 290610 96600 290660 96656
rect 290596 96596 290660 96600
rect 341380 96656 341444 96660
rect 341380 96600 341394 96656
rect 341394 96600 341444 96656
rect 341380 96596 341444 96600
rect 157380 70408 157444 70412
rect 157380 70352 157394 70408
rect 157394 70352 157444 70408
rect 157380 70348 157444 70352
rect 290412 67628 290476 67692
rect 157380 66328 157444 66332
rect 157380 66272 157394 66328
rect 157394 66272 157444 66328
rect 157380 66268 157444 66272
rect 290412 66328 290476 66332
rect 290412 66272 290462 66328
rect 290462 66272 290476 66328
rect 290412 66268 290476 66272
rect 420684 61432 420748 61436
rect 420684 61376 420698 61432
rect 420698 61376 420748 61432
rect 420684 61372 420748 61376
rect 420684 48316 420748 48380
rect 420684 42120 420748 42124
rect 420684 42064 420698 42120
rect 420698 42064 420748 42120
rect 420684 42060 420748 42064
rect 140820 38584 140884 38588
rect 140820 38528 140870 38584
rect 140870 38528 140884 38584
rect 140820 38524 140884 38528
rect 140820 29004 140884 29068
rect 420684 29004 420748 29068
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 679254 -7976 710862
rect -8576 679018 -8394 679254
rect -8158 679018 -7976 679254
rect -8576 678934 -7976 679018
rect -8576 678698 -8394 678934
rect -8158 678698 -7976 678934
rect -8576 643254 -7976 678698
rect -8576 643018 -8394 643254
rect -8158 643018 -7976 643254
rect -8576 642934 -7976 643018
rect -8576 642698 -8394 642934
rect -8158 642698 -7976 642934
rect -8576 607254 -7976 642698
rect -8576 607018 -8394 607254
rect -8158 607018 -7976 607254
rect -8576 606934 -7976 607018
rect -8576 606698 -8394 606934
rect -8158 606698 -7976 606934
rect -8576 571254 -7976 606698
rect -8576 571018 -8394 571254
rect -8158 571018 -7976 571254
rect -8576 570934 -7976 571018
rect -8576 570698 -8394 570934
rect -8158 570698 -7976 570934
rect -8576 535254 -7976 570698
rect -8576 535018 -8394 535254
rect -8158 535018 -7976 535254
rect -8576 534934 -7976 535018
rect -8576 534698 -8394 534934
rect -8158 534698 -7976 534934
rect -8576 499254 -7976 534698
rect -8576 499018 -8394 499254
rect -8158 499018 -7976 499254
rect -8576 498934 -7976 499018
rect -8576 498698 -8394 498934
rect -8158 498698 -7976 498934
rect -8576 463254 -7976 498698
rect -8576 463018 -8394 463254
rect -8158 463018 -7976 463254
rect -8576 462934 -7976 463018
rect -8576 462698 -8394 462934
rect -8158 462698 -7976 462934
rect -8576 427254 -7976 462698
rect -8576 427018 -8394 427254
rect -8158 427018 -7976 427254
rect -8576 426934 -7976 427018
rect -8576 426698 -8394 426934
rect -8158 426698 -7976 426934
rect -8576 391254 -7976 426698
rect -8576 391018 -8394 391254
rect -8158 391018 -7976 391254
rect -8576 390934 -7976 391018
rect -8576 390698 -8394 390934
rect -8158 390698 -7976 390934
rect -8576 355254 -7976 390698
rect -8576 355018 -8394 355254
rect -8158 355018 -7976 355254
rect -8576 354934 -7976 355018
rect -8576 354698 -8394 354934
rect -8158 354698 -7976 354934
rect -8576 319254 -7976 354698
rect -8576 319018 -8394 319254
rect -8158 319018 -7976 319254
rect -8576 318934 -7976 319018
rect -8576 318698 -8394 318934
rect -8158 318698 -7976 318934
rect -8576 283254 -7976 318698
rect -8576 283018 -8394 283254
rect -8158 283018 -7976 283254
rect -8576 282934 -7976 283018
rect -8576 282698 -8394 282934
rect -8158 282698 -7976 282934
rect -8576 247254 -7976 282698
rect -8576 247018 -8394 247254
rect -8158 247018 -7976 247254
rect -8576 246934 -7976 247018
rect -8576 246698 -8394 246934
rect -8158 246698 -7976 246934
rect -8576 211254 -7976 246698
rect -8576 211018 -8394 211254
rect -8158 211018 -7976 211254
rect -8576 210934 -7976 211018
rect -8576 210698 -8394 210934
rect -8158 210698 -7976 210934
rect -8576 175254 -7976 210698
rect -8576 175018 -8394 175254
rect -8158 175018 -7976 175254
rect -8576 174934 -7976 175018
rect -8576 174698 -8394 174934
rect -8158 174698 -7976 174934
rect -8576 139254 -7976 174698
rect -8576 139018 -8394 139254
rect -8158 139018 -7976 139254
rect -8576 138934 -7976 139018
rect -8576 138698 -8394 138934
rect -8158 138698 -7976 138934
rect -8576 103254 -7976 138698
rect -8576 103018 -8394 103254
rect -8158 103018 -7976 103254
rect -8576 102934 -7976 103018
rect -8576 102698 -8394 102934
rect -8158 102698 -7976 102934
rect -8576 67254 -7976 102698
rect -8576 67018 -8394 67254
rect -8158 67018 -7976 67254
rect -8576 66934 -7976 67018
rect -8576 66698 -8394 66934
rect -8158 66698 -7976 66934
rect -8576 31254 -7976 66698
rect -8576 31018 -8394 31254
rect -8158 31018 -7976 31254
rect -8576 30934 -7976 31018
rect -8576 30698 -8394 30934
rect -8158 30698 -7976 30934
rect -8576 -6926 -7976 30698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 697254 -7036 709922
rect 11604 710478 12204 711440
rect 11604 710242 11786 710478
rect 12022 710242 12204 710478
rect 11604 710158 12204 710242
rect 11604 709922 11786 710158
rect 12022 709922 12204 710158
rect -7636 697018 -7454 697254
rect -7218 697018 -7036 697254
rect -7636 696934 -7036 697018
rect -7636 696698 -7454 696934
rect -7218 696698 -7036 696934
rect -7636 661254 -7036 696698
rect -7636 661018 -7454 661254
rect -7218 661018 -7036 661254
rect -7636 660934 -7036 661018
rect -7636 660698 -7454 660934
rect -7218 660698 -7036 660934
rect -7636 625254 -7036 660698
rect -7636 625018 -7454 625254
rect -7218 625018 -7036 625254
rect -7636 624934 -7036 625018
rect -7636 624698 -7454 624934
rect -7218 624698 -7036 624934
rect -7636 589254 -7036 624698
rect -7636 589018 -7454 589254
rect -7218 589018 -7036 589254
rect -7636 588934 -7036 589018
rect -7636 588698 -7454 588934
rect -7218 588698 -7036 588934
rect -7636 553254 -7036 588698
rect -7636 553018 -7454 553254
rect -7218 553018 -7036 553254
rect -7636 552934 -7036 553018
rect -7636 552698 -7454 552934
rect -7218 552698 -7036 552934
rect -7636 517254 -7036 552698
rect -7636 517018 -7454 517254
rect -7218 517018 -7036 517254
rect -7636 516934 -7036 517018
rect -7636 516698 -7454 516934
rect -7218 516698 -7036 516934
rect -7636 481254 -7036 516698
rect -7636 481018 -7454 481254
rect -7218 481018 -7036 481254
rect -7636 480934 -7036 481018
rect -7636 480698 -7454 480934
rect -7218 480698 -7036 480934
rect -7636 445254 -7036 480698
rect -7636 445018 -7454 445254
rect -7218 445018 -7036 445254
rect -7636 444934 -7036 445018
rect -7636 444698 -7454 444934
rect -7218 444698 -7036 444934
rect -7636 409254 -7036 444698
rect -7636 409018 -7454 409254
rect -7218 409018 -7036 409254
rect -7636 408934 -7036 409018
rect -7636 408698 -7454 408934
rect -7218 408698 -7036 408934
rect -7636 373254 -7036 408698
rect -7636 373018 -7454 373254
rect -7218 373018 -7036 373254
rect -7636 372934 -7036 373018
rect -7636 372698 -7454 372934
rect -7218 372698 -7036 372934
rect -7636 337254 -7036 372698
rect -7636 337018 -7454 337254
rect -7218 337018 -7036 337254
rect -7636 336934 -7036 337018
rect -7636 336698 -7454 336934
rect -7218 336698 -7036 336934
rect -7636 301254 -7036 336698
rect -7636 301018 -7454 301254
rect -7218 301018 -7036 301254
rect -7636 300934 -7036 301018
rect -7636 300698 -7454 300934
rect -7218 300698 -7036 300934
rect -7636 265254 -7036 300698
rect -7636 265018 -7454 265254
rect -7218 265018 -7036 265254
rect -7636 264934 -7036 265018
rect -7636 264698 -7454 264934
rect -7218 264698 -7036 264934
rect -7636 229254 -7036 264698
rect -7636 229018 -7454 229254
rect -7218 229018 -7036 229254
rect -7636 228934 -7036 229018
rect -7636 228698 -7454 228934
rect -7218 228698 -7036 228934
rect -7636 193254 -7036 228698
rect -7636 193018 -7454 193254
rect -7218 193018 -7036 193254
rect -7636 192934 -7036 193018
rect -7636 192698 -7454 192934
rect -7218 192698 -7036 192934
rect -7636 157254 -7036 192698
rect -7636 157018 -7454 157254
rect -7218 157018 -7036 157254
rect -7636 156934 -7036 157018
rect -7636 156698 -7454 156934
rect -7218 156698 -7036 156934
rect -7636 121254 -7036 156698
rect -7636 121018 -7454 121254
rect -7218 121018 -7036 121254
rect -7636 120934 -7036 121018
rect -7636 120698 -7454 120934
rect -7218 120698 -7036 120934
rect -7636 85254 -7036 120698
rect -7636 85018 -7454 85254
rect -7218 85018 -7036 85254
rect -7636 84934 -7036 85018
rect -7636 84698 -7454 84934
rect -7218 84698 -7036 84934
rect -7636 49254 -7036 84698
rect -7636 49018 -7454 49254
rect -7218 49018 -7036 49254
rect -7636 48934 -7036 49018
rect -7636 48698 -7454 48934
rect -7218 48698 -7036 48934
rect -7636 13254 -7036 48698
rect -7636 13018 -7454 13254
rect -7218 13018 -7036 13254
rect -7636 12934 -7036 13018
rect -7636 12698 -7454 12934
rect -7218 12698 -7036 12934
rect -7636 -5986 -7036 12698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 675654 -6096 708982
rect -6696 675418 -6514 675654
rect -6278 675418 -6096 675654
rect -6696 675334 -6096 675418
rect -6696 675098 -6514 675334
rect -6278 675098 -6096 675334
rect -6696 639654 -6096 675098
rect -6696 639418 -6514 639654
rect -6278 639418 -6096 639654
rect -6696 639334 -6096 639418
rect -6696 639098 -6514 639334
rect -6278 639098 -6096 639334
rect -6696 603654 -6096 639098
rect -6696 603418 -6514 603654
rect -6278 603418 -6096 603654
rect -6696 603334 -6096 603418
rect -6696 603098 -6514 603334
rect -6278 603098 -6096 603334
rect -6696 567654 -6096 603098
rect -6696 567418 -6514 567654
rect -6278 567418 -6096 567654
rect -6696 567334 -6096 567418
rect -6696 567098 -6514 567334
rect -6278 567098 -6096 567334
rect -6696 531654 -6096 567098
rect -6696 531418 -6514 531654
rect -6278 531418 -6096 531654
rect -6696 531334 -6096 531418
rect -6696 531098 -6514 531334
rect -6278 531098 -6096 531334
rect -6696 495654 -6096 531098
rect -6696 495418 -6514 495654
rect -6278 495418 -6096 495654
rect -6696 495334 -6096 495418
rect -6696 495098 -6514 495334
rect -6278 495098 -6096 495334
rect -6696 459654 -6096 495098
rect -6696 459418 -6514 459654
rect -6278 459418 -6096 459654
rect -6696 459334 -6096 459418
rect -6696 459098 -6514 459334
rect -6278 459098 -6096 459334
rect -6696 423654 -6096 459098
rect -6696 423418 -6514 423654
rect -6278 423418 -6096 423654
rect -6696 423334 -6096 423418
rect -6696 423098 -6514 423334
rect -6278 423098 -6096 423334
rect -6696 387654 -6096 423098
rect -6696 387418 -6514 387654
rect -6278 387418 -6096 387654
rect -6696 387334 -6096 387418
rect -6696 387098 -6514 387334
rect -6278 387098 -6096 387334
rect -6696 351654 -6096 387098
rect -6696 351418 -6514 351654
rect -6278 351418 -6096 351654
rect -6696 351334 -6096 351418
rect -6696 351098 -6514 351334
rect -6278 351098 -6096 351334
rect -6696 315654 -6096 351098
rect -6696 315418 -6514 315654
rect -6278 315418 -6096 315654
rect -6696 315334 -6096 315418
rect -6696 315098 -6514 315334
rect -6278 315098 -6096 315334
rect -6696 279654 -6096 315098
rect -6696 279418 -6514 279654
rect -6278 279418 -6096 279654
rect -6696 279334 -6096 279418
rect -6696 279098 -6514 279334
rect -6278 279098 -6096 279334
rect -6696 243654 -6096 279098
rect -6696 243418 -6514 243654
rect -6278 243418 -6096 243654
rect -6696 243334 -6096 243418
rect -6696 243098 -6514 243334
rect -6278 243098 -6096 243334
rect -6696 207654 -6096 243098
rect -6696 207418 -6514 207654
rect -6278 207418 -6096 207654
rect -6696 207334 -6096 207418
rect -6696 207098 -6514 207334
rect -6278 207098 -6096 207334
rect -6696 171654 -6096 207098
rect -6696 171418 -6514 171654
rect -6278 171418 -6096 171654
rect -6696 171334 -6096 171418
rect -6696 171098 -6514 171334
rect -6278 171098 -6096 171334
rect -6696 135654 -6096 171098
rect -6696 135418 -6514 135654
rect -6278 135418 -6096 135654
rect -6696 135334 -6096 135418
rect -6696 135098 -6514 135334
rect -6278 135098 -6096 135334
rect -6696 99654 -6096 135098
rect -6696 99418 -6514 99654
rect -6278 99418 -6096 99654
rect -6696 99334 -6096 99418
rect -6696 99098 -6514 99334
rect -6278 99098 -6096 99334
rect -6696 63654 -6096 99098
rect -6696 63418 -6514 63654
rect -6278 63418 -6096 63654
rect -6696 63334 -6096 63418
rect -6696 63098 -6514 63334
rect -6278 63098 -6096 63334
rect -6696 27654 -6096 63098
rect -6696 27418 -6514 27654
rect -6278 27418 -6096 27654
rect -6696 27334 -6096 27418
rect -6696 27098 -6514 27334
rect -6278 27098 -6096 27334
rect -6696 -5046 -6096 27098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 693654 -5156 708042
rect 8004 708598 8604 709560
rect 8004 708362 8186 708598
rect 8422 708362 8604 708598
rect 8004 708278 8604 708362
rect 8004 708042 8186 708278
rect 8422 708042 8604 708278
rect -5756 693418 -5574 693654
rect -5338 693418 -5156 693654
rect -5756 693334 -5156 693418
rect -5756 693098 -5574 693334
rect -5338 693098 -5156 693334
rect -5756 657654 -5156 693098
rect -5756 657418 -5574 657654
rect -5338 657418 -5156 657654
rect -5756 657334 -5156 657418
rect -5756 657098 -5574 657334
rect -5338 657098 -5156 657334
rect -5756 621654 -5156 657098
rect -5756 621418 -5574 621654
rect -5338 621418 -5156 621654
rect -5756 621334 -5156 621418
rect -5756 621098 -5574 621334
rect -5338 621098 -5156 621334
rect -5756 585654 -5156 621098
rect -5756 585418 -5574 585654
rect -5338 585418 -5156 585654
rect -5756 585334 -5156 585418
rect -5756 585098 -5574 585334
rect -5338 585098 -5156 585334
rect -5756 549654 -5156 585098
rect -5756 549418 -5574 549654
rect -5338 549418 -5156 549654
rect -5756 549334 -5156 549418
rect -5756 549098 -5574 549334
rect -5338 549098 -5156 549334
rect -5756 513654 -5156 549098
rect -5756 513418 -5574 513654
rect -5338 513418 -5156 513654
rect -5756 513334 -5156 513418
rect -5756 513098 -5574 513334
rect -5338 513098 -5156 513334
rect -5756 477654 -5156 513098
rect -5756 477418 -5574 477654
rect -5338 477418 -5156 477654
rect -5756 477334 -5156 477418
rect -5756 477098 -5574 477334
rect -5338 477098 -5156 477334
rect -5756 441654 -5156 477098
rect -5756 441418 -5574 441654
rect -5338 441418 -5156 441654
rect -5756 441334 -5156 441418
rect -5756 441098 -5574 441334
rect -5338 441098 -5156 441334
rect -5756 405654 -5156 441098
rect -5756 405418 -5574 405654
rect -5338 405418 -5156 405654
rect -5756 405334 -5156 405418
rect -5756 405098 -5574 405334
rect -5338 405098 -5156 405334
rect -5756 369654 -5156 405098
rect -5756 369418 -5574 369654
rect -5338 369418 -5156 369654
rect -5756 369334 -5156 369418
rect -5756 369098 -5574 369334
rect -5338 369098 -5156 369334
rect -5756 333654 -5156 369098
rect -5756 333418 -5574 333654
rect -5338 333418 -5156 333654
rect -5756 333334 -5156 333418
rect -5756 333098 -5574 333334
rect -5338 333098 -5156 333334
rect -5756 297654 -5156 333098
rect -5756 297418 -5574 297654
rect -5338 297418 -5156 297654
rect -5756 297334 -5156 297418
rect -5756 297098 -5574 297334
rect -5338 297098 -5156 297334
rect -5756 261654 -5156 297098
rect -5756 261418 -5574 261654
rect -5338 261418 -5156 261654
rect -5756 261334 -5156 261418
rect -5756 261098 -5574 261334
rect -5338 261098 -5156 261334
rect -5756 225654 -5156 261098
rect -5756 225418 -5574 225654
rect -5338 225418 -5156 225654
rect -5756 225334 -5156 225418
rect -5756 225098 -5574 225334
rect -5338 225098 -5156 225334
rect -5756 189654 -5156 225098
rect -5756 189418 -5574 189654
rect -5338 189418 -5156 189654
rect -5756 189334 -5156 189418
rect -5756 189098 -5574 189334
rect -5338 189098 -5156 189334
rect -5756 153654 -5156 189098
rect -5756 153418 -5574 153654
rect -5338 153418 -5156 153654
rect -5756 153334 -5156 153418
rect -5756 153098 -5574 153334
rect -5338 153098 -5156 153334
rect -5756 117654 -5156 153098
rect -5756 117418 -5574 117654
rect -5338 117418 -5156 117654
rect -5756 117334 -5156 117418
rect -5756 117098 -5574 117334
rect -5338 117098 -5156 117334
rect -5756 81654 -5156 117098
rect -5756 81418 -5574 81654
rect -5338 81418 -5156 81654
rect -5756 81334 -5156 81418
rect -5756 81098 -5574 81334
rect -5338 81098 -5156 81334
rect -5756 45654 -5156 81098
rect -5756 45418 -5574 45654
rect -5338 45418 -5156 45654
rect -5756 45334 -5156 45418
rect -5756 45098 -5574 45334
rect -5338 45098 -5156 45334
rect -5756 9654 -5156 45098
rect -5756 9418 -5574 9654
rect -5338 9418 -5156 9654
rect -5756 9334 -5156 9418
rect -5756 9098 -5574 9334
rect -5338 9098 -5156 9334
rect -5756 -4106 -5156 9098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 672054 -4216 707102
rect -4816 671818 -4634 672054
rect -4398 671818 -4216 672054
rect -4816 671734 -4216 671818
rect -4816 671498 -4634 671734
rect -4398 671498 -4216 671734
rect -4816 636054 -4216 671498
rect -4816 635818 -4634 636054
rect -4398 635818 -4216 636054
rect -4816 635734 -4216 635818
rect -4816 635498 -4634 635734
rect -4398 635498 -4216 635734
rect -4816 600054 -4216 635498
rect -4816 599818 -4634 600054
rect -4398 599818 -4216 600054
rect -4816 599734 -4216 599818
rect -4816 599498 -4634 599734
rect -4398 599498 -4216 599734
rect -4816 564054 -4216 599498
rect -4816 563818 -4634 564054
rect -4398 563818 -4216 564054
rect -4816 563734 -4216 563818
rect -4816 563498 -4634 563734
rect -4398 563498 -4216 563734
rect -4816 528054 -4216 563498
rect -4816 527818 -4634 528054
rect -4398 527818 -4216 528054
rect -4816 527734 -4216 527818
rect -4816 527498 -4634 527734
rect -4398 527498 -4216 527734
rect -4816 492054 -4216 527498
rect -4816 491818 -4634 492054
rect -4398 491818 -4216 492054
rect -4816 491734 -4216 491818
rect -4816 491498 -4634 491734
rect -4398 491498 -4216 491734
rect -4816 456054 -4216 491498
rect -4816 455818 -4634 456054
rect -4398 455818 -4216 456054
rect -4816 455734 -4216 455818
rect -4816 455498 -4634 455734
rect -4398 455498 -4216 455734
rect -4816 420054 -4216 455498
rect -4816 419818 -4634 420054
rect -4398 419818 -4216 420054
rect -4816 419734 -4216 419818
rect -4816 419498 -4634 419734
rect -4398 419498 -4216 419734
rect -4816 384054 -4216 419498
rect -4816 383818 -4634 384054
rect -4398 383818 -4216 384054
rect -4816 383734 -4216 383818
rect -4816 383498 -4634 383734
rect -4398 383498 -4216 383734
rect -4816 348054 -4216 383498
rect -4816 347818 -4634 348054
rect -4398 347818 -4216 348054
rect -4816 347734 -4216 347818
rect -4816 347498 -4634 347734
rect -4398 347498 -4216 347734
rect -4816 312054 -4216 347498
rect -4816 311818 -4634 312054
rect -4398 311818 -4216 312054
rect -4816 311734 -4216 311818
rect -4816 311498 -4634 311734
rect -4398 311498 -4216 311734
rect -4816 276054 -4216 311498
rect -4816 275818 -4634 276054
rect -4398 275818 -4216 276054
rect -4816 275734 -4216 275818
rect -4816 275498 -4634 275734
rect -4398 275498 -4216 275734
rect -4816 240054 -4216 275498
rect -4816 239818 -4634 240054
rect -4398 239818 -4216 240054
rect -4816 239734 -4216 239818
rect -4816 239498 -4634 239734
rect -4398 239498 -4216 239734
rect -4816 204054 -4216 239498
rect -4816 203818 -4634 204054
rect -4398 203818 -4216 204054
rect -4816 203734 -4216 203818
rect -4816 203498 -4634 203734
rect -4398 203498 -4216 203734
rect -4816 168054 -4216 203498
rect -4816 167818 -4634 168054
rect -4398 167818 -4216 168054
rect -4816 167734 -4216 167818
rect -4816 167498 -4634 167734
rect -4398 167498 -4216 167734
rect -4816 132054 -4216 167498
rect -4816 131818 -4634 132054
rect -4398 131818 -4216 132054
rect -4816 131734 -4216 131818
rect -4816 131498 -4634 131734
rect -4398 131498 -4216 131734
rect -4816 96054 -4216 131498
rect -4816 95818 -4634 96054
rect -4398 95818 -4216 96054
rect -4816 95734 -4216 95818
rect -4816 95498 -4634 95734
rect -4398 95498 -4216 95734
rect -4816 60054 -4216 95498
rect -4816 59818 -4634 60054
rect -4398 59818 -4216 60054
rect -4816 59734 -4216 59818
rect -4816 59498 -4634 59734
rect -4398 59498 -4216 59734
rect -4816 24054 -4216 59498
rect -4816 23818 -4634 24054
rect -4398 23818 -4216 24054
rect -4816 23734 -4216 23818
rect -4816 23498 -4634 23734
rect -4398 23498 -4216 23734
rect -4816 -3166 -4216 23498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 690054 -3276 706162
rect 4404 706718 5004 707680
rect 4404 706482 4586 706718
rect 4822 706482 5004 706718
rect 4404 706398 5004 706482
rect 4404 706162 4586 706398
rect 4822 706162 5004 706398
rect -3876 689818 -3694 690054
rect -3458 689818 -3276 690054
rect -3876 689734 -3276 689818
rect -3876 689498 -3694 689734
rect -3458 689498 -3276 689734
rect -3876 654054 -3276 689498
rect -3876 653818 -3694 654054
rect -3458 653818 -3276 654054
rect -3876 653734 -3276 653818
rect -3876 653498 -3694 653734
rect -3458 653498 -3276 653734
rect -3876 618054 -3276 653498
rect -3876 617818 -3694 618054
rect -3458 617818 -3276 618054
rect -3876 617734 -3276 617818
rect -3876 617498 -3694 617734
rect -3458 617498 -3276 617734
rect -3876 582054 -3276 617498
rect -3876 581818 -3694 582054
rect -3458 581818 -3276 582054
rect -3876 581734 -3276 581818
rect -3876 581498 -3694 581734
rect -3458 581498 -3276 581734
rect -3876 546054 -3276 581498
rect -3876 545818 -3694 546054
rect -3458 545818 -3276 546054
rect -3876 545734 -3276 545818
rect -3876 545498 -3694 545734
rect -3458 545498 -3276 545734
rect -3876 510054 -3276 545498
rect -3876 509818 -3694 510054
rect -3458 509818 -3276 510054
rect -3876 509734 -3276 509818
rect -3876 509498 -3694 509734
rect -3458 509498 -3276 509734
rect -3876 474054 -3276 509498
rect -3876 473818 -3694 474054
rect -3458 473818 -3276 474054
rect -3876 473734 -3276 473818
rect -3876 473498 -3694 473734
rect -3458 473498 -3276 473734
rect -3876 438054 -3276 473498
rect -3876 437818 -3694 438054
rect -3458 437818 -3276 438054
rect -3876 437734 -3276 437818
rect -3876 437498 -3694 437734
rect -3458 437498 -3276 437734
rect -3876 402054 -3276 437498
rect -3876 401818 -3694 402054
rect -3458 401818 -3276 402054
rect -3876 401734 -3276 401818
rect -3876 401498 -3694 401734
rect -3458 401498 -3276 401734
rect -3876 366054 -3276 401498
rect -3876 365818 -3694 366054
rect -3458 365818 -3276 366054
rect -3876 365734 -3276 365818
rect -3876 365498 -3694 365734
rect -3458 365498 -3276 365734
rect -3876 330054 -3276 365498
rect -3876 329818 -3694 330054
rect -3458 329818 -3276 330054
rect -3876 329734 -3276 329818
rect -3876 329498 -3694 329734
rect -3458 329498 -3276 329734
rect -3876 294054 -3276 329498
rect -3876 293818 -3694 294054
rect -3458 293818 -3276 294054
rect -3876 293734 -3276 293818
rect -3876 293498 -3694 293734
rect -3458 293498 -3276 293734
rect -3876 258054 -3276 293498
rect -3876 257818 -3694 258054
rect -3458 257818 -3276 258054
rect -3876 257734 -3276 257818
rect -3876 257498 -3694 257734
rect -3458 257498 -3276 257734
rect -3876 222054 -3276 257498
rect -3876 221818 -3694 222054
rect -3458 221818 -3276 222054
rect -3876 221734 -3276 221818
rect -3876 221498 -3694 221734
rect -3458 221498 -3276 221734
rect -3876 186054 -3276 221498
rect -3876 185818 -3694 186054
rect -3458 185818 -3276 186054
rect -3876 185734 -3276 185818
rect -3876 185498 -3694 185734
rect -3458 185498 -3276 185734
rect -3876 150054 -3276 185498
rect -3876 149818 -3694 150054
rect -3458 149818 -3276 150054
rect -3876 149734 -3276 149818
rect -3876 149498 -3694 149734
rect -3458 149498 -3276 149734
rect -3876 114054 -3276 149498
rect -3876 113818 -3694 114054
rect -3458 113818 -3276 114054
rect -3876 113734 -3276 113818
rect -3876 113498 -3694 113734
rect -3458 113498 -3276 113734
rect -3876 78054 -3276 113498
rect -3876 77818 -3694 78054
rect -3458 77818 -3276 78054
rect -3876 77734 -3276 77818
rect -3876 77498 -3694 77734
rect -3458 77498 -3276 77734
rect -3876 42054 -3276 77498
rect -3876 41818 -3694 42054
rect -3458 41818 -3276 42054
rect -3876 41734 -3276 41818
rect -3876 41498 -3694 41734
rect -3458 41498 -3276 41734
rect -3876 6054 -3276 41498
rect -3876 5818 -3694 6054
rect -3458 5818 -3276 6054
rect -3876 5734 -3276 5818
rect -3876 5498 -3694 5734
rect -3458 5498 -3276 5734
rect -3876 -2226 -3276 5498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 4404 690054 5004 706162
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 4404 -2226 5004 5498
rect 4404 -2462 4586 -2226
rect 4822 -2462 5004 -2226
rect 4404 -2546 5004 -2462
rect 4404 -2782 4586 -2546
rect 4822 -2782 5004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 4404 -3744 5004 -2782
rect 8004 693654 8604 708042
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 8004 -4106 8604 9098
rect 8004 -4342 8186 -4106
rect 8422 -4342 8604 -4106
rect 8004 -4426 8604 -4342
rect 8004 -4662 8186 -4426
rect 8422 -4662 8604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 8004 -5624 8604 -4662
rect 11604 697254 12204 709922
rect 29604 711418 30204 711440
rect 29604 711182 29786 711418
rect 30022 711182 30204 711418
rect 29604 711098 30204 711182
rect 29604 710862 29786 711098
rect 30022 710862 30204 711098
rect 26004 709538 26604 709560
rect 26004 709302 26186 709538
rect 26422 709302 26604 709538
rect 26004 709218 26604 709302
rect 26004 708982 26186 709218
rect 26422 708982 26604 709218
rect 22404 707658 23004 707680
rect 22404 707422 22586 707658
rect 22822 707422 23004 707658
rect 22404 707338 23004 707422
rect 22404 707102 22586 707338
rect 22822 707102 23004 707338
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 11604 -5986 12204 12698
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 22404 672054 23004 707102
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3166 23004 23498
rect 22404 -3402 22586 -3166
rect 22822 -3402 23004 -3166
rect 22404 -3486 23004 -3402
rect 22404 -3722 22586 -3486
rect 22822 -3722 23004 -3486
rect 22404 -3744 23004 -3722
rect 26004 675654 26604 708982
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -5046 26604 27098
rect 26004 -5282 26186 -5046
rect 26422 -5282 26604 -5046
rect 26004 -5366 26604 -5282
rect 26004 -5602 26186 -5366
rect 26422 -5602 26604 -5366
rect 26004 -5624 26604 -5602
rect 29604 679254 30204 710862
rect 47604 710478 48204 711440
rect 47604 710242 47786 710478
rect 48022 710242 48204 710478
rect 47604 710158 48204 710242
rect 47604 709922 47786 710158
rect 48022 709922 48204 710158
rect 44004 708598 44604 709560
rect 44004 708362 44186 708598
rect 44422 708362 44604 708598
rect 44004 708278 44604 708362
rect 44004 708042 44186 708278
rect 44422 708042 44604 708278
rect 40404 706718 41004 707680
rect 40404 706482 40586 706718
rect 40822 706482 41004 706718
rect 40404 706398 41004 706482
rect 40404 706162 40586 706398
rect 40822 706162 41004 706398
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6222 11786 -5986
rect 12022 -6222 12204 -5986
rect 11604 -6306 12204 -6222
rect 11604 -6542 11786 -6306
rect 12022 -6542 12204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 11604 -7504 12204 -6542
rect 29604 -6926 30204 30698
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 40404 690054 41004 706162
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2226 41004 5498
rect 40404 -2462 40586 -2226
rect 40822 -2462 41004 -2226
rect 40404 -2546 41004 -2462
rect 40404 -2782 40586 -2546
rect 40822 -2782 41004 -2546
rect 40404 -3744 41004 -2782
rect 44004 693654 44604 708042
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4106 44604 9098
rect 44004 -4342 44186 -4106
rect 44422 -4342 44604 -4106
rect 44004 -4426 44604 -4342
rect 44004 -4662 44186 -4426
rect 44422 -4662 44604 -4426
rect 44004 -5624 44604 -4662
rect 47604 697254 48204 709922
rect 65604 711418 66204 711440
rect 65604 711182 65786 711418
rect 66022 711182 66204 711418
rect 65604 711098 66204 711182
rect 65604 710862 65786 711098
rect 66022 710862 66204 711098
rect 62004 709538 62604 709560
rect 62004 709302 62186 709538
rect 62422 709302 62604 709538
rect 62004 709218 62604 709302
rect 62004 708982 62186 709218
rect 62422 708982 62604 709218
rect 58404 707658 59004 707680
rect 58404 707422 58586 707658
rect 58822 707422 59004 707658
rect 58404 707338 59004 707422
rect 58404 707102 58586 707338
rect 58822 707102 59004 707338
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7162 29786 -6926
rect 30022 -7162 30204 -6926
rect 29604 -7246 30204 -7162
rect 29604 -7482 29786 -7246
rect 30022 -7482 30204 -7246
rect 29604 -7504 30204 -7482
rect 47604 -5986 48204 12698
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 58404 672054 59004 707102
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3166 59004 23498
rect 58404 -3402 58586 -3166
rect 58822 -3402 59004 -3166
rect 58404 -3486 59004 -3402
rect 58404 -3722 58586 -3486
rect 58822 -3722 59004 -3486
rect 58404 -3744 59004 -3722
rect 62004 675654 62604 708982
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -5046 62604 27098
rect 62004 -5282 62186 -5046
rect 62422 -5282 62604 -5046
rect 62004 -5366 62604 -5282
rect 62004 -5602 62186 -5366
rect 62422 -5602 62604 -5366
rect 62004 -5624 62604 -5602
rect 65604 679254 66204 710862
rect 83604 710478 84204 711440
rect 83604 710242 83786 710478
rect 84022 710242 84204 710478
rect 83604 710158 84204 710242
rect 83604 709922 83786 710158
rect 84022 709922 84204 710158
rect 80004 708598 80604 709560
rect 80004 708362 80186 708598
rect 80422 708362 80604 708598
rect 80004 708278 80604 708362
rect 80004 708042 80186 708278
rect 80422 708042 80604 708278
rect 76404 706718 77004 707680
rect 76404 706482 76586 706718
rect 76822 706482 77004 706718
rect 76404 706398 77004 706482
rect 76404 706162 76586 706398
rect 76822 706162 77004 706398
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 396550 73404 397898
rect 76404 690054 77004 706162
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 396550 77004 401498
rect 80004 693654 80604 708042
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 396550 80604 405098
rect 83604 697254 84204 709922
rect 101604 711418 102204 711440
rect 101604 711182 101786 711418
rect 102022 711182 102204 711418
rect 101604 711098 102204 711182
rect 101604 710862 101786 711098
rect 102022 710862 102204 711098
rect 98004 709538 98604 709560
rect 98004 709302 98186 709538
rect 98422 709302 98604 709538
rect 98004 709218 98604 709302
rect 98004 708982 98186 709218
rect 98422 708982 98604 709218
rect 94404 707658 95004 707680
rect 94404 707422 94586 707658
rect 94822 707422 95004 707658
rect 94404 707338 95004 707422
rect 94404 707102 94586 707338
rect 94822 707102 95004 707338
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 552104 91404 559898
rect 94404 672054 95004 707102
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 552104 95004 563498
rect 98004 675654 98604 708982
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 552104 98604 567098
rect 101604 679254 102204 710862
rect 119604 710478 120204 711440
rect 119604 710242 119786 710478
rect 120022 710242 120204 710478
rect 119604 710158 120204 710242
rect 119604 709922 119786 710158
rect 120022 709922 120204 710158
rect 116004 708598 116604 709560
rect 116004 708362 116186 708598
rect 116422 708362 116604 708598
rect 116004 708278 116604 708362
rect 116004 708042 116186 708278
rect 116422 708042 116604 708278
rect 112404 706718 113004 707680
rect 112404 706482 112586 706718
rect 112822 706482 113004 706718
rect 112404 706398 113004 706482
rect 112404 706162 112586 706398
rect 112822 706162 113004 706398
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 552104 102204 570698
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 552104 109404 577898
rect 112404 690054 113004 706162
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 552104 113004 581498
rect 116004 693654 116604 708042
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 91529 542454 91849 542476
rect 91529 542218 91571 542454
rect 91807 542218 91849 542454
rect 91529 542134 91849 542218
rect 91529 541898 91571 542134
rect 91807 541898 91849 542134
rect 91529 541876 91849 541898
rect 96113 524454 96433 524476
rect 96113 524218 96155 524454
rect 96391 524218 96433 524454
rect 96113 524134 96433 524218
rect 96113 523898 96155 524134
rect 96391 523898 96433 524134
rect 96113 523876 96433 523898
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 396550 84204 408698
rect 90804 488454 91404 519800
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 396550 91404 415898
rect 94404 492054 95004 519800
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 396550 95004 419498
rect 98004 495654 98604 519800
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 396550 98604 423098
rect 101604 499254 102204 519800
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 396550 102204 426698
rect 108804 506454 109404 519800
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 396550 109404 397898
rect 112404 510054 113004 519800
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 396550 113004 401498
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 396550 116604 405098
rect 119604 697254 120204 709922
rect 137604 711418 138204 711440
rect 137604 711182 137786 711418
rect 138022 711182 138204 711418
rect 137604 711098 138204 711182
rect 137604 710862 137786 711098
rect 138022 710862 138204 711098
rect 134004 709538 134604 709560
rect 134004 709302 134186 709538
rect 134422 709302 134604 709538
rect 134004 709218 134604 709302
rect 134004 708982 134186 709218
rect 134422 708982 134604 709218
rect 130404 707658 131004 707680
rect 130404 707422 130586 707658
rect 130822 707422 131004 707658
rect 130404 707338 131004 707422
rect 130404 707102 130586 707338
rect 130822 707102 131004 707338
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 553254 120204 588698
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 396550 120204 408698
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 91568 380454 91888 380476
rect 91568 380218 91610 380454
rect 91846 380218 91888 380454
rect 91568 380134 91888 380218
rect 91568 379898 91610 380134
rect 91846 379898 91888 380134
rect 91568 379876 91888 379898
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 76208 362454 76528 362476
rect 76208 362218 76250 362454
rect 76486 362218 76528 362454
rect 76208 362134 76528 362218
rect 76208 361898 76250 362134
rect 76486 361898 76528 362134
rect 76208 361876 76528 361898
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 91568 344454 91888 344476
rect 91568 344218 91610 344454
rect 91846 344218 91888 344454
rect 91568 344134 91888 344218
rect 91568 343898 91610 344134
rect 91846 343898 91888 344134
rect 91568 343876 91888 343898
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6222 47786 -5986
rect 48022 -6222 48204 -5986
rect 47604 -6306 48204 -6222
rect 47604 -6542 47786 -6306
rect 48022 -6542 48204 -6306
rect 47604 -7504 48204 -6542
rect 65604 -6926 66204 30698
rect 72804 326454 73404 339800
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 76404 330054 77004 339800
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2226 77004 5498
rect 76404 -2462 76586 -2226
rect 76822 -2462 77004 -2226
rect 76404 -2546 77004 -2462
rect 76404 -2782 76586 -2546
rect 76822 -2782 77004 -2546
rect 76404 -3744 77004 -2782
rect 80004 333654 80604 339800
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4106 80604 9098
rect 80004 -4342 80186 -4106
rect 80422 -4342 80604 -4106
rect 80004 -4426 80604 -4342
rect 80004 -4662 80186 -4426
rect 80422 -4662 80604 -4426
rect 80004 -5624 80604 -4662
rect 83604 337254 84204 339800
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7162 65786 -6926
rect 66022 -7162 66204 -6926
rect 65604 -7246 66204 -7162
rect 65604 -7482 65786 -7246
rect 66022 -7482 66204 -7246
rect 65604 -7504 66204 -7482
rect 83604 -5986 84204 12698
rect 90804 308454 91404 339800
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 94404 312054 95004 339800
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3166 95004 23498
rect 94404 -3402 94586 -3166
rect 94822 -3402 95004 -3166
rect 94404 -3486 95004 -3402
rect 94404 -3722 94586 -3486
rect 94822 -3722 95004 -3486
rect 94404 -3744 95004 -3722
rect 98004 315654 98604 339800
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -5046 98604 27098
rect 98004 -5282 98186 -5046
rect 98422 -5282 98604 -5046
rect 98004 -5366 98604 -5282
rect 98004 -5602 98186 -5366
rect 98422 -5602 98604 -5366
rect 98004 -5624 98604 -5602
rect 101604 319254 102204 339800
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6222 83786 -5986
rect 84022 -6222 84204 -5986
rect 83604 -6306 84204 -6222
rect 83604 -6542 83786 -6306
rect 84022 -6542 84204 -6306
rect 83604 -7504 84204 -6542
rect 101604 -6926 102204 30698
rect 108804 326454 109404 339800
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 112404 330054 113004 339800
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2226 113004 5498
rect 112404 -2462 112586 -2226
rect 112822 -2462 113004 -2226
rect 112404 -2546 113004 -2462
rect 112404 -2782 112586 -2546
rect 112822 -2782 113004 -2546
rect 112404 -3744 113004 -2782
rect 116004 333654 116604 339800
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4106 116604 9098
rect 116004 -4342 116186 -4106
rect 116422 -4342 116604 -4106
rect 116004 -4426 116604 -4342
rect 116004 -4662 116186 -4426
rect 116422 -4662 116604 -4426
rect 116004 -5624 116604 -4662
rect 119604 337254 120204 339800
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7162 101786 -6926
rect 102022 -7162 102204 -6926
rect 101604 -7246 102204 -7162
rect 101604 -7482 101786 -7246
rect 102022 -7482 102204 -7246
rect 101604 -7504 102204 -7482
rect 119604 -5986 120204 12698
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 130404 672054 131004 707102
rect 132171 700500 132237 700501
rect 132171 700436 132172 700500
rect 132236 700436 132237 700500
rect 132171 700435 132237 700436
rect 131987 685948 132053 685949
rect 131987 685884 131988 685948
rect 132052 685884 132053 685948
rect 131987 685883 132053 685884
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 131803 639028 131869 639029
rect 131803 638964 131804 639028
rect 131868 638964 131869 639028
rect 131803 638963 131869 638964
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 128859 299300 128925 299301
rect 128859 299236 128860 299300
rect 128924 299236 128925 299300
rect 128859 299235 128925 299236
rect 128862 289917 128922 299235
rect 128859 289916 128925 289917
rect 128859 289852 128860 289916
rect 128924 289852 128925 289916
rect 128859 289851 128925 289852
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 131806 134061 131866 638963
rect 131990 135149 132050 685883
rect 132174 137189 132234 700435
rect 132355 700364 132421 700365
rect 132355 700300 132356 700364
rect 132420 700300 132421 700364
rect 132355 700299 132421 700300
rect 132171 137188 132237 137189
rect 132171 137124 132172 137188
rect 132236 137124 132237 137188
rect 132171 137123 132237 137124
rect 132358 136237 132418 700299
rect 133643 697236 133709 697237
rect 133643 697172 133644 697236
rect 133708 697172 133709 697236
rect 133643 697171 133709 697172
rect 133459 650316 133525 650317
rect 133459 650252 133460 650316
rect 133524 650252 133525 650316
rect 133459 650251 133525 650252
rect 133091 603396 133157 603397
rect 133091 603332 133092 603396
rect 133156 603332 133157 603396
rect 133091 603331 133157 603332
rect 132907 200700 132973 200701
rect 132907 200636 132908 200700
rect 132972 200636 132973 200700
rect 132907 200635 132973 200636
rect 132910 176221 132970 200635
rect 132907 176220 132973 176221
rect 132907 176156 132908 176220
rect 132972 176156 132973 176220
rect 132907 176155 132973 176156
rect 133094 172957 133154 603331
rect 133275 592380 133341 592381
rect 133275 592316 133276 592380
rect 133340 592316 133341 592380
rect 133275 592315 133341 592316
rect 133091 172956 133157 172957
rect 133091 172892 133092 172956
rect 133156 172892 133157 172956
rect 133091 172891 133157 172892
rect 132355 136236 132421 136237
rect 132355 136172 132356 136236
rect 132420 136172 132421 136236
rect 132355 136171 132421 136172
rect 131987 135148 132053 135149
rect 131987 135084 131988 135148
rect 132052 135084 132053 135148
rect 131987 135083 132053 135084
rect 131803 134060 131869 134061
rect 131803 133996 131804 134060
rect 131868 133996 131869 134060
rect 131803 133995 131869 133996
rect 133278 132973 133338 592315
rect 133462 174045 133522 650251
rect 133646 175133 133706 697171
rect 134004 675654 134604 708982
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 134004 200200 134604 207098
rect 137604 679254 138204 710862
rect 155604 710478 156204 711440
rect 155604 710242 155786 710478
rect 156022 710242 156204 710478
rect 155604 710158 156204 710242
rect 155604 709922 155786 710158
rect 156022 709922 156204 710158
rect 152004 708598 152604 709560
rect 152004 708362 152186 708598
rect 152422 708362 152604 708598
rect 152004 708278 152604 708362
rect 152004 708042 152186 708278
rect 152422 708042 152604 708278
rect 148404 706718 149004 707680
rect 148404 706482 148586 706718
rect 148822 706482 149004 706718
rect 148404 706398 149004 706482
rect 148404 706162 148586 706398
rect 148822 706162 149004 706398
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 535254 138204 570698
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 200200 138204 210698
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 200200 145404 217898
rect 148404 690054 149004 706162
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 200200 149004 221498
rect 152004 693654 152604 708042
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 200200 152604 225098
rect 155604 697254 156204 709922
rect 173604 711418 174204 711440
rect 173604 711182 173786 711418
rect 174022 711182 174204 711418
rect 173604 711098 174204 711182
rect 173604 710862 173786 711098
rect 174022 710862 174204 711098
rect 170004 709538 170604 709560
rect 170004 709302 170186 709538
rect 170422 709302 170604 709538
rect 170004 709218 170604 709302
rect 170004 708982 170186 709218
rect 170422 708982 170604 709218
rect 166404 707658 167004 707680
rect 166404 707422 166586 707658
rect 166822 707422 167004 707658
rect 166404 707338 167004 707422
rect 166404 707102 166586 707338
rect 166822 707102 167004 707338
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 155604 409254 156204 444698
rect 155604 409018 155786 409254
rect 156022 409018 156204 409254
rect 155604 408934 156204 409018
rect 155604 408698 155786 408934
rect 156022 408698 156204 408934
rect 155604 373254 156204 408698
rect 155604 373018 155786 373254
rect 156022 373018 156204 373254
rect 155604 372934 156204 373018
rect 155604 372698 155786 372934
rect 156022 372698 156204 372934
rect 155604 337254 156204 372698
rect 155604 337018 155786 337254
rect 156022 337018 156204 337254
rect 155604 336934 156204 337018
rect 155604 336698 155786 336934
rect 156022 336698 156204 336934
rect 155604 301254 156204 336698
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 200200 156204 228698
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 164187 686492 164253 686493
rect 164187 686428 164188 686492
rect 164252 686428 164253 686492
rect 164187 686427 164253 686428
rect 164190 686221 164250 686427
rect 164187 686220 164253 686221
rect 164187 686156 164188 686220
rect 164252 686156 164253 686220
rect 164187 686155 164253 686156
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 166404 672054 167004 707102
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 164187 650588 164253 650589
rect 164187 650524 164188 650588
rect 164252 650524 164253 650588
rect 164187 650523 164253 650524
rect 164190 650317 164250 650523
rect 164187 650316 164253 650317
rect 164187 650252 164188 650316
rect 164252 650252 164253 650316
rect 164187 650251 164253 650252
rect 164187 639164 164253 639165
rect 164187 639100 164188 639164
rect 164252 639100 164253 639164
rect 164187 639099 164253 639100
rect 164190 638893 164250 639099
rect 164187 638892 164253 638893
rect 164187 638828 164188 638892
rect 164252 638828 164253 638892
rect 164187 638827 164253 638828
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 164187 603260 164253 603261
rect 164187 603196 164188 603260
rect 164252 603196 164253 603260
rect 164187 603195 164253 603196
rect 164190 602989 164250 603195
rect 164187 602988 164253 602989
rect 164187 602924 164188 602988
rect 164252 602924 164253 602988
rect 164187 602923 164253 602924
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 164187 592244 164253 592245
rect 164187 592180 164188 592244
rect 164252 592180 164253 592244
rect 164187 592179 164253 592180
rect 164190 591973 164250 592179
rect 164187 591972 164253 591973
rect 164187 591908 164188 591972
rect 164252 591908 164253 591972
rect 164187 591907 164253 591908
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200200 163404 235898
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 384054 167004 419498
rect 166404 383818 166586 384054
rect 166822 383818 167004 384054
rect 166404 383734 167004 383818
rect 166404 383498 166586 383734
rect 166822 383498 167004 383734
rect 166404 348054 167004 383498
rect 166404 347818 166586 348054
rect 166822 347818 167004 348054
rect 166404 347734 167004 347818
rect 166404 347498 166586 347734
rect 166822 347498 167004 347734
rect 166404 312054 167004 347498
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 200200 167004 203498
rect 170004 675654 170604 708982
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 387654 170604 423098
rect 170004 387418 170186 387654
rect 170422 387418 170604 387654
rect 170004 387334 170604 387418
rect 170004 387098 170186 387334
rect 170422 387098 170604 387334
rect 170004 351654 170604 387098
rect 170004 351418 170186 351654
rect 170422 351418 170604 351654
rect 170004 351334 170604 351418
rect 170004 351098 170186 351334
rect 170422 351098 170604 351334
rect 170004 315654 170604 351098
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 200200 170604 207098
rect 173604 679254 174204 710862
rect 191604 710478 192204 711440
rect 191604 710242 191786 710478
rect 192022 710242 192204 710478
rect 191604 710158 192204 710242
rect 191604 709922 191786 710158
rect 192022 709922 192204 710158
rect 188004 708598 188604 709560
rect 188004 708362 188186 708598
rect 188422 708362 188604 708598
rect 188004 708278 188604 708362
rect 188004 708042 188186 708278
rect 188422 708042 188604 708278
rect 184404 706718 185004 707680
rect 184404 706482 184586 706718
rect 184822 706482 185004 706718
rect 184404 706398 185004 706482
rect 184404 706162 184586 706398
rect 184822 706162 185004 706398
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 391254 174204 426698
rect 173604 391018 173786 391254
rect 174022 391018 174204 391254
rect 173604 390934 174204 391018
rect 173604 390698 173786 390934
rect 174022 390698 174204 390934
rect 173604 355254 174204 390698
rect 173604 355018 173786 355254
rect 174022 355018 174204 355254
rect 173604 354934 174204 355018
rect 173604 354698 173786 354934
rect 174022 354698 174204 354934
rect 173604 319254 174204 354698
rect 173604 319018 173786 319254
rect 174022 319018 174204 319254
rect 173604 318934 174204 319018
rect 173604 318698 173786 318934
rect 174022 318698 174204 318934
rect 173604 283254 174204 318698
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 200200 174204 210698
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 200200 181404 217898
rect 184404 690054 185004 706162
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 402054 185004 437498
rect 184404 401818 184586 402054
rect 184822 401818 185004 402054
rect 184404 401734 185004 401818
rect 184404 401498 184586 401734
rect 184822 401498 185004 401734
rect 184404 366054 185004 401498
rect 184404 365818 184586 366054
rect 184822 365818 185004 366054
rect 184404 365734 185004 365818
rect 184404 365498 184586 365734
rect 184822 365498 185004 365734
rect 184404 330054 185004 365498
rect 184404 329818 184586 330054
rect 184822 329818 185004 330054
rect 184404 329734 185004 329818
rect 184404 329498 184586 329734
rect 184822 329498 185004 329734
rect 184404 294054 185004 329498
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 200200 185004 221498
rect 188004 693654 188604 708042
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 405654 188604 441098
rect 188004 405418 188186 405654
rect 188422 405418 188604 405654
rect 188004 405334 188604 405418
rect 188004 405098 188186 405334
rect 188422 405098 188604 405334
rect 188004 369654 188604 405098
rect 188004 369418 188186 369654
rect 188422 369418 188604 369654
rect 188004 369334 188604 369418
rect 188004 369098 188186 369334
rect 188422 369098 188604 369334
rect 188004 333654 188604 369098
rect 188004 333418 188186 333654
rect 188422 333418 188604 333654
rect 188004 333334 188604 333418
rect 188004 333098 188186 333334
rect 188422 333098 188604 333334
rect 188004 297654 188604 333098
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 200200 188604 225098
rect 191604 697254 192204 709922
rect 209604 711418 210204 711440
rect 209604 711182 209786 711418
rect 210022 711182 210204 711418
rect 209604 711098 210204 711182
rect 209604 710862 209786 711098
rect 210022 710862 210204 711098
rect 206004 709538 206604 709560
rect 206004 709302 206186 709538
rect 206422 709302 206604 709538
rect 206004 709218 206604 709302
rect 206004 708982 206186 709218
rect 206422 708982 206604 709218
rect 202404 707658 203004 707680
rect 202404 707422 202586 707658
rect 202822 707422 203004 707658
rect 202404 707338 203004 707422
rect 202404 707102 202586 707338
rect 202822 707102 203004 707338
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 202404 672054 203004 707102
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 199699 561780 199765 561781
rect 199699 561716 199700 561780
rect 199764 561716 199765 561780
rect 199699 561715 199765 561716
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198595 556748 198661 556749
rect 198595 556684 198596 556748
rect 198660 556684 198661 556748
rect 198595 556683 198661 556684
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 198411 552124 198477 552125
rect 198411 552060 198412 552124
rect 198476 552060 198477 552124
rect 198411 552059 198477 552060
rect 198227 547908 198293 547909
rect 198227 547844 198228 547908
rect 198292 547844 198293 547908
rect 198227 547843 198293 547844
rect 198043 543828 198109 543829
rect 198043 543764 198044 543828
rect 198108 543764 198109 543828
rect 198043 543763 198109 543764
rect 197859 538524 197925 538525
rect 197859 538460 197860 538524
rect 197924 538460 197925 538524
rect 197859 538459 197925 538460
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 409254 192204 444698
rect 191604 409018 191786 409254
rect 192022 409018 192204 409254
rect 191604 408934 192204 409018
rect 191604 408698 191786 408934
rect 192022 408698 192204 408934
rect 191604 373254 192204 408698
rect 191604 373018 191786 373254
rect 192022 373018 192204 373254
rect 191604 372934 192204 373018
rect 191604 372698 191786 372934
rect 192022 372698 192204 372934
rect 191604 337254 192204 372698
rect 191604 337018 191786 337254
rect 192022 337018 192204 337254
rect 191604 336934 192204 337018
rect 191604 336698 191786 336934
rect 192022 336698 192204 336934
rect 191604 301254 192204 336698
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 200200 192204 228698
rect 197862 202605 197922 538459
rect 197859 202604 197925 202605
rect 197859 202540 197860 202604
rect 197924 202540 197925 202604
rect 197859 202539 197925 202540
rect 198046 201653 198106 543763
rect 198230 202333 198290 547843
rect 198227 202332 198293 202333
rect 198227 202268 198228 202332
rect 198292 202268 198293 202332
rect 198227 202267 198293 202268
rect 198414 201925 198474 552059
rect 198411 201924 198477 201925
rect 198411 201860 198412 201924
rect 198476 201860 198477 201924
rect 198411 201859 198477 201860
rect 198598 201789 198658 556683
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198595 201788 198661 201789
rect 198595 201724 198596 201788
rect 198660 201724 198661 201788
rect 198595 201723 198661 201724
rect 198043 201652 198109 201653
rect 198043 201588 198044 201652
rect 198108 201588 198109 201652
rect 198043 201587 198109 201588
rect 198804 200200 199404 235898
rect 199702 202061 199762 561715
rect 202404 560200 203004 563498
rect 206004 675654 206604 708982
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 560200 206604 567098
rect 209604 679254 210204 710862
rect 227604 710478 228204 711440
rect 227604 710242 227786 710478
rect 228022 710242 228204 710478
rect 227604 710158 228204 710242
rect 227604 709922 227786 710158
rect 228022 709922 228204 710158
rect 224004 708598 224604 709560
rect 224004 708362 224186 708598
rect 224422 708362 224604 708598
rect 224004 708278 224604 708362
rect 224004 708042 224186 708278
rect 224422 708042 224604 708278
rect 220404 706718 221004 707680
rect 220404 706482 220586 706718
rect 220822 706482 221004 706718
rect 220404 706398 221004 706482
rect 220404 706162 220586 706398
rect 220822 706162 221004 706398
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 560200 210204 570698
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 560200 217404 577898
rect 220404 690054 221004 706162
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 203909 542454 204229 542476
rect 203909 542218 203951 542454
rect 204187 542218 204229 542454
rect 203909 542134 204229 542218
rect 203909 541898 203951 542134
rect 204187 541898 204229 542134
rect 203909 541876 204229 541898
rect 206875 524454 207195 524476
rect 206875 524218 206917 524454
rect 207153 524218 207195 524454
rect 206875 524134 207195 524218
rect 206875 523898 206917 524134
rect 207153 523898 207195 524134
rect 206875 523876 207195 523898
rect 202404 492054 203004 519800
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 409022 203004 419498
rect 206004 495654 206604 519800
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 409022 206604 423098
rect 209604 499254 210204 519800
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 409022 210204 426698
rect 216804 506454 217404 519800
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 409022 217404 433898
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 409022 221004 437498
rect 224004 693654 224604 708042
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 549654 224604 585098
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 409022 224604 441098
rect 227604 697254 228204 709922
rect 245604 711418 246204 711440
rect 245604 711182 245786 711418
rect 246022 711182 246204 711418
rect 245604 711098 246204 711182
rect 245604 710862 245786 711098
rect 246022 710862 246204 711098
rect 242004 709538 242604 709560
rect 242004 709302 242186 709538
rect 242422 709302 242604 709538
rect 242004 709218 242604 709302
rect 242004 708982 242186 709218
rect 242422 708982 242604 709218
rect 238404 707658 239004 707680
rect 238404 707422 238586 707658
rect 238822 707422 239004 707658
rect 238404 707338 239004 707422
rect 238404 707102 238586 707338
rect 238822 707102 239004 707338
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 553254 228204 588698
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 409022 228204 444698
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 234804 409022 235404 415898
rect 238404 672054 239004 707102
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 564054 239004 599498
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 420054 239004 455498
rect 238404 419818 238586 420054
rect 238822 419818 239004 420054
rect 238404 419734 239004 419818
rect 238404 419498 238586 419734
rect 238822 419498 239004 419734
rect 238404 409022 239004 419498
rect 242004 675654 242604 708982
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 567654 242604 603098
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 242004 495654 242604 531098
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 242004 423654 242604 459098
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 242004 409022 242604 423098
rect 245604 679254 246204 710862
rect 263604 710478 264204 711440
rect 263604 710242 263786 710478
rect 264022 710242 264204 710478
rect 263604 710158 264204 710242
rect 263604 709922 263786 710158
rect 264022 709922 264204 710158
rect 260004 708598 260604 709560
rect 260004 708362 260186 708598
rect 260422 708362 260604 708598
rect 260004 708278 260604 708362
rect 260004 708042 260186 708278
rect 260422 708042 260604 708278
rect 256404 706718 257004 707680
rect 256404 706482 256586 706718
rect 256822 706482 257004 706718
rect 256404 706398 257004 706482
rect 256404 706162 256586 706398
rect 256822 706162 257004 706398
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 571254 246204 606698
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 535254 246204 570698
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 245604 499254 246204 534698
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 245604 427254 246204 462698
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 245604 409022 246204 426698
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 252804 409022 253404 433898
rect 256404 690054 257004 706162
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 409022 257004 437498
rect 260004 693654 260604 708042
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 477654 260604 513098
rect 260004 477418 260186 477654
rect 260422 477418 260604 477654
rect 260004 477334 260604 477418
rect 260004 477098 260186 477334
rect 260422 477098 260604 477334
rect 260004 441654 260604 477098
rect 260004 441418 260186 441654
rect 260422 441418 260604 441654
rect 260004 441334 260604 441418
rect 260004 441098 260186 441334
rect 260422 441098 260604 441334
rect 260004 409022 260604 441098
rect 263604 697254 264204 709922
rect 281604 711418 282204 711440
rect 281604 711182 281786 711418
rect 282022 711182 282204 711418
rect 281604 711098 282204 711182
rect 281604 710862 281786 711098
rect 282022 710862 282204 711098
rect 278004 709538 278604 709560
rect 278004 709302 278186 709538
rect 278422 709302 278604 709538
rect 278004 709218 278604 709302
rect 278004 708982 278186 709218
rect 278422 708982 278604 709218
rect 274404 707658 275004 707680
rect 274404 707422 274586 707658
rect 274822 707422 275004 707658
rect 274404 707338 275004 707422
rect 274404 707102 274586 707338
rect 274822 707102 275004 707338
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 517254 264204 552698
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 481254 264204 516698
rect 263604 481018 263786 481254
rect 264022 481018 264204 481254
rect 263604 480934 264204 481018
rect 263604 480698 263786 480934
rect 264022 480698 264204 480934
rect 263604 445254 264204 480698
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 409022 264204 444698
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 266859 410412 266925 410413
rect 266859 410348 266860 410412
rect 266924 410348 266925 410412
rect 266859 410347 266925 410348
rect 204208 398454 204528 398476
rect 204208 398218 204250 398454
rect 204486 398218 204528 398454
rect 204208 398134 204528 398218
rect 204208 397898 204250 398134
rect 204486 397898 204528 398134
rect 204208 397876 204528 397898
rect 219568 380454 219888 380476
rect 219568 380218 219610 380454
rect 219846 380218 219888 380454
rect 219568 380134 219888 380218
rect 219568 379898 219610 380134
rect 219846 379898 219888 380134
rect 219568 379876 219888 379898
rect 204208 362454 204528 362476
rect 204208 362218 204250 362454
rect 204486 362218 204528 362454
rect 204208 362134 204528 362218
rect 204208 361898 204250 362134
rect 204486 361898 204528 362134
rect 204208 361876 204528 361898
rect 219568 344454 219888 344476
rect 219568 344218 219610 344454
rect 219846 344218 219888 344454
rect 219568 344134 219888 344218
rect 219568 343898 219610 344134
rect 219846 343898 219888 344134
rect 219568 343876 219888 343898
rect 202404 312054 203004 339800
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 199699 202060 199765 202061
rect 199699 201996 199700 202060
rect 199764 201996 199765 202060
rect 199699 201995 199765 201996
rect 202404 200200 203004 203498
rect 206004 315654 206604 339800
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 200200 206604 207098
rect 209604 319254 210204 339800
rect 209604 319018 209786 319254
rect 210022 319018 210204 319254
rect 209604 318934 210204 319018
rect 209604 318698 209786 318934
rect 210022 318698 210204 318934
rect 209604 283254 210204 318698
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 200200 210204 210698
rect 216804 326454 217404 339800
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 200200 217404 217898
rect 220404 330054 221004 339800
rect 220404 329818 220586 330054
rect 220822 329818 221004 330054
rect 220404 329734 221004 329818
rect 220404 329498 220586 329734
rect 220822 329498 221004 329734
rect 220404 294054 221004 329498
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 200200 221004 221498
rect 224004 333654 224604 339800
rect 224004 333418 224186 333654
rect 224422 333418 224604 333654
rect 224004 333334 224604 333418
rect 224004 333098 224186 333334
rect 224422 333098 224604 333334
rect 224004 297654 224604 333098
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 200200 224604 225098
rect 227604 337254 228204 339800
rect 227604 337018 227786 337254
rect 228022 337018 228204 337254
rect 227604 336934 228204 337018
rect 227604 336698 227786 336934
rect 228022 336698 228204 336934
rect 227604 301254 228204 336698
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 200200 228204 228698
rect 234804 308454 235404 339800
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200200 235404 235898
rect 238404 312054 239004 339800
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 200200 239004 203498
rect 242004 315654 242604 339800
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 200200 242604 207098
rect 245604 319254 246204 339800
rect 245604 319018 245786 319254
rect 246022 319018 246204 319254
rect 245604 318934 246204 319018
rect 245604 318698 245786 318934
rect 246022 318698 246204 318934
rect 245604 283254 246204 318698
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 200200 246204 210698
rect 252804 326454 253404 339800
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 200200 253404 217898
rect 256404 330054 257004 339800
rect 256404 329818 256586 330054
rect 256822 329818 257004 330054
rect 256404 329734 257004 329818
rect 256404 329498 256586 329734
rect 256822 329498 257004 329734
rect 256404 294054 257004 329498
rect 260004 333654 260604 339800
rect 260004 333418 260186 333654
rect 260422 333418 260604 333654
rect 260004 333334 260604 333418
rect 260004 333098 260186 333334
rect 260422 333098 260604 333334
rect 257659 317388 257725 317389
rect 257659 317324 257660 317388
rect 257724 317324 257725 317388
rect 257659 317323 257725 317324
rect 257662 311813 257722 317323
rect 257659 311812 257725 311813
rect 257659 311748 257660 311812
rect 257724 311748 257725 311812
rect 257659 311747 257725 311748
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 200200 257004 221498
rect 260004 297654 260604 333098
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 200200 260604 225098
rect 263604 337254 264204 339800
rect 263604 337018 263786 337254
rect 264022 337018 264204 337254
rect 263604 336934 264204 337018
rect 263604 336698 263786 336934
rect 264022 336698 264204 336934
rect 263604 301254 264204 336698
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 200200 264204 228698
rect 266862 201517 266922 410347
rect 267963 410276 268029 410277
rect 267963 410212 267964 410276
rect 268028 410212 268029 410276
rect 267963 410211 268029 410212
rect 267779 410140 267845 410141
rect 267779 410076 267780 410140
rect 267844 410076 267845 410140
rect 267779 410075 267845 410076
rect 267782 201653 267842 410075
rect 267966 202197 268026 410211
rect 268147 410004 268213 410005
rect 268147 409940 268148 410004
rect 268212 409940 268213 410004
rect 268147 409939 268213 409940
rect 268150 338741 268210 409939
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 344454 271404 379898
rect 270804 344218 270986 344454
rect 271222 344218 271404 344454
rect 270804 344134 271404 344218
rect 270804 343898 270986 344134
rect 271222 343898 271404 344134
rect 268147 338740 268213 338741
rect 268147 338676 268148 338740
rect 268212 338676 268213 338740
rect 268147 338675 268213 338676
rect 270804 308454 271404 343898
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 267963 202196 268029 202197
rect 267963 202132 267964 202196
rect 268028 202132 268029 202196
rect 267963 202131 268029 202132
rect 267779 201652 267845 201653
rect 267779 201588 267780 201652
rect 267844 201588 267845 201652
rect 267779 201587 267845 201588
rect 266859 201516 266925 201517
rect 266859 201452 266860 201516
rect 266924 201452 266925 201516
rect 266859 201451 266925 201452
rect 270804 200200 271404 235898
rect 274404 672054 275004 707102
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 420054 275004 455498
rect 274404 419818 274586 420054
rect 274822 419818 275004 420054
rect 274404 419734 275004 419818
rect 274404 419498 274586 419734
rect 274822 419498 275004 419734
rect 274404 384054 275004 419498
rect 274404 383818 274586 384054
rect 274822 383818 275004 384054
rect 274404 383734 275004 383818
rect 274404 383498 274586 383734
rect 274822 383498 275004 383734
rect 274404 348054 275004 383498
rect 274404 347818 274586 348054
rect 274822 347818 275004 348054
rect 274404 347734 275004 347818
rect 274404 347498 274586 347734
rect 274822 347498 275004 347734
rect 274404 312054 275004 347498
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 200200 275004 203498
rect 278004 675654 278604 708982
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 459654 278604 495098
rect 278004 459418 278186 459654
rect 278422 459418 278604 459654
rect 278004 459334 278604 459418
rect 278004 459098 278186 459334
rect 278422 459098 278604 459334
rect 278004 423654 278604 459098
rect 278004 423418 278186 423654
rect 278422 423418 278604 423654
rect 278004 423334 278604 423418
rect 278004 423098 278186 423334
rect 278422 423098 278604 423334
rect 278004 387654 278604 423098
rect 278004 387418 278186 387654
rect 278422 387418 278604 387654
rect 278004 387334 278604 387418
rect 278004 387098 278186 387334
rect 278422 387098 278604 387334
rect 278004 351654 278604 387098
rect 278004 351418 278186 351654
rect 278422 351418 278604 351654
rect 278004 351334 278604 351418
rect 278004 351098 278186 351334
rect 278422 351098 278604 351334
rect 278004 315654 278604 351098
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 200200 278604 207098
rect 281604 679254 282204 710862
rect 299604 710478 300204 711440
rect 299604 710242 299786 710478
rect 300022 710242 300204 710478
rect 299604 710158 300204 710242
rect 299604 709922 299786 710158
rect 300022 709922 300204 710158
rect 296004 708598 296604 709560
rect 296004 708362 296186 708598
rect 296422 708362 296604 708598
rect 296004 708278 296604 708362
rect 296004 708042 296186 708278
rect 296422 708042 296604 708278
rect 292404 706718 293004 707680
rect 292404 706482 292586 706718
rect 292822 706482 293004 706718
rect 292404 706398 293004 706482
rect 292404 706162 292586 706398
rect 292822 706162 293004 706398
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 463254 282204 498698
rect 281604 463018 281786 463254
rect 282022 463018 282204 463254
rect 281604 462934 282204 463018
rect 281604 462698 281786 462934
rect 282022 462698 282204 462934
rect 281604 427254 282204 462698
rect 281604 427018 281786 427254
rect 282022 427018 282204 427254
rect 281604 426934 282204 427018
rect 281604 426698 281786 426934
rect 282022 426698 282204 426934
rect 281604 391254 282204 426698
rect 281604 391018 281786 391254
rect 282022 391018 282204 391254
rect 281604 390934 282204 391018
rect 281604 390698 281786 390934
rect 282022 390698 282204 390934
rect 281604 355254 282204 390698
rect 281604 355018 281786 355254
rect 282022 355018 282204 355254
rect 281604 354934 282204 355018
rect 281604 354698 281786 354934
rect 282022 354698 282204 354934
rect 281604 319254 282204 354698
rect 281604 319018 281786 319254
rect 282022 319018 282204 319254
rect 281604 318934 282204 319018
rect 281604 318698 281786 318934
rect 282022 318698 282204 318934
rect 281604 283254 282204 318698
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 200200 282204 210698
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 200200 289404 217898
rect 292404 690054 293004 706162
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 200200 293004 221498
rect 296004 693654 296604 708042
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 299604 697254 300204 709922
rect 317604 711418 318204 711440
rect 317604 711182 317786 711418
rect 318022 711182 318204 711418
rect 317604 711098 318204 711182
rect 317604 710862 317786 711098
rect 318022 710862 318204 711098
rect 314004 709538 314604 709560
rect 314004 709302 314186 709538
rect 314422 709302 314604 709538
rect 314004 709218 314604 709302
rect 314004 708982 314186 709218
rect 314422 708982 314604 709218
rect 310404 707658 311004 707680
rect 310404 707422 310586 707658
rect 310822 707422 311004 707658
rect 310404 707338 311004 707422
rect 310404 707102 310586 707338
rect 310822 707102 311004 707338
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 580211 300204 588698
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 580211 307404 595898
rect 310404 672054 311004 707102
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 580211 311004 599498
rect 314004 675654 314604 708982
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 580211 314604 603098
rect 317604 679254 318204 710862
rect 335604 710478 336204 711440
rect 335604 710242 335786 710478
rect 336022 710242 336204 710478
rect 335604 710158 336204 710242
rect 335604 709922 335786 710158
rect 336022 709922 336204 710158
rect 332004 708598 332604 709560
rect 332004 708362 332186 708598
rect 332422 708362 332604 708598
rect 332004 708278 332604 708362
rect 332004 708042 332186 708278
rect 332422 708042 332604 708278
rect 328404 706718 329004 707680
rect 328404 706482 328586 706718
rect 328822 706482 329004 706718
rect 328404 706398 329004 706482
rect 328404 706162 328586 706398
rect 328822 706162 329004 706398
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 580211 318204 606698
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 580211 325404 613898
rect 328404 690054 329004 706162
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 580211 329004 581498
rect 332004 693654 332604 708042
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 580211 332604 585098
rect 335604 697254 336204 709922
rect 353604 711418 354204 711440
rect 353604 711182 353786 711418
rect 354022 711182 354204 711418
rect 353604 711098 354204 711182
rect 353604 710862 353786 711098
rect 354022 710862 354204 711098
rect 350004 709538 350604 709560
rect 350004 709302 350186 709538
rect 350422 709302 350604 709538
rect 350004 709218 350604 709302
rect 350004 708982 350186 709218
rect 350422 708982 350604 709218
rect 346404 707658 347004 707680
rect 346404 707422 346586 707658
rect 346822 707422 347004 707658
rect 346404 707338 347004 707422
rect 346404 707102 346586 707338
rect 346822 707102 347004 707338
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 580211 336204 588698
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 580211 343404 595898
rect 346404 672054 347004 707102
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 580211 347004 599498
rect 350004 675654 350604 708982
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 580211 350604 603098
rect 353604 679254 354204 710862
rect 371604 710478 372204 711440
rect 371604 710242 371786 710478
rect 372022 710242 372204 710478
rect 371604 710158 372204 710242
rect 371604 709922 371786 710158
rect 372022 709922 372204 710158
rect 368004 708598 368604 709560
rect 368004 708362 368186 708598
rect 368422 708362 368604 708598
rect 368004 708278 368604 708362
rect 368004 708042 368186 708278
rect 368422 708042 368604 708278
rect 364404 706718 365004 707680
rect 364404 706482 364586 706718
rect 364822 706482 365004 706718
rect 364404 706398 365004 706482
rect 364404 706162 364586 706398
rect 364822 706162 365004 706398
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 580211 354204 606698
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 580211 361404 613898
rect 364404 690054 365004 706162
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 580211 365004 581498
rect 368004 693654 368604 708042
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 580211 368604 585098
rect 371604 697254 372204 709922
rect 389604 711418 390204 711440
rect 389604 711182 389786 711418
rect 390022 711182 390204 711418
rect 389604 711098 390204 711182
rect 389604 710862 389786 711098
rect 390022 710862 390204 711098
rect 386004 709538 386604 709560
rect 386004 709302 386186 709538
rect 386422 709302 386604 709538
rect 386004 709218 386604 709302
rect 386004 708982 386186 709218
rect 386422 708982 386604 709218
rect 382404 707658 383004 707680
rect 382404 707422 382586 707658
rect 382822 707422 383004 707658
rect 382404 707338 383004 707422
rect 382404 707102 382586 707338
rect 382822 707102 383004 707338
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 580211 372204 588698
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 319568 560454 319888 560476
rect 319568 560218 319610 560454
rect 319846 560218 319888 560454
rect 319568 560134 319888 560218
rect 319568 559898 319610 560134
rect 319846 559898 319888 560134
rect 319568 559876 319888 559898
rect 378804 560454 379404 595898
rect 382404 672054 383004 707102
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 379467 572116 379533 572117
rect 379467 572052 379468 572116
rect 379532 572052 379533 572116
rect 379467 572051 379533 572052
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 304208 542454 304528 542476
rect 304208 542218 304250 542454
rect 304486 542218 304528 542454
rect 304208 542134 304528 542218
rect 304208 541898 304250 542134
rect 304486 541898 304528 542134
rect 304208 541876 304528 541898
rect 319568 524454 319888 524476
rect 319568 524218 319610 524454
rect 319846 524218 319888 524454
rect 319568 524134 319888 524218
rect 319568 523898 319610 524134
rect 319846 523898 319888 524134
rect 319568 523876 319888 523898
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 304208 506454 304528 506476
rect 304208 506218 304250 506454
rect 304486 506218 304528 506454
rect 304208 506134 304528 506218
rect 304208 505898 304250 506134
rect 304486 505898 304528 506134
rect 304208 505876 304528 505898
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 200200 296604 225098
rect 299604 481254 300204 499800
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299604 301254 300204 336698
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 200200 300204 228698
rect 306804 488454 307404 499800
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200200 307404 235898
rect 310404 492054 311004 499800
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 200200 311004 203498
rect 314004 495654 314604 499800
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 200200 314604 207098
rect 317604 499254 318204 499800
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 200200 318204 210698
rect 324804 470454 325404 499800
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 200200 325404 217898
rect 328404 474054 329004 499800
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 294054 329004 329498
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 200200 329004 221498
rect 332004 477654 332604 499800
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 297654 332604 333098
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 200200 332604 225098
rect 335604 481254 336204 499800
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 335604 301254 336204 336698
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 200200 336204 228698
rect 342804 488454 343404 499800
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200200 343404 235898
rect 346404 492054 347004 499800
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 384054 347004 419498
rect 346404 383818 346586 384054
rect 346822 383818 347004 384054
rect 346404 383734 347004 383818
rect 346404 383498 346586 383734
rect 346822 383498 347004 383734
rect 346404 348054 347004 383498
rect 346404 347818 346586 348054
rect 346822 347818 347004 348054
rect 346404 347734 347004 347818
rect 346404 347498 346586 347734
rect 346822 347498 347004 347734
rect 346404 312054 347004 347498
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 200200 347004 203498
rect 350004 495654 350604 499800
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 387654 350604 423098
rect 350004 387418 350186 387654
rect 350422 387418 350604 387654
rect 350004 387334 350604 387418
rect 350004 387098 350186 387334
rect 350422 387098 350604 387334
rect 350004 351654 350604 387098
rect 350004 351418 350186 351654
rect 350422 351418 350604 351654
rect 350004 351334 350604 351418
rect 350004 351098 350186 351334
rect 350422 351098 350604 351334
rect 350004 315654 350604 351098
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 200200 350604 207098
rect 353604 499254 354204 499800
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 391254 354204 426698
rect 353604 391018 353786 391254
rect 354022 391018 354204 391254
rect 353604 390934 354204 391018
rect 353604 390698 353786 390934
rect 354022 390698 354204 390934
rect 353604 355254 354204 390698
rect 353604 355018 353786 355254
rect 354022 355018 354204 355254
rect 353604 354934 354204 355018
rect 353604 354698 353786 354934
rect 354022 354698 354204 354934
rect 353604 319254 354204 354698
rect 353604 319018 353786 319254
rect 354022 319018 354204 319254
rect 353604 318934 354204 319018
rect 353604 318698 353786 318934
rect 354022 318698 354204 318934
rect 353604 283254 354204 318698
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 200200 354204 210698
rect 360804 470454 361404 499800
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 200200 361404 217898
rect 364404 474054 365004 499800
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 402054 365004 437498
rect 364404 401818 364586 402054
rect 364822 401818 365004 402054
rect 364404 401734 365004 401818
rect 364404 401498 364586 401734
rect 364822 401498 365004 401734
rect 364404 366054 365004 401498
rect 364404 365818 364586 366054
rect 364822 365818 365004 366054
rect 364404 365734 365004 365818
rect 364404 365498 364586 365734
rect 364822 365498 365004 365734
rect 364404 330054 365004 365498
rect 364404 329818 364586 330054
rect 364822 329818 365004 330054
rect 364404 329734 365004 329818
rect 364404 329498 364586 329734
rect 364822 329498 365004 329734
rect 364404 294054 365004 329498
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 200200 365004 221498
rect 368004 477654 368604 499800
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 405654 368604 441098
rect 368004 405418 368186 405654
rect 368422 405418 368604 405654
rect 368004 405334 368604 405418
rect 368004 405098 368186 405334
rect 368422 405098 368604 405334
rect 368004 369654 368604 405098
rect 368004 369418 368186 369654
rect 368422 369418 368604 369654
rect 368004 369334 368604 369418
rect 368004 369098 368186 369334
rect 368422 369098 368604 369334
rect 368004 333654 368604 369098
rect 368004 333418 368186 333654
rect 368422 333418 368604 333654
rect 368004 333334 368604 333418
rect 368004 333098 368186 333334
rect 368422 333098 368604 333334
rect 368004 297654 368604 333098
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 200200 368604 225098
rect 371604 481254 372204 499800
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 409254 372204 444698
rect 371604 409018 371786 409254
rect 372022 409018 372204 409254
rect 371604 408934 372204 409018
rect 371604 408698 371786 408934
rect 372022 408698 372204 408934
rect 371604 373254 372204 408698
rect 371604 373018 371786 373254
rect 372022 373018 372204 373254
rect 371604 372934 372204 373018
rect 371604 372698 371786 372934
rect 372022 372698 372204 372934
rect 371604 337254 372204 372698
rect 371604 337018 371786 337254
rect 372022 337018 372204 337254
rect 371604 336934 372204 337018
rect 371604 336698 371786 336934
rect 372022 336698 372204 336934
rect 371604 301254 372204 336698
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 200200 372204 228698
rect 378804 488454 379404 523898
rect 379470 500309 379530 572051
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 379651 541108 379717 541109
rect 379651 541044 379652 541108
rect 379716 541044 379717 541108
rect 379651 541043 379717 541044
rect 379467 500308 379533 500309
rect 379467 500244 379468 500308
rect 379532 500244 379533 500308
rect 379467 500243 379533 500244
rect 379654 500173 379714 541043
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 379651 500172 379717 500173
rect 379651 500108 379652 500172
rect 379716 500108 379717 500172
rect 379651 500107 379717 500108
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200200 379404 235898
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 382404 384054 383004 419498
rect 382404 383818 382586 384054
rect 382822 383818 383004 384054
rect 382404 383734 383004 383818
rect 382404 383498 382586 383734
rect 382822 383498 383004 383734
rect 386004 675654 386604 708982
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 387654 386604 423098
rect 386004 387418 386186 387654
rect 386422 387418 386604 387654
rect 386004 387334 386604 387418
rect 386004 387098 386186 387334
rect 386422 387098 386604 387334
rect 386004 383619 386604 387098
rect 389604 679254 390204 710862
rect 407604 710478 408204 711440
rect 407604 710242 407786 710478
rect 408022 710242 408204 710478
rect 407604 710158 408204 710242
rect 407604 709922 407786 710158
rect 408022 709922 408204 710158
rect 404004 708598 404604 709560
rect 404004 708362 404186 708598
rect 404422 708362 404604 708598
rect 404004 708278 404604 708362
rect 404004 708042 404186 708278
rect 404422 708042 404604 708278
rect 400404 706718 401004 707680
rect 400404 706482 400586 706718
rect 400822 706482 401004 706718
rect 400404 706398 401004 706482
rect 400404 706162 400586 706398
rect 400822 706162 401004 706398
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 391254 390204 426698
rect 389604 391018 389786 391254
rect 390022 391018 390204 391254
rect 389604 390934 390204 391018
rect 389604 390698 389786 390934
rect 390022 390698 390204 390934
rect 389604 383619 390204 390698
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 383619 397404 397898
rect 400404 690054 401004 706162
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 383619 401004 401498
rect 404004 693654 404604 708042
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 383619 404604 405098
rect 407604 697254 408204 709922
rect 425604 711418 426204 711440
rect 425604 711182 425786 711418
rect 426022 711182 426204 711418
rect 425604 711098 426204 711182
rect 425604 710862 425786 711098
rect 426022 710862 426204 711098
rect 422004 709538 422604 709560
rect 422004 709302 422186 709538
rect 422422 709302 422604 709538
rect 422004 709218 422604 709302
rect 422004 708982 422186 709218
rect 422422 708982 422604 709218
rect 418404 707658 419004 707680
rect 418404 707422 418586 707658
rect 418822 707422 419004 707658
rect 418404 707338 419004 707422
rect 418404 707102 418586 707338
rect 418822 707102 419004 707338
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 383619 408204 408698
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 383619 415404 415898
rect 418404 672054 419004 707102
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 382404 348054 383004 383498
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 394604 380454 394924 380476
rect 394604 380218 394646 380454
rect 394882 380218 394924 380454
rect 394604 380134 394924 380218
rect 394604 379898 394646 380134
rect 394882 379898 394924 380134
rect 394604 379876 394924 379898
rect 389774 362454 390094 362476
rect 389774 362218 389816 362454
rect 390052 362218 390094 362454
rect 389774 362134 390094 362218
rect 389774 361898 389816 362134
rect 390052 361898 390094 362134
rect 389774 361876 390094 361898
rect 382404 347818 382586 348054
rect 382822 347818 383004 348054
rect 382404 347734 383004 347818
rect 382404 347498 382586 347734
rect 382822 347498 383004 347734
rect 382404 312054 383004 347498
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 200200 383004 203498
rect 386004 315654 386604 349800
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 200200 386604 207098
rect 389604 319254 390204 349800
rect 389604 319018 389786 319254
rect 390022 319018 390204 319254
rect 389604 318934 390204 319018
rect 389604 318698 389786 318934
rect 390022 318698 390204 318934
rect 389604 283254 390204 318698
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 200200 390204 210698
rect 396804 326454 397404 349800
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 200200 397404 217898
rect 400404 330054 401004 349800
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 200200 401004 221498
rect 404004 333654 404604 349800
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 297654 404604 333098
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 200200 404604 225098
rect 407604 337254 408204 349800
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 301254 408204 336698
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 200200 408204 228698
rect 414804 344454 415404 349800
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200200 415404 235898
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 200200 419004 203498
rect 422004 675654 422604 708982
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 200200 422604 207098
rect 425604 679254 426204 710862
rect 443604 710478 444204 711440
rect 443604 710242 443786 710478
rect 444022 710242 444204 710478
rect 443604 710158 444204 710242
rect 443604 709922 443786 710158
rect 444022 709922 444204 710158
rect 440004 708598 440604 709560
rect 440004 708362 440186 708598
rect 440422 708362 440604 708598
rect 440004 708278 440604 708362
rect 440004 708042 440186 708278
rect 440422 708042 440604 708278
rect 436404 706718 437004 707680
rect 436404 706482 436586 706718
rect 436822 706482 437004 706718
rect 436404 706398 437004 706482
rect 436404 706162 436586 706398
rect 436822 706162 437004 706398
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 200200 426204 210698
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 200200 433404 217898
rect 436404 690054 437004 706162
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 138208 182454 138528 182476
rect 138208 182218 138250 182454
rect 138486 182218 138528 182454
rect 138208 182134 138528 182218
rect 138208 181898 138250 182134
rect 138486 181898 138528 182134
rect 138208 181876 138528 181898
rect 133643 175132 133709 175133
rect 133643 175068 133644 175132
rect 133708 175068 133709 175132
rect 133643 175067 133709 175068
rect 133459 174044 133525 174045
rect 133459 173980 133460 174044
rect 133524 173980 133525 174044
rect 133459 173979 133525 173980
rect 153568 164454 153888 164476
rect 153568 164218 153610 164454
rect 153846 164218 153888 164454
rect 153568 164134 153888 164218
rect 153568 163898 153610 164134
rect 153846 163898 153888 164134
rect 153568 163876 153888 163898
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 138208 146454 138528 146476
rect 138208 146218 138250 146454
rect 138486 146218 138528 146454
rect 138208 146134 138528 146218
rect 138208 145898 138250 146134
rect 138486 145898 138528 146134
rect 138208 145876 138528 145898
rect 133275 132972 133341 132973
rect 133275 132908 133276 132972
rect 133340 132908 133341 132972
rect 133275 132907 133341 132908
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 153568 128454 153888 128476
rect 153568 128218 153610 128454
rect 153846 128218 153888 128454
rect 153568 128134 153888 128218
rect 153568 127898 153610 128134
rect 153846 127898 153888 128134
rect 153568 127876 153888 127898
rect 133827 119780 133893 119781
rect 133827 119716 133828 119780
rect 133892 119716 133893 119780
rect 133827 119715 133893 119716
rect 133830 117877 133890 119715
rect 133827 117876 133893 117877
rect 133827 117812 133828 117876
rect 133892 117812 133893 117876
rect 133827 117811 133893 117812
rect 133827 117604 133893 117605
rect 133827 117540 133828 117604
rect 133892 117540 133893 117604
rect 133827 117539 133893 117540
rect 133830 117469 133890 117539
rect 133827 117468 133893 117469
rect 133827 117404 133828 117468
rect 133892 117404 133893 117468
rect 133827 117403 133893 117404
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3166 131004 23498
rect 130404 -3402 130586 -3166
rect 130822 -3402 131004 -3166
rect 130404 -3486 131004 -3402
rect 130404 -3722 130586 -3486
rect 130822 -3722 131004 -3486
rect 130404 -3744 131004 -3722
rect 134004 99654 134604 119800
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -5046 134604 27098
rect 134004 -5282 134186 -5046
rect 134422 -5282 134604 -5046
rect 134004 -5366 134604 -5282
rect 134004 -5602 134186 -5366
rect 134422 -5602 134604 -5366
rect 134004 -5624 134604 -5602
rect 137604 103254 138204 119800
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 144804 110454 145404 119800
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 140819 38588 140885 38589
rect 140819 38524 140820 38588
rect 140884 38524 140885 38588
rect 140819 38523 140885 38524
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6222 119786 -5986
rect 120022 -6222 120204 -5986
rect 119604 -6306 120204 -6222
rect 119604 -6542 119786 -6306
rect 120022 -6542 120204 -6306
rect 119604 -7504 120204 -6542
rect 137604 -6926 138204 30698
rect 140822 29069 140882 38523
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 140819 29068 140885 29069
rect 140819 29004 140820 29068
rect 140884 29004 140885 29068
rect 140819 29003 140885 29004
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 148404 114054 149004 119800
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2226 149004 5498
rect 148404 -2462 148586 -2226
rect 148822 -2462 149004 -2226
rect 148404 -2546 149004 -2462
rect 148404 -2782 148586 -2546
rect 148822 -2782 149004 -2546
rect 148404 -3744 149004 -2782
rect 152004 117654 152604 119800
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4106 152604 9098
rect 152004 -4342 152186 -4106
rect 152422 -4342 152604 -4106
rect 152004 -4426 152604 -4342
rect 152004 -4662 152186 -4426
rect 152422 -4662 152604 -4426
rect 152004 -5624 152604 -4662
rect 155604 85254 156204 119800
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 162804 92454 163404 119800
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 157379 70412 157445 70413
rect 157379 70348 157380 70412
rect 157444 70348 157445 70412
rect 157379 70347 157445 70348
rect 157382 66333 157442 70347
rect 157379 66332 157445 66333
rect 157379 66268 157380 66332
rect 157444 66268 157445 66332
rect 157379 66267 157445 66268
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7162 137786 -6926
rect 138022 -7162 138204 -6926
rect 137604 -7246 138204 -7162
rect 137604 -7482 137786 -7246
rect 138022 -7482 138204 -7246
rect 137604 -7504 138204 -7482
rect 155604 -5986 156204 12698
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 166404 96054 167004 119800
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3166 167004 23498
rect 166404 -3402 166586 -3166
rect 166822 -3402 167004 -3166
rect 166404 -3486 167004 -3402
rect 166404 -3722 166586 -3486
rect 166822 -3722 167004 -3486
rect 166404 -3744 167004 -3722
rect 170004 99654 170604 119800
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -5046 170604 27098
rect 170004 -5282 170186 -5046
rect 170422 -5282 170604 -5046
rect 170004 -5366 170604 -5282
rect 170004 -5602 170186 -5366
rect 170422 -5602 170604 -5366
rect 170004 -5624 170604 -5602
rect 173604 103254 174204 119800
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6222 155786 -5986
rect 156022 -6222 156204 -5986
rect 155604 -6306 156204 -6222
rect 155604 -6542 155786 -6306
rect 156022 -6542 156204 -6306
rect 155604 -7504 156204 -6542
rect 173604 -6926 174204 30698
rect 180804 110454 181404 119800
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 184404 114054 185004 119800
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2226 185004 5498
rect 184404 -2462 184586 -2226
rect 184822 -2462 185004 -2226
rect 184404 -2546 185004 -2462
rect 184404 -2782 184586 -2546
rect 184822 -2782 185004 -2546
rect 184404 -3744 185004 -2782
rect 188004 117654 188604 119800
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4106 188604 9098
rect 188004 -4342 188186 -4106
rect 188422 -4342 188604 -4106
rect 188004 -4426 188604 -4342
rect 188004 -4662 188186 -4426
rect 188422 -4662 188604 -4426
rect 188004 -5624 188604 -4662
rect 191604 85254 192204 119800
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7162 173786 -6926
rect 174022 -7162 174204 -6926
rect 173604 -7246 174204 -7162
rect 173604 -7482 173786 -7246
rect 174022 -7482 174204 -7246
rect 173604 -7504 174204 -7482
rect 191604 -5986 192204 12698
rect 198804 92454 199404 119800
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 202404 96054 203004 119800
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3166 203004 23498
rect 202404 -3402 202586 -3166
rect 202822 -3402 203004 -3166
rect 202404 -3486 203004 -3402
rect 202404 -3722 202586 -3486
rect 202822 -3722 203004 -3486
rect 202404 -3744 203004 -3722
rect 206004 99654 206604 119800
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -5046 206604 27098
rect 206004 -5282 206186 -5046
rect 206422 -5282 206604 -5046
rect 206004 -5366 206604 -5282
rect 206004 -5602 206186 -5366
rect 206422 -5602 206604 -5366
rect 206004 -5624 206604 -5602
rect 209604 103254 210204 119800
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6222 191786 -5986
rect 192022 -6222 192204 -5986
rect 191604 -6306 192204 -6222
rect 191604 -6542 191786 -6306
rect 192022 -6542 192204 -6306
rect 191604 -7504 192204 -6542
rect 209604 -6926 210204 30698
rect 216804 110454 217404 119800
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 220404 114054 221004 119800
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2226 221004 5498
rect 220404 -2462 220586 -2226
rect 220822 -2462 221004 -2226
rect 220404 -2546 221004 -2462
rect 220404 -2782 220586 -2546
rect 220822 -2782 221004 -2546
rect 220404 -3744 221004 -2782
rect 224004 117654 224604 119800
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4106 224604 9098
rect 224004 -4342 224186 -4106
rect 224422 -4342 224604 -4106
rect 224004 -4426 224604 -4342
rect 224004 -4662 224186 -4426
rect 224422 -4662 224604 -4426
rect 224004 -5624 224604 -4662
rect 227604 85254 228204 119800
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7162 209786 -6926
rect 210022 -7162 210204 -6926
rect 209604 -7246 210204 -7162
rect 209604 -7482 209786 -7246
rect 210022 -7482 210204 -7246
rect 209604 -7504 210204 -7482
rect 227604 -5986 228204 12698
rect 234804 92454 235404 119800
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 238404 96054 239004 119800
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3166 239004 23498
rect 238404 -3402 238586 -3166
rect 238822 -3402 239004 -3166
rect 238404 -3486 239004 -3402
rect 238404 -3722 238586 -3486
rect 238822 -3722 239004 -3486
rect 238404 -3744 239004 -3722
rect 242004 99654 242604 119800
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -5046 242604 27098
rect 242004 -5282 242186 -5046
rect 242422 -5282 242604 -5046
rect 242004 -5366 242604 -5282
rect 242004 -5602 242186 -5366
rect 242422 -5602 242604 -5366
rect 242004 -5624 242604 -5602
rect 245604 103254 246204 119800
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6222 227786 -5986
rect 228022 -6222 228204 -5986
rect 227604 -6306 228204 -6222
rect 227604 -6542 227786 -6306
rect 228022 -6542 228204 -6306
rect 227604 -7504 228204 -6542
rect 245604 -6926 246204 30698
rect 252804 110454 253404 119800
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 256404 114054 257004 119800
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2226 257004 5498
rect 256404 -2462 256586 -2226
rect 256822 -2462 257004 -2226
rect 256404 -2546 257004 -2462
rect 256404 -2782 256586 -2546
rect 256822 -2782 257004 -2546
rect 256404 -3744 257004 -2782
rect 260004 117654 260604 119800
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4106 260604 9098
rect 260004 -4342 260186 -4106
rect 260422 -4342 260604 -4106
rect 260004 -4426 260604 -4342
rect 260004 -4662 260186 -4426
rect 260422 -4662 260604 -4426
rect 260004 -5624 260604 -4662
rect 263604 85254 264204 119800
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7162 245786 -6926
rect 246022 -7162 246204 -6926
rect 245604 -7246 246204 -7162
rect 245604 -7482 245786 -7246
rect 246022 -7482 246204 -7246
rect 245604 -7504 246204 -7482
rect 263604 -5986 264204 12698
rect 270804 92454 271404 119800
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 274404 96054 275004 119800
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3166 275004 23498
rect 274404 -3402 274586 -3166
rect 274822 -3402 275004 -3166
rect 274404 -3486 275004 -3402
rect 274404 -3722 274586 -3486
rect 274822 -3722 275004 -3486
rect 274404 -3744 275004 -3722
rect 278004 99654 278604 119800
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -5046 278604 27098
rect 278004 -5282 278186 -5046
rect 278422 -5282 278604 -5046
rect 278004 -5366 278604 -5282
rect 278004 -5602 278186 -5366
rect 278422 -5602 278604 -5366
rect 278004 -5624 278604 -5602
rect 281604 103254 282204 119800
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6222 263786 -5986
rect 264022 -6222 264204 -5986
rect 263604 -6306 264204 -6222
rect 263604 -6542 263786 -6306
rect 264022 -6542 264204 -6306
rect 263604 -7504 264204 -6542
rect 281604 -6926 282204 30698
rect 288804 110454 289404 119800
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 292404 114054 293004 119800
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 290595 99516 290661 99517
rect 290595 99452 290596 99516
rect 290660 99452 290661 99516
rect 290595 99451 290661 99452
rect 290598 96661 290658 99451
rect 290595 96660 290661 96661
rect 290595 96596 290596 96660
rect 290660 96596 290661 96660
rect 290595 96595 290661 96596
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 290411 67692 290477 67693
rect 290411 67628 290412 67692
rect 290476 67628 290477 67692
rect 290411 67627 290477 67628
rect 290414 66333 290474 67627
rect 290411 66332 290477 66333
rect 290411 66268 290412 66332
rect 290476 66268 290477 66332
rect 290411 66267 290477 66268
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2226 293004 5498
rect 292404 -2462 292586 -2226
rect 292822 -2462 293004 -2226
rect 292404 -2546 293004 -2462
rect 292404 -2782 292586 -2546
rect 292822 -2782 293004 -2546
rect 292404 -3744 293004 -2782
rect 296004 117654 296604 119800
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4106 296604 9098
rect 296004 -4342 296186 -4106
rect 296422 -4342 296604 -4106
rect 296004 -4426 296604 -4342
rect 296004 -4662 296186 -4426
rect 296422 -4662 296604 -4426
rect 296004 -5624 296604 -4662
rect 299604 85254 300204 119800
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7162 281786 -6926
rect 282022 -7162 282204 -6926
rect 281604 -7246 282204 -7162
rect 281604 -7482 281786 -7246
rect 282022 -7482 282204 -7246
rect 281604 -7504 282204 -7482
rect 299604 -5986 300204 12698
rect 306804 92454 307404 119800
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 310404 96054 311004 119800
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3166 311004 23498
rect 310404 -3402 310586 -3166
rect 310822 -3402 311004 -3166
rect 310404 -3486 311004 -3402
rect 310404 -3722 310586 -3486
rect 310822 -3722 311004 -3486
rect 310404 -3744 311004 -3722
rect 314004 99654 314604 119800
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -5046 314604 27098
rect 314004 -5282 314186 -5046
rect 314422 -5282 314604 -5046
rect 314004 -5366 314604 -5282
rect 314004 -5602 314186 -5366
rect 314422 -5602 314604 -5366
rect 314004 -5624 314604 -5602
rect 317604 103254 318204 119800
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6222 299786 -5986
rect 300022 -6222 300204 -5986
rect 299604 -6306 300204 -6222
rect 299604 -6542 299786 -6306
rect 300022 -6542 300204 -6306
rect 299604 -7504 300204 -6542
rect 317604 -6926 318204 30698
rect 324804 110454 325404 119800
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 328404 114054 329004 119800
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2226 329004 5498
rect 328404 -2462 328586 -2226
rect 328822 -2462 329004 -2226
rect 328404 -2546 329004 -2462
rect 328404 -2782 328586 -2546
rect 328822 -2782 329004 -2546
rect 328404 -3744 329004 -2782
rect 332004 117654 332604 119800
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4106 332604 9098
rect 332004 -4342 332186 -4106
rect 332422 -4342 332604 -4106
rect 332004 -4426 332604 -4342
rect 332004 -4662 332186 -4426
rect 332422 -4662 332604 -4426
rect 332004 -5624 332604 -4662
rect 335604 85254 336204 119800
rect 341379 99516 341445 99517
rect 341379 99452 341380 99516
rect 341444 99452 341445 99516
rect 341379 99451 341445 99452
rect 341382 96661 341442 99451
rect 341379 96660 341445 96661
rect 341379 96596 341380 96660
rect 341444 96596 341445 96660
rect 341379 96595 341445 96596
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7162 317786 -6926
rect 318022 -7162 318204 -6926
rect 317604 -7246 318204 -7162
rect 317604 -7482 317786 -7246
rect 318022 -7482 318204 -7246
rect 317604 -7504 318204 -7482
rect 335604 -5986 336204 12698
rect 342804 92454 343404 119800
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 346404 96054 347004 119800
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3166 347004 23498
rect 346404 -3402 346586 -3166
rect 346822 -3402 347004 -3166
rect 346404 -3486 347004 -3402
rect 346404 -3722 346586 -3486
rect 346822 -3722 347004 -3486
rect 346404 -3744 347004 -3722
rect 350004 99654 350604 119800
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -5046 350604 27098
rect 350004 -5282 350186 -5046
rect 350422 -5282 350604 -5046
rect 350004 -5366 350604 -5282
rect 350004 -5602 350186 -5366
rect 350422 -5602 350604 -5366
rect 350004 -5624 350604 -5602
rect 353604 103254 354204 119800
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6222 335786 -5986
rect 336022 -6222 336204 -5986
rect 335604 -6306 336204 -6222
rect 335604 -6542 335786 -6306
rect 336022 -6542 336204 -6306
rect 335604 -7504 336204 -6542
rect 353604 -6926 354204 30698
rect 360804 110454 361404 119800
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 364404 114054 365004 119800
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2226 365004 5498
rect 364404 -2462 364586 -2226
rect 364822 -2462 365004 -2226
rect 364404 -2546 365004 -2462
rect 364404 -2782 364586 -2546
rect 364822 -2782 365004 -2546
rect 364404 -3744 365004 -2782
rect 368004 117654 368604 119800
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4106 368604 9098
rect 368004 -4342 368186 -4106
rect 368422 -4342 368604 -4106
rect 368004 -4426 368604 -4342
rect 368004 -4662 368186 -4426
rect 368422 -4662 368604 -4426
rect 368004 -5624 368604 -4662
rect 371604 85254 372204 119800
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7162 353786 -6926
rect 354022 -7162 354204 -6926
rect 353604 -7246 354204 -7162
rect 353604 -7482 353786 -7246
rect 354022 -7482 354204 -7246
rect 353604 -7504 354204 -7482
rect 371604 -5986 372204 12698
rect 378804 92454 379404 119800
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 382404 96054 383004 119800
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3166 383004 23498
rect 382404 -3402 382586 -3166
rect 382822 -3402 383004 -3166
rect 382404 -3486 383004 -3402
rect 382404 -3722 382586 -3486
rect 382822 -3722 383004 -3486
rect 382404 -3744 383004 -3722
rect 386004 99654 386604 119800
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -5046 386604 27098
rect 386004 -5282 386186 -5046
rect 386422 -5282 386604 -5046
rect 386004 -5366 386604 -5282
rect 386004 -5602 386186 -5366
rect 386422 -5602 386604 -5366
rect 386004 -5624 386604 -5602
rect 389604 103254 390204 119800
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6222 371786 -5986
rect 372022 -6222 372204 -5986
rect 371604 -6306 372204 -6222
rect 371604 -6542 371786 -6306
rect 372022 -6542 372204 -6306
rect 371604 -7504 372204 -6542
rect 389604 -6926 390204 30698
rect 396804 110454 397404 119800
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 400404 114054 401004 119800
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2226 401004 5498
rect 400404 -2462 400586 -2226
rect 400822 -2462 401004 -2226
rect 400404 -2546 401004 -2462
rect 400404 -2782 400586 -2546
rect 400822 -2782 401004 -2546
rect 400404 -3744 401004 -2782
rect 404004 117654 404604 119800
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4106 404604 9098
rect 404004 -4342 404186 -4106
rect 404422 -4342 404604 -4106
rect 404004 -4426 404604 -4342
rect 404004 -4662 404186 -4426
rect 404422 -4662 404604 -4426
rect 404004 -5624 404604 -4662
rect 407604 85254 408204 119800
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7162 389786 -6926
rect 390022 -7162 390204 -6926
rect 389604 -7246 390204 -7162
rect 389604 -7482 389786 -7246
rect 390022 -7482 390204 -7246
rect 389604 -7504 390204 -7482
rect 407604 -5986 408204 12698
rect 414804 92454 415404 119800
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 418404 96054 419004 119800
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 422004 99654 422604 119800
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 420683 61436 420749 61437
rect 420683 61372 420684 61436
rect 420748 61372 420749 61436
rect 420683 61371 420749 61372
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 420686 48381 420746 61371
rect 420683 48380 420749 48381
rect 420683 48316 420684 48380
rect 420748 48316 420749 48380
rect 420683 48315 420749 48316
rect 420683 42124 420749 42125
rect 420683 42060 420684 42124
rect 420748 42060 420749 42124
rect 420683 42059 420749 42060
rect 420686 29069 420746 42059
rect 420683 29068 420749 29069
rect 420683 29004 420684 29068
rect 420748 29004 420749 29068
rect 420683 29003 420749 29004
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3166 419004 23498
rect 418404 -3402 418586 -3166
rect 418822 -3402 419004 -3166
rect 418404 -3486 419004 -3402
rect 418404 -3722 418586 -3486
rect 418822 -3722 419004 -3486
rect 418404 -3744 419004 -3722
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -5046 422604 27098
rect 422004 -5282 422186 -5046
rect 422422 -5282 422604 -5046
rect 422004 -5366 422604 -5282
rect 422004 -5602 422186 -5366
rect 422422 -5602 422604 -5366
rect 422004 -5624 422604 -5602
rect 425604 103254 426204 119800
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6222 407786 -5986
rect 408022 -6222 408204 -5986
rect 407604 -6306 408204 -6222
rect 407604 -6542 407786 -6306
rect 408022 -6542 408204 -6306
rect 407604 -7504 408204 -6542
rect 425604 -6926 426204 30698
rect 432804 110454 433404 119800
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2226 437004 5498
rect 436404 -2462 436586 -2226
rect 436822 -2462 437004 -2226
rect 436404 -2546 437004 -2462
rect 436404 -2782 436586 -2546
rect 436822 -2782 437004 -2546
rect 436404 -3744 437004 -2782
rect 440004 693654 440604 708042
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4106 440604 9098
rect 440004 -4342 440186 -4106
rect 440422 -4342 440604 -4106
rect 440004 -4426 440604 -4342
rect 440004 -4662 440186 -4426
rect 440422 -4662 440604 -4426
rect 440004 -5624 440604 -4662
rect 443604 697254 444204 709922
rect 461604 711418 462204 711440
rect 461604 711182 461786 711418
rect 462022 711182 462204 711418
rect 461604 711098 462204 711182
rect 461604 710862 461786 711098
rect 462022 710862 462204 711098
rect 458004 709538 458604 709560
rect 458004 709302 458186 709538
rect 458422 709302 458604 709538
rect 458004 709218 458604 709302
rect 458004 708982 458186 709218
rect 458422 708982 458604 709218
rect 454404 707658 455004 707680
rect 454404 707422 454586 707658
rect 454822 707422 455004 707658
rect 454404 707338 455004 707422
rect 454404 707102 454586 707338
rect 454822 707102 455004 707338
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7162 425786 -6926
rect 426022 -7162 426204 -6926
rect 425604 -7246 426204 -7162
rect 425604 -7482 425786 -7246
rect 426022 -7482 426204 -7246
rect 425604 -7504 426204 -7482
rect 443604 -5986 444204 12698
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 454404 672054 455004 707102
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3166 455004 23498
rect 454404 -3402 454586 -3166
rect 454822 -3402 455004 -3166
rect 454404 -3486 455004 -3402
rect 454404 -3722 454586 -3486
rect 454822 -3722 455004 -3486
rect 454404 -3744 455004 -3722
rect 458004 675654 458604 708982
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 461604 679254 462204 710862
rect 479604 710478 480204 711440
rect 479604 710242 479786 710478
rect 480022 710242 480204 710478
rect 479604 710158 480204 710242
rect 479604 709922 479786 710158
rect 480022 709922 480204 710158
rect 476004 708598 476604 709560
rect 476004 708362 476186 708598
rect 476422 708362 476604 708598
rect 476004 708278 476604 708362
rect 476004 708042 476186 708278
rect 476422 708042 476604 708278
rect 472404 706718 473004 707680
rect 472404 706482 472586 706718
rect 472822 706482 473004 706718
rect 472404 706398 473004 706482
rect 472404 706162 472586 706398
rect 472822 706162 473004 706398
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 387749 462204 390698
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 387749 469404 397898
rect 472404 690054 473004 706162
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 387749 473004 401498
rect 476004 693654 476604 708042
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 479604 697254 480204 709922
rect 497604 711418 498204 711440
rect 497604 711182 497786 711418
rect 498022 711182 498204 711418
rect 497604 711098 498204 711182
rect 497604 710862 497786 711098
rect 498022 710862 498204 711098
rect 494004 709538 494604 709560
rect 494004 709302 494186 709538
rect 494422 709302 494604 709538
rect 494004 709218 494604 709302
rect 494004 708982 494186 709218
rect 494422 708982 494604 709218
rect 490404 707658 491004 707680
rect 490404 707422 490586 707658
rect 490822 707422 491004 707658
rect 490404 707338 491004 707422
rect 490404 707102 490586 707338
rect 490822 707102 491004 707338
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 554964 480204 588698
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 554964 487404 559898
rect 490404 672054 491004 707102
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 554964 491004 563498
rect 494004 675654 494604 708982
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 554964 494604 567098
rect 497604 679254 498204 710862
rect 515604 710478 516204 711440
rect 515604 710242 515786 710478
rect 516022 710242 516204 710478
rect 515604 710158 516204 710242
rect 515604 709922 515786 710158
rect 516022 709922 516204 710158
rect 512004 708598 512604 709560
rect 512004 708362 512186 708598
rect 512422 708362 512604 708598
rect 512004 708278 512604 708362
rect 512004 708042 512186 708278
rect 512422 708042 512604 708278
rect 508404 706718 509004 707680
rect 508404 706482 508586 706718
rect 508822 706482 509004 706718
rect 508404 706398 509004 706482
rect 508404 706162 508586 706398
rect 508822 706162 509004 706398
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 554964 498204 570698
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 554964 505404 577898
rect 508404 690054 509004 706162
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 554964 509004 581498
rect 512004 693654 512604 708042
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 485438 542454 485758 542476
rect 485438 542218 485480 542454
rect 485716 542218 485758 542454
rect 485438 542134 485758 542218
rect 485438 541898 485480 542134
rect 485716 541898 485758 542134
rect 485438 541876 485758 541898
rect 490498 524454 490818 524476
rect 490498 524218 490540 524454
rect 490776 524218 490818 524454
rect 490498 524134 490818 524218
rect 490498 523898 490540 524134
rect 490776 523898 490818 524134
rect 490498 523876 490818 523898
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 387749 476604 405098
rect 479604 517254 480204 519800
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 387749 480204 408698
rect 486804 488454 487404 519800
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 387749 487404 415898
rect 490404 492054 491004 519800
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 387749 491004 419498
rect 494004 495654 494604 519800
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387749 494604 423098
rect 497604 499254 498204 519800
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 387749 498204 390698
rect 504804 506454 505404 519800
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 387749 505404 397898
rect 508404 510054 509004 519800
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 479568 380454 479888 380476
rect 479568 380218 479610 380454
rect 479846 380218 479888 380454
rect 479568 380134 479888 380218
rect 479568 379898 479610 380134
rect 479846 379898 479888 380134
rect 479568 379876 479888 379898
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 464208 362454 464528 362476
rect 464208 362218 464250 362454
rect 464486 362218 464528 362454
rect 464208 362134 464528 362218
rect 464208 361898 464250 362134
rect 464486 361898 464528 362134
rect 464208 361876 464528 361898
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 479568 344454 479888 344476
rect 479568 344218 479610 344454
rect 479846 344218 479888 344454
rect 479568 344134 479888 344218
rect 479568 343898 479610 344134
rect 479846 343898 479888 344134
rect 479568 343876 479888 343898
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -5046 458604 27098
rect 458004 -5282 458186 -5046
rect 458422 -5282 458604 -5046
rect 458004 -5366 458604 -5282
rect 458004 -5602 458186 -5366
rect 458422 -5602 458604 -5366
rect 458004 -5624 458604 -5602
rect 461604 319254 462204 339800
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6222 443786 -5986
rect 444022 -6222 444204 -5986
rect 443604 -6306 444204 -6222
rect 443604 -6542 443786 -6306
rect 444022 -6542 444204 -6306
rect 443604 -7504 444204 -6542
rect 461604 -6926 462204 30698
rect 468804 326454 469404 339800
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 472404 330054 473004 339800
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2226 473004 5498
rect 472404 -2462 472586 -2226
rect 472822 -2462 473004 -2226
rect 472404 -2546 473004 -2462
rect 472404 -2782 472586 -2546
rect 472822 -2782 473004 -2546
rect 472404 -3744 473004 -2782
rect 476004 333654 476604 339800
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4106 476604 9098
rect 476004 -4342 476186 -4106
rect 476422 -4342 476604 -4106
rect 476004 -4426 476604 -4342
rect 476004 -4662 476186 -4426
rect 476422 -4662 476604 -4426
rect 476004 -5624 476604 -4662
rect 479604 337254 480204 339800
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7162 461786 -6926
rect 462022 -7162 462204 -6926
rect 461604 -7246 462204 -7162
rect 461604 -7482 461786 -7246
rect 462022 -7482 462204 -7246
rect 461604 -7504 462204 -7482
rect 479604 -5986 480204 12698
rect 486804 308454 487404 339800
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 490404 312054 491004 339800
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3166 491004 23498
rect 490404 -3402 490586 -3166
rect 490822 -3402 491004 -3166
rect 490404 -3486 491004 -3402
rect 490404 -3722 490586 -3486
rect 490822 -3722 491004 -3486
rect 490404 -3744 491004 -3722
rect 494004 315654 494604 339800
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -5046 494604 27098
rect 494004 -5282 494186 -5046
rect 494422 -5282 494604 -5046
rect 494004 -5366 494604 -5282
rect 494004 -5602 494186 -5366
rect 494422 -5602 494604 -5366
rect 494004 -5624 494604 -5602
rect 497604 319254 498204 339800
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6222 479786 -5986
rect 480022 -6222 480204 -5986
rect 479604 -6306 480204 -6222
rect 479604 -6542 479786 -6306
rect 480022 -6542 480204 -6306
rect 479604 -7504 480204 -6542
rect 497604 -6926 498204 30698
rect 504804 326454 505404 339800
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2226 509004 5498
rect 508404 -2462 508586 -2226
rect 508822 -2462 509004 -2226
rect 508404 -2546 509004 -2462
rect 508404 -2782 508586 -2546
rect 508822 -2782 509004 -2546
rect 508404 -3744 509004 -2782
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4106 512604 9098
rect 512004 -4342 512186 -4106
rect 512422 -4342 512604 -4106
rect 512004 -4426 512604 -4342
rect 512004 -4662 512186 -4426
rect 512422 -4662 512604 -4426
rect 512004 -5624 512604 -4662
rect 515604 697254 516204 709922
rect 533604 711418 534204 711440
rect 533604 711182 533786 711418
rect 534022 711182 534204 711418
rect 533604 711098 534204 711182
rect 533604 710862 533786 711098
rect 534022 710862 534204 711098
rect 530004 709538 530604 709560
rect 530004 709302 530186 709538
rect 530422 709302 530604 709538
rect 530004 709218 530604 709302
rect 530004 708982 530186 709218
rect 530422 708982 530604 709218
rect 526404 707658 527004 707680
rect 526404 707422 526586 707658
rect 526822 707422 527004 707658
rect 526404 707338 527004 707422
rect 526404 707102 526586 707338
rect 526822 707102 527004 707338
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7162 497786 -6926
rect 498022 -7162 498204 -6926
rect 497604 -7246 498204 -7162
rect 497604 -7482 497786 -7246
rect 498022 -7482 498204 -7246
rect 497604 -7504 498204 -7482
rect 515604 -5986 516204 12698
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 526404 672054 527004 707102
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3166 527004 23498
rect 526404 -3402 526586 -3166
rect 526822 -3402 527004 -3166
rect 526404 -3486 527004 -3402
rect 526404 -3722 526586 -3486
rect 526822 -3722 527004 -3486
rect 526404 -3744 527004 -3722
rect 530004 675654 530604 708982
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -5046 530604 27098
rect 530004 -5282 530186 -5046
rect 530422 -5282 530604 -5046
rect 530004 -5366 530604 -5282
rect 530004 -5602 530186 -5366
rect 530422 -5602 530604 -5366
rect 530004 -5624 530604 -5602
rect 533604 679254 534204 710862
rect 551604 710478 552204 711440
rect 551604 710242 551786 710478
rect 552022 710242 552204 710478
rect 551604 710158 552204 710242
rect 551604 709922 551786 710158
rect 552022 709922 552204 710158
rect 548004 708598 548604 709560
rect 548004 708362 548186 708598
rect 548422 708362 548604 708598
rect 548004 708278 548604 708362
rect 548004 708042 548186 708278
rect 548422 708042 548604 708278
rect 544404 706718 545004 707680
rect 544404 706482 544586 706718
rect 544822 706482 545004 706718
rect 544404 706398 545004 706482
rect 544404 706162 544586 706398
rect 544822 706162 545004 706398
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6222 515786 -5986
rect 516022 -6222 516204 -5986
rect 515604 -6306 516204 -6222
rect 515604 -6542 515786 -6306
rect 516022 -6542 516204 -6306
rect 515604 -7504 516204 -6542
rect 533604 -6926 534204 30698
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 544404 690054 545004 706162
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2226 545004 5498
rect 544404 -2462 544586 -2226
rect 544822 -2462 545004 -2226
rect 544404 -2546 545004 -2462
rect 544404 -2782 544586 -2546
rect 544822 -2782 545004 -2546
rect 544404 -3744 545004 -2782
rect 548004 693654 548604 708042
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4106 548604 9098
rect 548004 -4342 548186 -4106
rect 548422 -4342 548604 -4106
rect 548004 -4426 548604 -4342
rect 548004 -4662 548186 -4426
rect 548422 -4662 548604 -4426
rect 548004 -5624 548604 -4662
rect 551604 697254 552204 709922
rect 569604 711418 570204 711440
rect 569604 711182 569786 711418
rect 570022 711182 570204 711418
rect 569604 711098 570204 711182
rect 569604 710862 569786 711098
rect 570022 710862 570204 711098
rect 566004 709538 566604 709560
rect 566004 709302 566186 709538
rect 566422 709302 566604 709538
rect 566004 709218 566604 709302
rect 566004 708982 566186 709218
rect 566422 708982 566604 709218
rect 562404 707658 563004 707680
rect 562404 707422 562586 707658
rect 562822 707422 563004 707658
rect 562404 707338 563004 707422
rect 562404 707102 562586 707338
rect 562822 707102 563004 707338
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7162 533786 -6926
rect 534022 -7162 534204 -6926
rect 533604 -7246 534204 -7162
rect 533604 -7482 533786 -7246
rect 534022 -7482 534204 -7246
rect 533604 -7504 534204 -7482
rect 551604 -5986 552204 12698
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 562404 672054 563004 707102
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3166 563004 23498
rect 562404 -3402 562586 -3166
rect 562822 -3402 563004 -3166
rect 562404 -3486 563004 -3402
rect 562404 -3722 562586 -3486
rect 562822 -3722 563004 -3486
rect 562404 -3744 563004 -3722
rect 566004 675654 566604 708982
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -5046 566604 27098
rect 566004 -5282 566186 -5046
rect 566422 -5282 566604 -5046
rect 566004 -5366 566604 -5282
rect 566004 -5602 566186 -5366
rect 566422 -5602 566604 -5366
rect 566004 -5624 566604 -5602
rect 569604 679254 570204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 580404 706718 581004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 580404 706482 580586 706718
rect 580822 706482 581004 706718
rect 580404 706398 581004 706482
rect 580404 706162 580586 706398
rect 580822 706162 581004 706398
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6222 551786 -5986
rect 552022 -6222 552204 -5986
rect 551604 -6306 552204 -6222
rect 551604 -6542 551786 -6306
rect 552022 -6542 552204 -6306
rect 551604 -7504 552204 -6542
rect 569604 -6926 570204 30698
rect 576804 704838 577404 705800
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 580404 690054 581004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2226 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 690054 587800 706162
rect 587200 689818 587382 690054
rect 587618 689818 587800 690054
rect 587200 689734 587800 689818
rect 587200 689498 587382 689734
rect 587618 689498 587800 689734
rect 587200 654054 587800 689498
rect 587200 653818 587382 654054
rect 587618 653818 587800 654054
rect 587200 653734 587800 653818
rect 587200 653498 587382 653734
rect 587618 653498 587800 653734
rect 587200 618054 587800 653498
rect 587200 617818 587382 618054
rect 587618 617818 587800 618054
rect 587200 617734 587800 617818
rect 587200 617498 587382 617734
rect 587618 617498 587800 617734
rect 587200 582054 587800 617498
rect 587200 581818 587382 582054
rect 587618 581818 587800 582054
rect 587200 581734 587800 581818
rect 587200 581498 587382 581734
rect 587618 581498 587800 581734
rect 587200 546054 587800 581498
rect 587200 545818 587382 546054
rect 587618 545818 587800 546054
rect 587200 545734 587800 545818
rect 587200 545498 587382 545734
rect 587618 545498 587800 545734
rect 587200 510054 587800 545498
rect 587200 509818 587382 510054
rect 587618 509818 587800 510054
rect 587200 509734 587800 509818
rect 587200 509498 587382 509734
rect 587618 509498 587800 509734
rect 587200 474054 587800 509498
rect 587200 473818 587382 474054
rect 587618 473818 587800 474054
rect 587200 473734 587800 473818
rect 587200 473498 587382 473734
rect 587618 473498 587800 473734
rect 587200 438054 587800 473498
rect 587200 437818 587382 438054
rect 587618 437818 587800 438054
rect 587200 437734 587800 437818
rect 587200 437498 587382 437734
rect 587618 437498 587800 437734
rect 587200 402054 587800 437498
rect 587200 401818 587382 402054
rect 587618 401818 587800 402054
rect 587200 401734 587800 401818
rect 587200 401498 587382 401734
rect 587618 401498 587800 401734
rect 587200 366054 587800 401498
rect 587200 365818 587382 366054
rect 587618 365818 587800 366054
rect 587200 365734 587800 365818
rect 587200 365498 587382 365734
rect 587618 365498 587800 365734
rect 587200 330054 587800 365498
rect 587200 329818 587382 330054
rect 587618 329818 587800 330054
rect 587200 329734 587800 329818
rect 587200 329498 587382 329734
rect 587618 329498 587800 329734
rect 587200 294054 587800 329498
rect 587200 293818 587382 294054
rect 587618 293818 587800 294054
rect 587200 293734 587800 293818
rect 587200 293498 587382 293734
rect 587618 293498 587800 293734
rect 587200 258054 587800 293498
rect 587200 257818 587382 258054
rect 587618 257818 587800 258054
rect 587200 257734 587800 257818
rect 587200 257498 587382 257734
rect 587618 257498 587800 257734
rect 587200 222054 587800 257498
rect 587200 221818 587382 222054
rect 587618 221818 587800 222054
rect 587200 221734 587800 221818
rect 587200 221498 587382 221734
rect 587618 221498 587800 221734
rect 587200 186054 587800 221498
rect 587200 185818 587382 186054
rect 587618 185818 587800 186054
rect 587200 185734 587800 185818
rect 587200 185498 587382 185734
rect 587618 185498 587800 185734
rect 587200 150054 587800 185498
rect 587200 149818 587382 150054
rect 587618 149818 587800 150054
rect 587200 149734 587800 149818
rect 587200 149498 587382 149734
rect 587618 149498 587800 149734
rect 587200 114054 587800 149498
rect 587200 113818 587382 114054
rect 587618 113818 587800 114054
rect 587200 113734 587800 113818
rect 587200 113498 587382 113734
rect 587618 113498 587800 113734
rect 587200 78054 587800 113498
rect 587200 77818 587382 78054
rect 587618 77818 587800 78054
rect 587200 77734 587800 77818
rect 587200 77498 587382 77734
rect 587618 77498 587800 77734
rect 587200 42054 587800 77498
rect 587200 41818 587382 42054
rect 587618 41818 587800 42054
rect 587200 41734 587800 41818
rect 587200 41498 587382 41734
rect 587618 41498 587800 41734
rect 587200 6054 587800 41498
rect 587200 5818 587382 6054
rect 587618 5818 587800 6054
rect 587200 5734 587800 5818
rect 587200 5498 587382 5734
rect 587618 5498 587800 5734
rect 580404 -2462 580586 -2226
rect 580822 -2462 581004 -2226
rect 580404 -2546 581004 -2462
rect 580404 -2782 580586 -2546
rect 580822 -2782 581004 -2546
rect 580404 -3744 581004 -2782
rect 587200 -2226 587800 5498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 672054 588740 707102
rect 588140 671818 588322 672054
rect 588558 671818 588740 672054
rect 588140 671734 588740 671818
rect 588140 671498 588322 671734
rect 588558 671498 588740 671734
rect 588140 636054 588740 671498
rect 588140 635818 588322 636054
rect 588558 635818 588740 636054
rect 588140 635734 588740 635818
rect 588140 635498 588322 635734
rect 588558 635498 588740 635734
rect 588140 600054 588740 635498
rect 588140 599818 588322 600054
rect 588558 599818 588740 600054
rect 588140 599734 588740 599818
rect 588140 599498 588322 599734
rect 588558 599498 588740 599734
rect 588140 564054 588740 599498
rect 588140 563818 588322 564054
rect 588558 563818 588740 564054
rect 588140 563734 588740 563818
rect 588140 563498 588322 563734
rect 588558 563498 588740 563734
rect 588140 528054 588740 563498
rect 588140 527818 588322 528054
rect 588558 527818 588740 528054
rect 588140 527734 588740 527818
rect 588140 527498 588322 527734
rect 588558 527498 588740 527734
rect 588140 492054 588740 527498
rect 588140 491818 588322 492054
rect 588558 491818 588740 492054
rect 588140 491734 588740 491818
rect 588140 491498 588322 491734
rect 588558 491498 588740 491734
rect 588140 456054 588740 491498
rect 588140 455818 588322 456054
rect 588558 455818 588740 456054
rect 588140 455734 588740 455818
rect 588140 455498 588322 455734
rect 588558 455498 588740 455734
rect 588140 420054 588740 455498
rect 588140 419818 588322 420054
rect 588558 419818 588740 420054
rect 588140 419734 588740 419818
rect 588140 419498 588322 419734
rect 588558 419498 588740 419734
rect 588140 384054 588740 419498
rect 588140 383818 588322 384054
rect 588558 383818 588740 384054
rect 588140 383734 588740 383818
rect 588140 383498 588322 383734
rect 588558 383498 588740 383734
rect 588140 348054 588740 383498
rect 588140 347818 588322 348054
rect 588558 347818 588740 348054
rect 588140 347734 588740 347818
rect 588140 347498 588322 347734
rect 588558 347498 588740 347734
rect 588140 312054 588740 347498
rect 588140 311818 588322 312054
rect 588558 311818 588740 312054
rect 588140 311734 588740 311818
rect 588140 311498 588322 311734
rect 588558 311498 588740 311734
rect 588140 276054 588740 311498
rect 588140 275818 588322 276054
rect 588558 275818 588740 276054
rect 588140 275734 588740 275818
rect 588140 275498 588322 275734
rect 588558 275498 588740 275734
rect 588140 240054 588740 275498
rect 588140 239818 588322 240054
rect 588558 239818 588740 240054
rect 588140 239734 588740 239818
rect 588140 239498 588322 239734
rect 588558 239498 588740 239734
rect 588140 204054 588740 239498
rect 588140 203818 588322 204054
rect 588558 203818 588740 204054
rect 588140 203734 588740 203818
rect 588140 203498 588322 203734
rect 588558 203498 588740 203734
rect 588140 168054 588740 203498
rect 588140 167818 588322 168054
rect 588558 167818 588740 168054
rect 588140 167734 588740 167818
rect 588140 167498 588322 167734
rect 588558 167498 588740 167734
rect 588140 132054 588740 167498
rect 588140 131818 588322 132054
rect 588558 131818 588740 132054
rect 588140 131734 588740 131818
rect 588140 131498 588322 131734
rect 588558 131498 588740 131734
rect 588140 96054 588740 131498
rect 588140 95818 588322 96054
rect 588558 95818 588740 96054
rect 588140 95734 588740 95818
rect 588140 95498 588322 95734
rect 588558 95498 588740 95734
rect 588140 60054 588740 95498
rect 588140 59818 588322 60054
rect 588558 59818 588740 60054
rect 588140 59734 588740 59818
rect 588140 59498 588322 59734
rect 588558 59498 588740 59734
rect 588140 24054 588740 59498
rect 588140 23818 588322 24054
rect 588558 23818 588740 24054
rect 588140 23734 588740 23818
rect 588140 23498 588322 23734
rect 588558 23498 588740 23734
rect 588140 -3166 588740 23498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 693654 589680 708042
rect 589080 693418 589262 693654
rect 589498 693418 589680 693654
rect 589080 693334 589680 693418
rect 589080 693098 589262 693334
rect 589498 693098 589680 693334
rect 589080 657654 589680 693098
rect 589080 657418 589262 657654
rect 589498 657418 589680 657654
rect 589080 657334 589680 657418
rect 589080 657098 589262 657334
rect 589498 657098 589680 657334
rect 589080 621654 589680 657098
rect 589080 621418 589262 621654
rect 589498 621418 589680 621654
rect 589080 621334 589680 621418
rect 589080 621098 589262 621334
rect 589498 621098 589680 621334
rect 589080 585654 589680 621098
rect 589080 585418 589262 585654
rect 589498 585418 589680 585654
rect 589080 585334 589680 585418
rect 589080 585098 589262 585334
rect 589498 585098 589680 585334
rect 589080 549654 589680 585098
rect 589080 549418 589262 549654
rect 589498 549418 589680 549654
rect 589080 549334 589680 549418
rect 589080 549098 589262 549334
rect 589498 549098 589680 549334
rect 589080 513654 589680 549098
rect 589080 513418 589262 513654
rect 589498 513418 589680 513654
rect 589080 513334 589680 513418
rect 589080 513098 589262 513334
rect 589498 513098 589680 513334
rect 589080 477654 589680 513098
rect 589080 477418 589262 477654
rect 589498 477418 589680 477654
rect 589080 477334 589680 477418
rect 589080 477098 589262 477334
rect 589498 477098 589680 477334
rect 589080 441654 589680 477098
rect 589080 441418 589262 441654
rect 589498 441418 589680 441654
rect 589080 441334 589680 441418
rect 589080 441098 589262 441334
rect 589498 441098 589680 441334
rect 589080 405654 589680 441098
rect 589080 405418 589262 405654
rect 589498 405418 589680 405654
rect 589080 405334 589680 405418
rect 589080 405098 589262 405334
rect 589498 405098 589680 405334
rect 589080 369654 589680 405098
rect 589080 369418 589262 369654
rect 589498 369418 589680 369654
rect 589080 369334 589680 369418
rect 589080 369098 589262 369334
rect 589498 369098 589680 369334
rect 589080 333654 589680 369098
rect 589080 333418 589262 333654
rect 589498 333418 589680 333654
rect 589080 333334 589680 333418
rect 589080 333098 589262 333334
rect 589498 333098 589680 333334
rect 589080 297654 589680 333098
rect 589080 297418 589262 297654
rect 589498 297418 589680 297654
rect 589080 297334 589680 297418
rect 589080 297098 589262 297334
rect 589498 297098 589680 297334
rect 589080 261654 589680 297098
rect 589080 261418 589262 261654
rect 589498 261418 589680 261654
rect 589080 261334 589680 261418
rect 589080 261098 589262 261334
rect 589498 261098 589680 261334
rect 589080 225654 589680 261098
rect 589080 225418 589262 225654
rect 589498 225418 589680 225654
rect 589080 225334 589680 225418
rect 589080 225098 589262 225334
rect 589498 225098 589680 225334
rect 589080 189654 589680 225098
rect 589080 189418 589262 189654
rect 589498 189418 589680 189654
rect 589080 189334 589680 189418
rect 589080 189098 589262 189334
rect 589498 189098 589680 189334
rect 589080 153654 589680 189098
rect 589080 153418 589262 153654
rect 589498 153418 589680 153654
rect 589080 153334 589680 153418
rect 589080 153098 589262 153334
rect 589498 153098 589680 153334
rect 589080 117654 589680 153098
rect 589080 117418 589262 117654
rect 589498 117418 589680 117654
rect 589080 117334 589680 117418
rect 589080 117098 589262 117334
rect 589498 117098 589680 117334
rect 589080 81654 589680 117098
rect 589080 81418 589262 81654
rect 589498 81418 589680 81654
rect 589080 81334 589680 81418
rect 589080 81098 589262 81334
rect 589498 81098 589680 81334
rect 589080 45654 589680 81098
rect 589080 45418 589262 45654
rect 589498 45418 589680 45654
rect 589080 45334 589680 45418
rect 589080 45098 589262 45334
rect 589498 45098 589680 45334
rect 589080 9654 589680 45098
rect 589080 9418 589262 9654
rect 589498 9418 589680 9654
rect 589080 9334 589680 9418
rect 589080 9098 589262 9334
rect 589498 9098 589680 9334
rect 589080 -4106 589680 9098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 675654 590620 708982
rect 590020 675418 590202 675654
rect 590438 675418 590620 675654
rect 590020 675334 590620 675418
rect 590020 675098 590202 675334
rect 590438 675098 590620 675334
rect 590020 639654 590620 675098
rect 590020 639418 590202 639654
rect 590438 639418 590620 639654
rect 590020 639334 590620 639418
rect 590020 639098 590202 639334
rect 590438 639098 590620 639334
rect 590020 603654 590620 639098
rect 590020 603418 590202 603654
rect 590438 603418 590620 603654
rect 590020 603334 590620 603418
rect 590020 603098 590202 603334
rect 590438 603098 590620 603334
rect 590020 567654 590620 603098
rect 590020 567418 590202 567654
rect 590438 567418 590620 567654
rect 590020 567334 590620 567418
rect 590020 567098 590202 567334
rect 590438 567098 590620 567334
rect 590020 531654 590620 567098
rect 590020 531418 590202 531654
rect 590438 531418 590620 531654
rect 590020 531334 590620 531418
rect 590020 531098 590202 531334
rect 590438 531098 590620 531334
rect 590020 495654 590620 531098
rect 590020 495418 590202 495654
rect 590438 495418 590620 495654
rect 590020 495334 590620 495418
rect 590020 495098 590202 495334
rect 590438 495098 590620 495334
rect 590020 459654 590620 495098
rect 590020 459418 590202 459654
rect 590438 459418 590620 459654
rect 590020 459334 590620 459418
rect 590020 459098 590202 459334
rect 590438 459098 590620 459334
rect 590020 423654 590620 459098
rect 590020 423418 590202 423654
rect 590438 423418 590620 423654
rect 590020 423334 590620 423418
rect 590020 423098 590202 423334
rect 590438 423098 590620 423334
rect 590020 387654 590620 423098
rect 590020 387418 590202 387654
rect 590438 387418 590620 387654
rect 590020 387334 590620 387418
rect 590020 387098 590202 387334
rect 590438 387098 590620 387334
rect 590020 351654 590620 387098
rect 590020 351418 590202 351654
rect 590438 351418 590620 351654
rect 590020 351334 590620 351418
rect 590020 351098 590202 351334
rect 590438 351098 590620 351334
rect 590020 315654 590620 351098
rect 590020 315418 590202 315654
rect 590438 315418 590620 315654
rect 590020 315334 590620 315418
rect 590020 315098 590202 315334
rect 590438 315098 590620 315334
rect 590020 279654 590620 315098
rect 590020 279418 590202 279654
rect 590438 279418 590620 279654
rect 590020 279334 590620 279418
rect 590020 279098 590202 279334
rect 590438 279098 590620 279334
rect 590020 243654 590620 279098
rect 590020 243418 590202 243654
rect 590438 243418 590620 243654
rect 590020 243334 590620 243418
rect 590020 243098 590202 243334
rect 590438 243098 590620 243334
rect 590020 207654 590620 243098
rect 590020 207418 590202 207654
rect 590438 207418 590620 207654
rect 590020 207334 590620 207418
rect 590020 207098 590202 207334
rect 590438 207098 590620 207334
rect 590020 171654 590620 207098
rect 590020 171418 590202 171654
rect 590438 171418 590620 171654
rect 590020 171334 590620 171418
rect 590020 171098 590202 171334
rect 590438 171098 590620 171334
rect 590020 135654 590620 171098
rect 590020 135418 590202 135654
rect 590438 135418 590620 135654
rect 590020 135334 590620 135418
rect 590020 135098 590202 135334
rect 590438 135098 590620 135334
rect 590020 99654 590620 135098
rect 590020 99418 590202 99654
rect 590438 99418 590620 99654
rect 590020 99334 590620 99418
rect 590020 99098 590202 99334
rect 590438 99098 590620 99334
rect 590020 63654 590620 99098
rect 590020 63418 590202 63654
rect 590438 63418 590620 63654
rect 590020 63334 590620 63418
rect 590020 63098 590202 63334
rect 590438 63098 590620 63334
rect 590020 27654 590620 63098
rect 590020 27418 590202 27654
rect 590438 27418 590620 27654
rect 590020 27334 590620 27418
rect 590020 27098 590202 27334
rect 590438 27098 590620 27334
rect 590020 -5046 590620 27098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 697254 591560 709922
rect 590960 697018 591142 697254
rect 591378 697018 591560 697254
rect 590960 696934 591560 697018
rect 590960 696698 591142 696934
rect 591378 696698 591560 696934
rect 590960 661254 591560 696698
rect 590960 661018 591142 661254
rect 591378 661018 591560 661254
rect 590960 660934 591560 661018
rect 590960 660698 591142 660934
rect 591378 660698 591560 660934
rect 590960 625254 591560 660698
rect 590960 625018 591142 625254
rect 591378 625018 591560 625254
rect 590960 624934 591560 625018
rect 590960 624698 591142 624934
rect 591378 624698 591560 624934
rect 590960 589254 591560 624698
rect 590960 589018 591142 589254
rect 591378 589018 591560 589254
rect 590960 588934 591560 589018
rect 590960 588698 591142 588934
rect 591378 588698 591560 588934
rect 590960 553254 591560 588698
rect 590960 553018 591142 553254
rect 591378 553018 591560 553254
rect 590960 552934 591560 553018
rect 590960 552698 591142 552934
rect 591378 552698 591560 552934
rect 590960 517254 591560 552698
rect 590960 517018 591142 517254
rect 591378 517018 591560 517254
rect 590960 516934 591560 517018
rect 590960 516698 591142 516934
rect 591378 516698 591560 516934
rect 590960 481254 591560 516698
rect 590960 481018 591142 481254
rect 591378 481018 591560 481254
rect 590960 480934 591560 481018
rect 590960 480698 591142 480934
rect 591378 480698 591560 480934
rect 590960 445254 591560 480698
rect 590960 445018 591142 445254
rect 591378 445018 591560 445254
rect 590960 444934 591560 445018
rect 590960 444698 591142 444934
rect 591378 444698 591560 444934
rect 590960 409254 591560 444698
rect 590960 409018 591142 409254
rect 591378 409018 591560 409254
rect 590960 408934 591560 409018
rect 590960 408698 591142 408934
rect 591378 408698 591560 408934
rect 590960 373254 591560 408698
rect 590960 373018 591142 373254
rect 591378 373018 591560 373254
rect 590960 372934 591560 373018
rect 590960 372698 591142 372934
rect 591378 372698 591560 372934
rect 590960 337254 591560 372698
rect 590960 337018 591142 337254
rect 591378 337018 591560 337254
rect 590960 336934 591560 337018
rect 590960 336698 591142 336934
rect 591378 336698 591560 336934
rect 590960 301254 591560 336698
rect 590960 301018 591142 301254
rect 591378 301018 591560 301254
rect 590960 300934 591560 301018
rect 590960 300698 591142 300934
rect 591378 300698 591560 300934
rect 590960 265254 591560 300698
rect 590960 265018 591142 265254
rect 591378 265018 591560 265254
rect 590960 264934 591560 265018
rect 590960 264698 591142 264934
rect 591378 264698 591560 264934
rect 590960 229254 591560 264698
rect 590960 229018 591142 229254
rect 591378 229018 591560 229254
rect 590960 228934 591560 229018
rect 590960 228698 591142 228934
rect 591378 228698 591560 228934
rect 590960 193254 591560 228698
rect 590960 193018 591142 193254
rect 591378 193018 591560 193254
rect 590960 192934 591560 193018
rect 590960 192698 591142 192934
rect 591378 192698 591560 192934
rect 590960 157254 591560 192698
rect 590960 157018 591142 157254
rect 591378 157018 591560 157254
rect 590960 156934 591560 157018
rect 590960 156698 591142 156934
rect 591378 156698 591560 156934
rect 590960 121254 591560 156698
rect 590960 121018 591142 121254
rect 591378 121018 591560 121254
rect 590960 120934 591560 121018
rect 590960 120698 591142 120934
rect 591378 120698 591560 120934
rect 590960 85254 591560 120698
rect 590960 85018 591142 85254
rect 591378 85018 591560 85254
rect 590960 84934 591560 85018
rect 590960 84698 591142 84934
rect 591378 84698 591560 84934
rect 590960 49254 591560 84698
rect 590960 49018 591142 49254
rect 591378 49018 591560 49254
rect 590960 48934 591560 49018
rect 590960 48698 591142 48934
rect 591378 48698 591560 48934
rect 590960 13254 591560 48698
rect 590960 13018 591142 13254
rect 591378 13018 591560 13254
rect 590960 12934 591560 13018
rect 590960 12698 591142 12934
rect 591378 12698 591560 12934
rect 590960 -5986 591560 12698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 679254 592500 710862
rect 591900 679018 592082 679254
rect 592318 679018 592500 679254
rect 591900 678934 592500 679018
rect 591900 678698 592082 678934
rect 592318 678698 592500 678934
rect 591900 643254 592500 678698
rect 591900 643018 592082 643254
rect 592318 643018 592500 643254
rect 591900 642934 592500 643018
rect 591900 642698 592082 642934
rect 592318 642698 592500 642934
rect 591900 607254 592500 642698
rect 591900 607018 592082 607254
rect 592318 607018 592500 607254
rect 591900 606934 592500 607018
rect 591900 606698 592082 606934
rect 592318 606698 592500 606934
rect 591900 571254 592500 606698
rect 591900 571018 592082 571254
rect 592318 571018 592500 571254
rect 591900 570934 592500 571018
rect 591900 570698 592082 570934
rect 592318 570698 592500 570934
rect 591900 535254 592500 570698
rect 591900 535018 592082 535254
rect 592318 535018 592500 535254
rect 591900 534934 592500 535018
rect 591900 534698 592082 534934
rect 592318 534698 592500 534934
rect 591900 499254 592500 534698
rect 591900 499018 592082 499254
rect 592318 499018 592500 499254
rect 591900 498934 592500 499018
rect 591900 498698 592082 498934
rect 592318 498698 592500 498934
rect 591900 463254 592500 498698
rect 591900 463018 592082 463254
rect 592318 463018 592500 463254
rect 591900 462934 592500 463018
rect 591900 462698 592082 462934
rect 592318 462698 592500 462934
rect 591900 427254 592500 462698
rect 591900 427018 592082 427254
rect 592318 427018 592500 427254
rect 591900 426934 592500 427018
rect 591900 426698 592082 426934
rect 592318 426698 592500 426934
rect 591900 391254 592500 426698
rect 591900 391018 592082 391254
rect 592318 391018 592500 391254
rect 591900 390934 592500 391018
rect 591900 390698 592082 390934
rect 592318 390698 592500 390934
rect 591900 355254 592500 390698
rect 591900 355018 592082 355254
rect 592318 355018 592500 355254
rect 591900 354934 592500 355018
rect 591900 354698 592082 354934
rect 592318 354698 592500 354934
rect 591900 319254 592500 354698
rect 591900 319018 592082 319254
rect 592318 319018 592500 319254
rect 591900 318934 592500 319018
rect 591900 318698 592082 318934
rect 592318 318698 592500 318934
rect 591900 283254 592500 318698
rect 591900 283018 592082 283254
rect 592318 283018 592500 283254
rect 591900 282934 592500 283018
rect 591900 282698 592082 282934
rect 592318 282698 592500 282934
rect 591900 247254 592500 282698
rect 591900 247018 592082 247254
rect 592318 247018 592500 247254
rect 591900 246934 592500 247018
rect 591900 246698 592082 246934
rect 592318 246698 592500 246934
rect 591900 211254 592500 246698
rect 591900 211018 592082 211254
rect 592318 211018 592500 211254
rect 591900 210934 592500 211018
rect 591900 210698 592082 210934
rect 592318 210698 592500 210934
rect 591900 175254 592500 210698
rect 591900 175018 592082 175254
rect 592318 175018 592500 175254
rect 591900 174934 592500 175018
rect 591900 174698 592082 174934
rect 592318 174698 592500 174934
rect 591900 139254 592500 174698
rect 591900 139018 592082 139254
rect 592318 139018 592500 139254
rect 591900 138934 592500 139018
rect 591900 138698 592082 138934
rect 592318 138698 592500 138934
rect 591900 103254 592500 138698
rect 591900 103018 592082 103254
rect 592318 103018 592500 103254
rect 591900 102934 592500 103018
rect 591900 102698 592082 102934
rect 592318 102698 592500 102934
rect 591900 67254 592500 102698
rect 591900 67018 592082 67254
rect 592318 67018 592500 67254
rect 591900 66934 592500 67018
rect 591900 66698 592082 66934
rect 592318 66698 592500 66934
rect 591900 31254 592500 66698
rect 591900 31018 592082 31254
rect 592318 31018 592500 31254
rect 591900 30934 592500 31018
rect 591900 30698 592082 30934
rect 592318 30698 592500 30934
rect 569604 -7162 569786 -6926
rect 570022 -7162 570204 -6926
rect 569604 -7246 570204 -7162
rect 569604 -7482 569786 -7246
rect 570022 -7482 570204 -7246
rect 569604 -7504 570204 -7482
rect 591900 -6926 592500 30698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 679018 -8158 679254
rect -8394 678698 -8158 678934
rect -8394 643018 -8158 643254
rect -8394 642698 -8158 642934
rect -8394 607018 -8158 607254
rect -8394 606698 -8158 606934
rect -8394 571018 -8158 571254
rect -8394 570698 -8158 570934
rect -8394 535018 -8158 535254
rect -8394 534698 -8158 534934
rect -8394 499018 -8158 499254
rect -8394 498698 -8158 498934
rect -8394 463018 -8158 463254
rect -8394 462698 -8158 462934
rect -8394 427018 -8158 427254
rect -8394 426698 -8158 426934
rect -8394 391018 -8158 391254
rect -8394 390698 -8158 390934
rect -8394 355018 -8158 355254
rect -8394 354698 -8158 354934
rect -8394 319018 -8158 319254
rect -8394 318698 -8158 318934
rect -8394 283018 -8158 283254
rect -8394 282698 -8158 282934
rect -8394 247018 -8158 247254
rect -8394 246698 -8158 246934
rect -8394 211018 -8158 211254
rect -8394 210698 -8158 210934
rect -8394 175018 -8158 175254
rect -8394 174698 -8158 174934
rect -8394 139018 -8158 139254
rect -8394 138698 -8158 138934
rect -8394 103018 -8158 103254
rect -8394 102698 -8158 102934
rect -8394 67018 -8158 67254
rect -8394 66698 -8158 66934
rect -8394 31018 -8158 31254
rect -8394 30698 -8158 30934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 11786 710242 12022 710478
rect 11786 709922 12022 710158
rect -7454 697018 -7218 697254
rect -7454 696698 -7218 696934
rect -7454 661018 -7218 661254
rect -7454 660698 -7218 660934
rect -7454 625018 -7218 625254
rect -7454 624698 -7218 624934
rect -7454 589018 -7218 589254
rect -7454 588698 -7218 588934
rect -7454 553018 -7218 553254
rect -7454 552698 -7218 552934
rect -7454 517018 -7218 517254
rect -7454 516698 -7218 516934
rect -7454 481018 -7218 481254
rect -7454 480698 -7218 480934
rect -7454 445018 -7218 445254
rect -7454 444698 -7218 444934
rect -7454 409018 -7218 409254
rect -7454 408698 -7218 408934
rect -7454 373018 -7218 373254
rect -7454 372698 -7218 372934
rect -7454 337018 -7218 337254
rect -7454 336698 -7218 336934
rect -7454 301018 -7218 301254
rect -7454 300698 -7218 300934
rect -7454 265018 -7218 265254
rect -7454 264698 -7218 264934
rect -7454 229018 -7218 229254
rect -7454 228698 -7218 228934
rect -7454 193018 -7218 193254
rect -7454 192698 -7218 192934
rect -7454 157018 -7218 157254
rect -7454 156698 -7218 156934
rect -7454 121018 -7218 121254
rect -7454 120698 -7218 120934
rect -7454 85018 -7218 85254
rect -7454 84698 -7218 84934
rect -7454 49018 -7218 49254
rect -7454 48698 -7218 48934
rect -7454 13018 -7218 13254
rect -7454 12698 -7218 12934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 675418 -6278 675654
rect -6514 675098 -6278 675334
rect -6514 639418 -6278 639654
rect -6514 639098 -6278 639334
rect -6514 603418 -6278 603654
rect -6514 603098 -6278 603334
rect -6514 567418 -6278 567654
rect -6514 567098 -6278 567334
rect -6514 531418 -6278 531654
rect -6514 531098 -6278 531334
rect -6514 495418 -6278 495654
rect -6514 495098 -6278 495334
rect -6514 459418 -6278 459654
rect -6514 459098 -6278 459334
rect -6514 423418 -6278 423654
rect -6514 423098 -6278 423334
rect -6514 387418 -6278 387654
rect -6514 387098 -6278 387334
rect -6514 351418 -6278 351654
rect -6514 351098 -6278 351334
rect -6514 315418 -6278 315654
rect -6514 315098 -6278 315334
rect -6514 279418 -6278 279654
rect -6514 279098 -6278 279334
rect -6514 243418 -6278 243654
rect -6514 243098 -6278 243334
rect -6514 207418 -6278 207654
rect -6514 207098 -6278 207334
rect -6514 171418 -6278 171654
rect -6514 171098 -6278 171334
rect -6514 135418 -6278 135654
rect -6514 135098 -6278 135334
rect -6514 99418 -6278 99654
rect -6514 99098 -6278 99334
rect -6514 63418 -6278 63654
rect -6514 63098 -6278 63334
rect -6514 27418 -6278 27654
rect -6514 27098 -6278 27334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 8186 708362 8422 708598
rect 8186 708042 8422 708278
rect -5574 693418 -5338 693654
rect -5574 693098 -5338 693334
rect -5574 657418 -5338 657654
rect -5574 657098 -5338 657334
rect -5574 621418 -5338 621654
rect -5574 621098 -5338 621334
rect -5574 585418 -5338 585654
rect -5574 585098 -5338 585334
rect -5574 549418 -5338 549654
rect -5574 549098 -5338 549334
rect -5574 513418 -5338 513654
rect -5574 513098 -5338 513334
rect -5574 477418 -5338 477654
rect -5574 477098 -5338 477334
rect -5574 441418 -5338 441654
rect -5574 441098 -5338 441334
rect -5574 405418 -5338 405654
rect -5574 405098 -5338 405334
rect -5574 369418 -5338 369654
rect -5574 369098 -5338 369334
rect -5574 333418 -5338 333654
rect -5574 333098 -5338 333334
rect -5574 297418 -5338 297654
rect -5574 297098 -5338 297334
rect -5574 261418 -5338 261654
rect -5574 261098 -5338 261334
rect -5574 225418 -5338 225654
rect -5574 225098 -5338 225334
rect -5574 189418 -5338 189654
rect -5574 189098 -5338 189334
rect -5574 153418 -5338 153654
rect -5574 153098 -5338 153334
rect -5574 117418 -5338 117654
rect -5574 117098 -5338 117334
rect -5574 81418 -5338 81654
rect -5574 81098 -5338 81334
rect -5574 45418 -5338 45654
rect -5574 45098 -5338 45334
rect -5574 9418 -5338 9654
rect -5574 9098 -5338 9334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 671818 -4398 672054
rect -4634 671498 -4398 671734
rect -4634 635818 -4398 636054
rect -4634 635498 -4398 635734
rect -4634 599818 -4398 600054
rect -4634 599498 -4398 599734
rect -4634 563818 -4398 564054
rect -4634 563498 -4398 563734
rect -4634 527818 -4398 528054
rect -4634 527498 -4398 527734
rect -4634 491818 -4398 492054
rect -4634 491498 -4398 491734
rect -4634 455818 -4398 456054
rect -4634 455498 -4398 455734
rect -4634 419818 -4398 420054
rect -4634 419498 -4398 419734
rect -4634 383818 -4398 384054
rect -4634 383498 -4398 383734
rect -4634 347818 -4398 348054
rect -4634 347498 -4398 347734
rect -4634 311818 -4398 312054
rect -4634 311498 -4398 311734
rect -4634 275818 -4398 276054
rect -4634 275498 -4398 275734
rect -4634 239818 -4398 240054
rect -4634 239498 -4398 239734
rect -4634 203818 -4398 204054
rect -4634 203498 -4398 203734
rect -4634 167818 -4398 168054
rect -4634 167498 -4398 167734
rect -4634 131818 -4398 132054
rect -4634 131498 -4398 131734
rect -4634 95818 -4398 96054
rect -4634 95498 -4398 95734
rect -4634 59818 -4398 60054
rect -4634 59498 -4398 59734
rect -4634 23818 -4398 24054
rect -4634 23498 -4398 23734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 4586 706482 4822 706718
rect 4586 706162 4822 706398
rect -3694 689818 -3458 690054
rect -3694 689498 -3458 689734
rect -3694 653818 -3458 654054
rect -3694 653498 -3458 653734
rect -3694 617818 -3458 618054
rect -3694 617498 -3458 617734
rect -3694 581818 -3458 582054
rect -3694 581498 -3458 581734
rect -3694 545818 -3458 546054
rect -3694 545498 -3458 545734
rect -3694 509818 -3458 510054
rect -3694 509498 -3458 509734
rect -3694 473818 -3458 474054
rect -3694 473498 -3458 473734
rect -3694 437818 -3458 438054
rect -3694 437498 -3458 437734
rect -3694 401818 -3458 402054
rect -3694 401498 -3458 401734
rect -3694 365818 -3458 366054
rect -3694 365498 -3458 365734
rect -3694 329818 -3458 330054
rect -3694 329498 -3458 329734
rect -3694 293818 -3458 294054
rect -3694 293498 -3458 293734
rect -3694 257818 -3458 258054
rect -3694 257498 -3458 257734
rect -3694 221818 -3458 222054
rect -3694 221498 -3458 221734
rect -3694 185818 -3458 186054
rect -3694 185498 -3458 185734
rect -3694 149818 -3458 150054
rect -3694 149498 -3458 149734
rect -3694 113818 -3458 114054
rect -3694 113498 -3458 113734
rect -3694 77818 -3458 78054
rect -3694 77498 -3458 77734
rect -3694 41818 -3458 42054
rect -3694 41498 -3458 41734
rect -3694 5818 -3458 6054
rect -3694 5498 -3458 5734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 4586 -2462 4822 -2226
rect 4586 -2782 4822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 8186 -4342 8422 -4106
rect 8186 -4662 8422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 29786 711182 30022 711418
rect 29786 710862 30022 711098
rect 26186 709302 26422 709538
rect 26186 708982 26422 709218
rect 22586 707422 22822 707658
rect 22586 707102 22822 707338
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3402 22822 -3166
rect 22586 -3722 22822 -3486
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5282 26422 -5046
rect 26186 -5602 26422 -5366
rect 47786 710242 48022 710478
rect 47786 709922 48022 710158
rect 44186 708362 44422 708598
rect 44186 708042 44422 708278
rect 40586 706482 40822 706718
rect 40586 706162 40822 706398
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6222 12022 -5986
rect 11786 -6542 12022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2462 40822 -2226
rect 40586 -2782 40822 -2546
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4342 44422 -4106
rect 44186 -4662 44422 -4426
rect 65786 711182 66022 711418
rect 65786 710862 66022 711098
rect 62186 709302 62422 709538
rect 62186 708982 62422 709218
rect 58586 707422 58822 707658
rect 58586 707102 58822 707338
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7162 30022 -6926
rect 29786 -7482 30022 -7246
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3402 58822 -3166
rect 58586 -3722 58822 -3486
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5282 62422 -5046
rect 62186 -5602 62422 -5366
rect 83786 710242 84022 710478
rect 83786 709922 84022 710158
rect 80186 708362 80422 708598
rect 80186 708042 80422 708278
rect 76586 706482 76822 706718
rect 76586 706162 76822 706398
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 101786 711182 102022 711418
rect 101786 710862 102022 711098
rect 98186 709302 98422 709538
rect 98186 708982 98422 709218
rect 94586 707422 94822 707658
rect 94586 707102 94822 707338
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 119786 710242 120022 710478
rect 119786 709922 120022 710158
rect 116186 708362 116422 708598
rect 116186 708042 116422 708278
rect 112586 706482 112822 706718
rect 112586 706162 112822 706398
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 91571 542218 91807 542454
rect 91571 541898 91807 542134
rect 96155 524218 96391 524454
rect 96155 523898 96391 524134
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 137786 711182 138022 711418
rect 137786 710862 138022 711098
rect 134186 709302 134422 709538
rect 134186 708982 134422 709218
rect 130586 707422 130822 707658
rect 130586 707102 130822 707338
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 91610 380218 91846 380454
rect 91610 379898 91846 380134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 76250 362218 76486 362454
rect 76250 361898 76486 362134
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 91610 344218 91846 344454
rect 91610 343898 91846 344134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6222 48022 -5986
rect 47786 -6542 48022 -6306
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2462 76822 -2226
rect 76586 -2782 76822 -2546
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4342 80422 -4106
rect 80186 -4662 80422 -4426
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7162 66022 -6926
rect 65786 -7482 66022 -7246
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3402 94822 -3166
rect 94586 -3722 94822 -3486
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5282 98422 -5046
rect 98186 -5602 98422 -5366
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6222 84022 -5986
rect 83786 -6542 84022 -6306
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2462 112822 -2226
rect 112586 -2782 112822 -2546
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4342 116422 -4106
rect 116186 -4662 116422 -4426
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7162 102022 -6926
rect 101786 -7482 102022 -7246
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 155786 710242 156022 710478
rect 155786 709922 156022 710158
rect 152186 708362 152422 708598
rect 152186 708042 152422 708278
rect 148586 706482 148822 706718
rect 148586 706162 148822 706398
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 173786 711182 174022 711418
rect 173786 710862 174022 711098
rect 170186 709302 170422 709538
rect 170186 708982 170422 709218
rect 166586 707422 166822 707658
rect 166586 707102 166822 707338
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 155786 409018 156022 409254
rect 155786 408698 156022 408934
rect 155786 373018 156022 373254
rect 155786 372698 156022 372934
rect 155786 337018 156022 337254
rect 155786 336698 156022 336934
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 166586 383818 166822 384054
rect 166586 383498 166822 383734
rect 166586 347818 166822 348054
rect 166586 347498 166822 347734
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 170186 387418 170422 387654
rect 170186 387098 170422 387334
rect 170186 351418 170422 351654
rect 170186 351098 170422 351334
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 191786 710242 192022 710478
rect 191786 709922 192022 710158
rect 188186 708362 188422 708598
rect 188186 708042 188422 708278
rect 184586 706482 184822 706718
rect 184586 706162 184822 706398
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 173786 391018 174022 391254
rect 173786 390698 174022 390934
rect 173786 355018 174022 355254
rect 173786 354698 174022 354934
rect 173786 319018 174022 319254
rect 173786 318698 174022 318934
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 184586 401818 184822 402054
rect 184586 401498 184822 401734
rect 184586 365818 184822 366054
rect 184586 365498 184822 365734
rect 184586 329818 184822 330054
rect 184586 329498 184822 329734
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 188186 405418 188422 405654
rect 188186 405098 188422 405334
rect 188186 369418 188422 369654
rect 188186 369098 188422 369334
rect 188186 333418 188422 333654
rect 188186 333098 188422 333334
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 209786 711182 210022 711418
rect 209786 710862 210022 711098
rect 206186 709302 206422 709538
rect 206186 708982 206422 709218
rect 202586 707422 202822 707658
rect 202586 707102 202822 707338
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 191786 409018 192022 409254
rect 191786 408698 192022 408934
rect 191786 373018 192022 373254
rect 191786 372698 192022 372934
rect 191786 337018 192022 337254
rect 191786 336698 192022 336934
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 227786 710242 228022 710478
rect 227786 709922 228022 710158
rect 224186 708362 224422 708598
rect 224186 708042 224422 708278
rect 220586 706482 220822 706718
rect 220586 706162 220822 706398
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 203951 542218 204187 542454
rect 203951 541898 204187 542134
rect 206917 524218 207153 524454
rect 206917 523898 207153 524134
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 245786 711182 246022 711418
rect 245786 710862 246022 711098
rect 242186 709302 242422 709538
rect 242186 708982 242422 709218
rect 238586 707422 238822 707658
rect 238586 707102 238822 707338
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 238586 419818 238822 420054
rect 238586 419498 238822 419734
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 242186 423418 242422 423654
rect 242186 423098 242422 423334
rect 263786 710242 264022 710478
rect 263786 709922 264022 710158
rect 260186 708362 260422 708598
rect 260186 708042 260422 708278
rect 256586 706482 256822 706718
rect 256586 706162 256822 706398
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 260186 477418 260422 477654
rect 260186 477098 260422 477334
rect 260186 441418 260422 441654
rect 260186 441098 260422 441334
rect 281786 711182 282022 711418
rect 281786 710862 282022 711098
rect 278186 709302 278422 709538
rect 278186 708982 278422 709218
rect 274586 707422 274822 707658
rect 274586 707102 274822 707338
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 263786 481018 264022 481254
rect 263786 480698 264022 480934
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 204250 398218 204486 398454
rect 204250 397898 204486 398134
rect 219610 380218 219846 380454
rect 219610 379898 219846 380134
rect 204250 362218 204486 362454
rect 204250 361898 204486 362134
rect 219610 344218 219846 344454
rect 219610 343898 219846 344134
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 209786 319018 210022 319254
rect 209786 318698 210022 318934
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 220586 329818 220822 330054
rect 220586 329498 220822 329734
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 224186 333418 224422 333654
rect 224186 333098 224422 333334
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 227786 337018 228022 337254
rect 227786 336698 228022 336934
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 245786 319018 246022 319254
rect 245786 318698 246022 318934
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 256586 329818 256822 330054
rect 256586 329498 256822 329734
rect 260186 333418 260422 333654
rect 260186 333098 260422 333334
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 263786 337018 264022 337254
rect 263786 336698 264022 336934
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 270986 344218 271222 344454
rect 270986 343898 271222 344134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 274586 419818 274822 420054
rect 274586 419498 274822 419734
rect 274586 383818 274822 384054
rect 274586 383498 274822 383734
rect 274586 347818 274822 348054
rect 274586 347498 274822 347734
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 278186 459418 278422 459654
rect 278186 459098 278422 459334
rect 278186 423418 278422 423654
rect 278186 423098 278422 423334
rect 278186 387418 278422 387654
rect 278186 387098 278422 387334
rect 278186 351418 278422 351654
rect 278186 351098 278422 351334
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 299786 710242 300022 710478
rect 299786 709922 300022 710158
rect 296186 708362 296422 708598
rect 296186 708042 296422 708278
rect 292586 706482 292822 706718
rect 292586 706162 292822 706398
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 281786 463018 282022 463254
rect 281786 462698 282022 462934
rect 281786 427018 282022 427254
rect 281786 426698 282022 426934
rect 281786 391018 282022 391254
rect 281786 390698 282022 390934
rect 281786 355018 282022 355254
rect 281786 354698 282022 354934
rect 281786 319018 282022 319254
rect 281786 318698 282022 318934
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 317786 711182 318022 711418
rect 317786 710862 318022 711098
rect 314186 709302 314422 709538
rect 314186 708982 314422 709218
rect 310586 707422 310822 707658
rect 310586 707102 310822 707338
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 335786 710242 336022 710478
rect 335786 709922 336022 710158
rect 332186 708362 332422 708598
rect 332186 708042 332422 708278
rect 328586 706482 328822 706718
rect 328586 706162 328822 706398
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 353786 711182 354022 711418
rect 353786 710862 354022 711098
rect 350186 709302 350422 709538
rect 350186 708982 350422 709218
rect 346586 707422 346822 707658
rect 346586 707102 346822 707338
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 371786 710242 372022 710478
rect 371786 709922 372022 710158
rect 368186 708362 368422 708598
rect 368186 708042 368422 708278
rect 364586 706482 364822 706718
rect 364586 706162 364822 706398
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 389786 711182 390022 711418
rect 389786 710862 390022 711098
rect 386186 709302 386422 709538
rect 386186 708982 386422 709218
rect 382586 707422 382822 707658
rect 382586 707102 382822 707338
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 319610 560218 319846 560454
rect 319610 559898 319846 560134
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 304250 542218 304486 542454
rect 304250 541898 304486 542134
rect 319610 524218 319846 524454
rect 319610 523898 319846 524134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 304250 506218 304486 506454
rect 304250 505898 304486 506134
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 346586 383818 346822 384054
rect 346586 383498 346822 383734
rect 346586 347818 346822 348054
rect 346586 347498 346822 347734
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 350186 387418 350422 387654
rect 350186 387098 350422 387334
rect 350186 351418 350422 351654
rect 350186 351098 350422 351334
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 353786 391018 354022 391254
rect 353786 390698 354022 390934
rect 353786 355018 354022 355254
rect 353786 354698 354022 354934
rect 353786 319018 354022 319254
rect 353786 318698 354022 318934
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 364586 401818 364822 402054
rect 364586 401498 364822 401734
rect 364586 365818 364822 366054
rect 364586 365498 364822 365734
rect 364586 329818 364822 330054
rect 364586 329498 364822 329734
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 368186 405418 368422 405654
rect 368186 405098 368422 405334
rect 368186 369418 368422 369654
rect 368186 369098 368422 369334
rect 368186 333418 368422 333654
rect 368186 333098 368422 333334
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 371786 409018 372022 409254
rect 371786 408698 372022 408934
rect 371786 373018 372022 373254
rect 371786 372698 372022 372934
rect 371786 337018 372022 337254
rect 371786 336698 372022 336934
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 382586 383818 382822 384054
rect 382586 383498 382822 383734
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 386186 387418 386422 387654
rect 386186 387098 386422 387334
rect 407786 710242 408022 710478
rect 407786 709922 408022 710158
rect 404186 708362 404422 708598
rect 404186 708042 404422 708278
rect 400586 706482 400822 706718
rect 400586 706162 400822 706398
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 389786 391018 390022 391254
rect 389786 390698 390022 390934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 425786 711182 426022 711418
rect 425786 710862 426022 711098
rect 422186 709302 422422 709538
rect 422186 708982 422422 709218
rect 418586 707422 418822 707658
rect 418586 707102 418822 707338
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 394646 380218 394882 380454
rect 394646 379898 394882 380134
rect 389816 362218 390052 362454
rect 389816 361898 390052 362134
rect 382586 347818 382822 348054
rect 382586 347498 382822 347734
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 389786 319018 390022 319254
rect 389786 318698 390022 318934
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 443786 710242 444022 710478
rect 443786 709922 444022 710158
rect 440186 708362 440422 708598
rect 440186 708042 440422 708278
rect 436586 706482 436822 706718
rect 436586 706162 436822 706398
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 138250 182218 138486 182454
rect 138250 181898 138486 182134
rect 153610 164218 153846 164454
rect 153610 163898 153846 164134
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 138250 146218 138486 146454
rect 138250 145898 138486 146134
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 153610 128218 153846 128454
rect 153610 127898 153846 128134
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3402 130822 -3166
rect 130586 -3722 130822 -3486
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5282 134422 -5046
rect 134186 -5602 134422 -5366
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6222 120022 -5986
rect 119786 -6542 120022 -6306
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2462 148822 -2226
rect 148586 -2782 148822 -2546
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4342 152422 -4106
rect 152186 -4662 152422 -4426
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7162 138022 -6926
rect 137786 -7482 138022 -7246
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3402 166822 -3166
rect 166586 -3722 166822 -3486
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5282 170422 -5046
rect 170186 -5602 170422 -5366
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6222 156022 -5986
rect 155786 -6542 156022 -6306
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2462 184822 -2226
rect 184586 -2782 184822 -2546
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4342 188422 -4106
rect 188186 -4662 188422 -4426
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7162 174022 -6926
rect 173786 -7482 174022 -7246
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3402 202822 -3166
rect 202586 -3722 202822 -3486
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5282 206422 -5046
rect 206186 -5602 206422 -5366
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6222 192022 -5986
rect 191786 -6542 192022 -6306
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2462 220822 -2226
rect 220586 -2782 220822 -2546
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4342 224422 -4106
rect 224186 -4662 224422 -4426
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7162 210022 -6926
rect 209786 -7482 210022 -7246
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3402 238822 -3166
rect 238586 -3722 238822 -3486
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5282 242422 -5046
rect 242186 -5602 242422 -5366
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6222 228022 -5986
rect 227786 -6542 228022 -6306
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2462 256822 -2226
rect 256586 -2782 256822 -2546
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4342 260422 -4106
rect 260186 -4662 260422 -4426
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7162 246022 -6926
rect 245786 -7482 246022 -7246
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3402 274822 -3166
rect 274586 -3722 274822 -3486
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5282 278422 -5046
rect 278186 -5602 278422 -5366
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6222 264022 -5986
rect 263786 -6542 264022 -6306
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2462 292822 -2226
rect 292586 -2782 292822 -2546
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4342 296422 -4106
rect 296186 -4662 296422 -4426
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7162 282022 -6926
rect 281786 -7482 282022 -7246
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3402 310822 -3166
rect 310586 -3722 310822 -3486
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5282 314422 -5046
rect 314186 -5602 314422 -5366
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6222 300022 -5986
rect 299786 -6542 300022 -6306
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2462 328822 -2226
rect 328586 -2782 328822 -2546
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4342 332422 -4106
rect 332186 -4662 332422 -4426
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7162 318022 -6926
rect 317786 -7482 318022 -7246
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3402 346822 -3166
rect 346586 -3722 346822 -3486
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5282 350422 -5046
rect 350186 -5602 350422 -5366
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6222 336022 -5986
rect 335786 -6542 336022 -6306
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2462 364822 -2226
rect 364586 -2782 364822 -2546
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4342 368422 -4106
rect 368186 -4662 368422 -4426
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7162 354022 -6926
rect 353786 -7482 354022 -7246
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3402 382822 -3166
rect 382586 -3722 382822 -3486
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5282 386422 -5046
rect 386186 -5602 386422 -5366
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6222 372022 -5986
rect 371786 -6542 372022 -6306
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2462 400822 -2226
rect 400586 -2782 400822 -2546
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4342 404422 -4106
rect 404186 -4662 404422 -4426
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7162 390022 -6926
rect 389786 -7482 390022 -7246
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3402 418822 -3166
rect 418586 -3722 418822 -3486
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5282 422422 -5046
rect 422186 -5602 422422 -5366
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6222 408022 -5986
rect 407786 -6542 408022 -6306
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2462 436822 -2226
rect 436586 -2782 436822 -2546
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4342 440422 -4106
rect 440186 -4662 440422 -4426
rect 461786 711182 462022 711418
rect 461786 710862 462022 711098
rect 458186 709302 458422 709538
rect 458186 708982 458422 709218
rect 454586 707422 454822 707658
rect 454586 707102 454822 707338
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7162 426022 -6926
rect 425786 -7482 426022 -7246
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3402 454822 -3166
rect 454586 -3722 454822 -3486
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 479786 710242 480022 710478
rect 479786 709922 480022 710158
rect 476186 708362 476422 708598
rect 476186 708042 476422 708278
rect 472586 706482 472822 706718
rect 472586 706162 472822 706398
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 497786 711182 498022 711418
rect 497786 710862 498022 711098
rect 494186 709302 494422 709538
rect 494186 708982 494422 709218
rect 490586 707422 490822 707658
rect 490586 707102 490822 707338
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 515786 710242 516022 710478
rect 515786 709922 516022 710158
rect 512186 708362 512422 708598
rect 512186 708042 512422 708278
rect 508586 706482 508822 706718
rect 508586 706162 508822 706398
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 485480 542218 485716 542454
rect 485480 541898 485716 542134
rect 490540 524218 490776 524454
rect 490540 523898 490776 524134
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 479610 380218 479846 380454
rect 479610 379898 479846 380134
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 464250 362218 464486 362454
rect 464250 361898 464486 362134
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 479610 344218 479846 344454
rect 479610 343898 479846 344134
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5282 458422 -5046
rect 458186 -5602 458422 -5366
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6222 444022 -5986
rect 443786 -6542 444022 -6306
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2462 472822 -2226
rect 472586 -2782 472822 -2546
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4342 476422 -4106
rect 476186 -4662 476422 -4426
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7162 462022 -6926
rect 461786 -7482 462022 -7246
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3402 490822 -3166
rect 490586 -3722 490822 -3486
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5282 494422 -5046
rect 494186 -5602 494422 -5366
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6222 480022 -5986
rect 479786 -6542 480022 -6306
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2462 508822 -2226
rect 508586 -2782 508822 -2546
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4342 512422 -4106
rect 512186 -4662 512422 -4426
rect 533786 711182 534022 711418
rect 533786 710862 534022 711098
rect 530186 709302 530422 709538
rect 530186 708982 530422 709218
rect 526586 707422 526822 707658
rect 526586 707102 526822 707338
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7162 498022 -6926
rect 497786 -7482 498022 -7246
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3402 526822 -3166
rect 526586 -3722 526822 -3486
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5282 530422 -5046
rect 530186 -5602 530422 -5366
rect 551786 710242 552022 710478
rect 551786 709922 552022 710158
rect 548186 708362 548422 708598
rect 548186 708042 548422 708278
rect 544586 706482 544822 706718
rect 544586 706162 544822 706398
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6222 516022 -5986
rect 515786 -6542 516022 -6306
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2462 544822 -2226
rect 544586 -2782 544822 -2546
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4342 548422 -4106
rect 548186 -4662 548422 -4426
rect 569786 711182 570022 711418
rect 569786 710862 570022 711098
rect 566186 709302 566422 709538
rect 566186 708982 566422 709218
rect 562586 707422 562822 707658
rect 562586 707102 562822 707338
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7162 534022 -6926
rect 533786 -7482 534022 -7246
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3402 562822 -3166
rect 562586 -3722 562822 -3486
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5282 566422 -5046
rect 566186 -5602 566422 -5366
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 580586 706482 580822 706718
rect 580586 706162 580822 706398
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6222 552022 -5986
rect 551786 -6542 552022 -6306
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 689818 587618 690054
rect 587382 689498 587618 689734
rect 587382 653818 587618 654054
rect 587382 653498 587618 653734
rect 587382 617818 587618 618054
rect 587382 617498 587618 617734
rect 587382 581818 587618 582054
rect 587382 581498 587618 581734
rect 587382 545818 587618 546054
rect 587382 545498 587618 545734
rect 587382 509818 587618 510054
rect 587382 509498 587618 509734
rect 587382 473818 587618 474054
rect 587382 473498 587618 473734
rect 587382 437818 587618 438054
rect 587382 437498 587618 437734
rect 587382 401818 587618 402054
rect 587382 401498 587618 401734
rect 587382 365818 587618 366054
rect 587382 365498 587618 365734
rect 587382 329818 587618 330054
rect 587382 329498 587618 329734
rect 587382 293818 587618 294054
rect 587382 293498 587618 293734
rect 587382 257818 587618 258054
rect 587382 257498 587618 257734
rect 587382 221818 587618 222054
rect 587382 221498 587618 221734
rect 587382 185818 587618 186054
rect 587382 185498 587618 185734
rect 587382 149818 587618 150054
rect 587382 149498 587618 149734
rect 587382 113818 587618 114054
rect 587382 113498 587618 113734
rect 587382 77818 587618 78054
rect 587382 77498 587618 77734
rect 587382 41818 587618 42054
rect 587382 41498 587618 41734
rect 587382 5818 587618 6054
rect 587382 5498 587618 5734
rect 580586 -2462 580822 -2226
rect 580586 -2782 580822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 671818 588558 672054
rect 588322 671498 588558 671734
rect 588322 635818 588558 636054
rect 588322 635498 588558 635734
rect 588322 599818 588558 600054
rect 588322 599498 588558 599734
rect 588322 563818 588558 564054
rect 588322 563498 588558 563734
rect 588322 527818 588558 528054
rect 588322 527498 588558 527734
rect 588322 491818 588558 492054
rect 588322 491498 588558 491734
rect 588322 455818 588558 456054
rect 588322 455498 588558 455734
rect 588322 419818 588558 420054
rect 588322 419498 588558 419734
rect 588322 383818 588558 384054
rect 588322 383498 588558 383734
rect 588322 347818 588558 348054
rect 588322 347498 588558 347734
rect 588322 311818 588558 312054
rect 588322 311498 588558 311734
rect 588322 275818 588558 276054
rect 588322 275498 588558 275734
rect 588322 239818 588558 240054
rect 588322 239498 588558 239734
rect 588322 203818 588558 204054
rect 588322 203498 588558 203734
rect 588322 167818 588558 168054
rect 588322 167498 588558 167734
rect 588322 131818 588558 132054
rect 588322 131498 588558 131734
rect 588322 95818 588558 96054
rect 588322 95498 588558 95734
rect 588322 59818 588558 60054
rect 588322 59498 588558 59734
rect 588322 23818 588558 24054
rect 588322 23498 588558 23734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 693418 589498 693654
rect 589262 693098 589498 693334
rect 589262 657418 589498 657654
rect 589262 657098 589498 657334
rect 589262 621418 589498 621654
rect 589262 621098 589498 621334
rect 589262 585418 589498 585654
rect 589262 585098 589498 585334
rect 589262 549418 589498 549654
rect 589262 549098 589498 549334
rect 589262 513418 589498 513654
rect 589262 513098 589498 513334
rect 589262 477418 589498 477654
rect 589262 477098 589498 477334
rect 589262 441418 589498 441654
rect 589262 441098 589498 441334
rect 589262 405418 589498 405654
rect 589262 405098 589498 405334
rect 589262 369418 589498 369654
rect 589262 369098 589498 369334
rect 589262 333418 589498 333654
rect 589262 333098 589498 333334
rect 589262 297418 589498 297654
rect 589262 297098 589498 297334
rect 589262 261418 589498 261654
rect 589262 261098 589498 261334
rect 589262 225418 589498 225654
rect 589262 225098 589498 225334
rect 589262 189418 589498 189654
rect 589262 189098 589498 189334
rect 589262 153418 589498 153654
rect 589262 153098 589498 153334
rect 589262 117418 589498 117654
rect 589262 117098 589498 117334
rect 589262 81418 589498 81654
rect 589262 81098 589498 81334
rect 589262 45418 589498 45654
rect 589262 45098 589498 45334
rect 589262 9418 589498 9654
rect 589262 9098 589498 9334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 675418 590438 675654
rect 590202 675098 590438 675334
rect 590202 639418 590438 639654
rect 590202 639098 590438 639334
rect 590202 603418 590438 603654
rect 590202 603098 590438 603334
rect 590202 567418 590438 567654
rect 590202 567098 590438 567334
rect 590202 531418 590438 531654
rect 590202 531098 590438 531334
rect 590202 495418 590438 495654
rect 590202 495098 590438 495334
rect 590202 459418 590438 459654
rect 590202 459098 590438 459334
rect 590202 423418 590438 423654
rect 590202 423098 590438 423334
rect 590202 387418 590438 387654
rect 590202 387098 590438 387334
rect 590202 351418 590438 351654
rect 590202 351098 590438 351334
rect 590202 315418 590438 315654
rect 590202 315098 590438 315334
rect 590202 279418 590438 279654
rect 590202 279098 590438 279334
rect 590202 243418 590438 243654
rect 590202 243098 590438 243334
rect 590202 207418 590438 207654
rect 590202 207098 590438 207334
rect 590202 171418 590438 171654
rect 590202 171098 590438 171334
rect 590202 135418 590438 135654
rect 590202 135098 590438 135334
rect 590202 99418 590438 99654
rect 590202 99098 590438 99334
rect 590202 63418 590438 63654
rect 590202 63098 590438 63334
rect 590202 27418 590438 27654
rect 590202 27098 590438 27334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 697018 591378 697254
rect 591142 696698 591378 696934
rect 591142 661018 591378 661254
rect 591142 660698 591378 660934
rect 591142 625018 591378 625254
rect 591142 624698 591378 624934
rect 591142 589018 591378 589254
rect 591142 588698 591378 588934
rect 591142 553018 591378 553254
rect 591142 552698 591378 552934
rect 591142 517018 591378 517254
rect 591142 516698 591378 516934
rect 591142 481018 591378 481254
rect 591142 480698 591378 480934
rect 591142 445018 591378 445254
rect 591142 444698 591378 444934
rect 591142 409018 591378 409254
rect 591142 408698 591378 408934
rect 591142 373018 591378 373254
rect 591142 372698 591378 372934
rect 591142 337018 591378 337254
rect 591142 336698 591378 336934
rect 591142 301018 591378 301254
rect 591142 300698 591378 300934
rect 591142 265018 591378 265254
rect 591142 264698 591378 264934
rect 591142 229018 591378 229254
rect 591142 228698 591378 228934
rect 591142 193018 591378 193254
rect 591142 192698 591378 192934
rect 591142 157018 591378 157254
rect 591142 156698 591378 156934
rect 591142 121018 591378 121254
rect 591142 120698 591378 120934
rect 591142 85018 591378 85254
rect 591142 84698 591378 84934
rect 591142 49018 591378 49254
rect 591142 48698 591378 48934
rect 591142 13018 591378 13254
rect 591142 12698 591378 12934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 679018 592318 679254
rect 592082 678698 592318 678934
rect 592082 643018 592318 643254
rect 592082 642698 592318 642934
rect 592082 607018 592318 607254
rect 592082 606698 592318 606934
rect 592082 571018 592318 571254
rect 592082 570698 592318 570934
rect 592082 535018 592318 535254
rect 592082 534698 592318 534934
rect 592082 499018 592318 499254
rect 592082 498698 592318 498934
rect 592082 463018 592318 463254
rect 592082 462698 592318 462934
rect 592082 427018 592318 427254
rect 592082 426698 592318 426934
rect 592082 391018 592318 391254
rect 592082 390698 592318 390934
rect 592082 355018 592318 355254
rect 592082 354698 592318 354934
rect 592082 319018 592318 319254
rect 592082 318698 592318 318934
rect 592082 283018 592318 283254
rect 592082 282698 592318 282934
rect 592082 247018 592318 247254
rect 592082 246698 592318 246934
rect 592082 211018 592318 211254
rect 592082 210698 592318 210934
rect 592082 175018 592318 175254
rect 592082 174698 592318 174934
rect 592082 139018 592318 139254
rect 592082 138698 592318 138934
rect 592082 103018 592318 103254
rect 592082 102698 592318 102934
rect 592082 67018 592318 67254
rect 592082 66698 592318 66934
rect 592082 31018 592318 31254
rect 592082 30698 592318 30934
rect 569786 -7162 570022 -6926
rect 569786 -7482 570022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 29786 711418
rect 30022 711182 65786 711418
rect 66022 711182 101786 711418
rect 102022 711182 137786 711418
rect 138022 711182 173786 711418
rect 174022 711182 209786 711418
rect 210022 711182 245786 711418
rect 246022 711182 281786 711418
rect 282022 711182 317786 711418
rect 318022 711182 353786 711418
rect 354022 711182 389786 711418
rect 390022 711182 425786 711418
rect 426022 711182 461786 711418
rect 462022 711182 497786 711418
rect 498022 711182 533786 711418
rect 534022 711182 569786 711418
rect 570022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 29786 711098
rect 30022 710862 65786 711098
rect 66022 710862 101786 711098
rect 102022 710862 137786 711098
rect 138022 710862 173786 711098
rect 174022 710862 209786 711098
rect 210022 710862 245786 711098
rect 246022 710862 281786 711098
rect 282022 710862 317786 711098
rect 318022 710862 353786 711098
rect 354022 710862 389786 711098
rect 390022 710862 425786 711098
rect 426022 710862 461786 711098
rect 462022 710862 497786 711098
rect 498022 710862 533786 711098
rect 534022 710862 569786 711098
rect 570022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 11786 710478
rect 12022 710242 47786 710478
rect 48022 710242 83786 710478
rect 84022 710242 119786 710478
rect 120022 710242 155786 710478
rect 156022 710242 191786 710478
rect 192022 710242 227786 710478
rect 228022 710242 263786 710478
rect 264022 710242 299786 710478
rect 300022 710242 335786 710478
rect 336022 710242 371786 710478
rect 372022 710242 407786 710478
rect 408022 710242 443786 710478
rect 444022 710242 479786 710478
rect 480022 710242 515786 710478
rect 516022 710242 551786 710478
rect 552022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 11786 710158
rect 12022 709922 47786 710158
rect 48022 709922 83786 710158
rect 84022 709922 119786 710158
rect 120022 709922 155786 710158
rect 156022 709922 191786 710158
rect 192022 709922 227786 710158
rect 228022 709922 263786 710158
rect 264022 709922 299786 710158
rect 300022 709922 335786 710158
rect 336022 709922 371786 710158
rect 372022 709922 407786 710158
rect 408022 709922 443786 710158
rect 444022 709922 479786 710158
rect 480022 709922 515786 710158
rect 516022 709922 551786 710158
rect 552022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 26186 709538
rect 26422 709302 62186 709538
rect 62422 709302 98186 709538
rect 98422 709302 134186 709538
rect 134422 709302 170186 709538
rect 170422 709302 206186 709538
rect 206422 709302 242186 709538
rect 242422 709302 278186 709538
rect 278422 709302 314186 709538
rect 314422 709302 350186 709538
rect 350422 709302 386186 709538
rect 386422 709302 422186 709538
rect 422422 709302 458186 709538
rect 458422 709302 494186 709538
rect 494422 709302 530186 709538
rect 530422 709302 566186 709538
rect 566422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 26186 709218
rect 26422 708982 62186 709218
rect 62422 708982 98186 709218
rect 98422 708982 134186 709218
rect 134422 708982 170186 709218
rect 170422 708982 206186 709218
rect 206422 708982 242186 709218
rect 242422 708982 278186 709218
rect 278422 708982 314186 709218
rect 314422 708982 350186 709218
rect 350422 708982 386186 709218
rect 386422 708982 422186 709218
rect 422422 708982 458186 709218
rect 458422 708982 494186 709218
rect 494422 708982 530186 709218
rect 530422 708982 566186 709218
rect 566422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 8186 708598
rect 8422 708362 44186 708598
rect 44422 708362 80186 708598
rect 80422 708362 116186 708598
rect 116422 708362 152186 708598
rect 152422 708362 188186 708598
rect 188422 708362 224186 708598
rect 224422 708362 260186 708598
rect 260422 708362 296186 708598
rect 296422 708362 332186 708598
rect 332422 708362 368186 708598
rect 368422 708362 404186 708598
rect 404422 708362 440186 708598
rect 440422 708362 476186 708598
rect 476422 708362 512186 708598
rect 512422 708362 548186 708598
rect 548422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 8186 708278
rect 8422 708042 44186 708278
rect 44422 708042 80186 708278
rect 80422 708042 116186 708278
rect 116422 708042 152186 708278
rect 152422 708042 188186 708278
rect 188422 708042 224186 708278
rect 224422 708042 260186 708278
rect 260422 708042 296186 708278
rect 296422 708042 332186 708278
rect 332422 708042 368186 708278
rect 368422 708042 404186 708278
rect 404422 708042 440186 708278
rect 440422 708042 476186 708278
rect 476422 708042 512186 708278
rect 512422 708042 548186 708278
rect 548422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 22586 707658
rect 22822 707422 58586 707658
rect 58822 707422 94586 707658
rect 94822 707422 130586 707658
rect 130822 707422 166586 707658
rect 166822 707422 202586 707658
rect 202822 707422 238586 707658
rect 238822 707422 274586 707658
rect 274822 707422 310586 707658
rect 310822 707422 346586 707658
rect 346822 707422 382586 707658
rect 382822 707422 418586 707658
rect 418822 707422 454586 707658
rect 454822 707422 490586 707658
rect 490822 707422 526586 707658
rect 526822 707422 562586 707658
rect 562822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 22586 707338
rect 22822 707102 58586 707338
rect 58822 707102 94586 707338
rect 94822 707102 130586 707338
rect 130822 707102 166586 707338
rect 166822 707102 202586 707338
rect 202822 707102 238586 707338
rect 238822 707102 274586 707338
rect 274822 707102 310586 707338
rect 310822 707102 346586 707338
rect 346822 707102 382586 707338
rect 382822 707102 418586 707338
rect 418822 707102 454586 707338
rect 454822 707102 490586 707338
rect 490822 707102 526586 707338
rect 526822 707102 562586 707338
rect 562822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 4586 706718
rect 4822 706482 40586 706718
rect 40822 706482 76586 706718
rect 76822 706482 112586 706718
rect 112822 706482 148586 706718
rect 148822 706482 184586 706718
rect 184822 706482 220586 706718
rect 220822 706482 256586 706718
rect 256822 706482 292586 706718
rect 292822 706482 328586 706718
rect 328822 706482 364586 706718
rect 364822 706482 400586 706718
rect 400822 706482 436586 706718
rect 436822 706482 472586 706718
rect 472822 706482 508586 706718
rect 508822 706482 544586 706718
rect 544822 706482 580586 706718
rect 580822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 4586 706398
rect 4822 706162 40586 706398
rect 40822 706162 76586 706398
rect 76822 706162 112586 706398
rect 112822 706162 148586 706398
rect 148822 706162 184586 706398
rect 184822 706162 220586 706398
rect 220822 706162 256586 706398
rect 256822 706162 292586 706398
rect 292822 706162 328586 706398
rect 328822 706162 364586 706398
rect 364822 706162 400586 706398
rect 400822 706162 436586 706398
rect 436822 706162 472586 706398
rect 472822 706162 508586 706398
rect 508822 706162 544586 706398
rect 544822 706162 580586 706398
rect 580822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7636 697276 -7036 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590960 697276 591560 697278
rect -8576 697254 592500 697276
rect -8576 697018 -7454 697254
rect -7218 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591142 697254
rect 591378 697018 592500 697254
rect -8576 696934 592500 697018
rect -8576 696698 -7454 696934
rect -7218 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591142 696934
rect 591378 696698 592500 696934
rect -8576 696676 592500 696698
rect -7636 696674 -7036 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590960 696674 591560 696676
rect -5756 693676 -5156 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589080 693676 589680 693678
rect -6696 693654 590620 693676
rect -6696 693418 -5574 693654
rect -5338 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589262 693654
rect 589498 693418 590620 693654
rect -6696 693334 590620 693418
rect -6696 693098 -5574 693334
rect -5338 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589262 693334
rect 589498 693098 590620 693334
rect -6696 693076 590620 693098
rect -5756 693074 -5156 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589080 693074 589680 693076
rect -3876 690076 -3276 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587200 690076 587800 690078
rect -4816 690054 588740 690076
rect -4816 689818 -3694 690054
rect -3458 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587382 690054
rect 587618 689818 588740 690054
rect -4816 689734 588740 689818
rect -4816 689498 -3694 689734
rect -3458 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587382 689734
rect 587618 689498 588740 689734
rect -4816 689476 588740 689498
rect -3876 689474 -3276 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587200 689474 587800 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8576 679276 -7976 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591900 679276 592500 679278
rect -8576 679254 592500 679276
rect -8576 679018 -8394 679254
rect -8158 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 592082 679254
rect 592318 679018 592500 679254
rect -8576 678934 592500 679018
rect -8576 678698 -8394 678934
rect -8158 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 592082 678934
rect 592318 678698 592500 678934
rect -8576 678676 592500 678698
rect -8576 678674 -7976 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591900 678674 592500 678676
rect -6696 675676 -6096 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 590020 675676 590620 675678
rect -6696 675654 590620 675676
rect -6696 675418 -6514 675654
rect -6278 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590202 675654
rect 590438 675418 590620 675654
rect -6696 675334 590620 675418
rect -6696 675098 -6514 675334
rect -6278 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590202 675334
rect 590438 675098 590620 675334
rect -6696 675076 590620 675098
rect -6696 675074 -6096 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 590020 675074 590620 675076
rect -4816 672076 -4216 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588140 672076 588740 672078
rect -4816 672054 588740 672076
rect -4816 671818 -4634 672054
rect -4398 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588322 672054
rect 588558 671818 588740 672054
rect -4816 671734 588740 671818
rect -4816 671498 -4634 671734
rect -4398 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588322 671734
rect 588558 671498 588740 671734
rect -4816 671476 588740 671498
rect -4816 671474 -4216 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588140 671474 588740 671476
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -7636 661276 -7036 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590960 661276 591560 661278
rect -8576 661254 592500 661276
rect -8576 661018 -7454 661254
rect -7218 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591142 661254
rect 591378 661018 592500 661254
rect -8576 660934 592500 661018
rect -8576 660698 -7454 660934
rect -7218 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591142 660934
rect 591378 660698 592500 660934
rect -8576 660676 592500 660698
rect -7636 660674 -7036 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590960 660674 591560 660676
rect -5756 657676 -5156 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589080 657676 589680 657678
rect -6696 657654 590620 657676
rect -6696 657418 -5574 657654
rect -5338 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589262 657654
rect 589498 657418 590620 657654
rect -6696 657334 590620 657418
rect -6696 657098 -5574 657334
rect -5338 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589262 657334
rect 589498 657098 590620 657334
rect -6696 657076 590620 657098
rect -5756 657074 -5156 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589080 657074 589680 657076
rect -3876 654076 -3276 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587200 654076 587800 654078
rect -4816 654054 588740 654076
rect -4816 653818 -3694 654054
rect -3458 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587382 654054
rect 587618 653818 588740 654054
rect -4816 653734 588740 653818
rect -4816 653498 -3694 653734
rect -3458 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587382 653734
rect 587618 653498 588740 653734
rect -4816 653476 588740 653498
rect -3876 653474 -3276 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587200 653474 587800 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8576 643276 -7976 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591900 643276 592500 643278
rect -8576 643254 592500 643276
rect -8576 643018 -8394 643254
rect -8158 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 592082 643254
rect 592318 643018 592500 643254
rect -8576 642934 592500 643018
rect -8576 642698 -8394 642934
rect -8158 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 592082 642934
rect 592318 642698 592500 642934
rect -8576 642676 592500 642698
rect -8576 642674 -7976 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591900 642674 592500 642676
rect -6696 639676 -6096 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 590020 639676 590620 639678
rect -6696 639654 590620 639676
rect -6696 639418 -6514 639654
rect -6278 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590202 639654
rect 590438 639418 590620 639654
rect -6696 639334 590620 639418
rect -6696 639098 -6514 639334
rect -6278 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590202 639334
rect 590438 639098 590620 639334
rect -6696 639076 590620 639098
rect -6696 639074 -6096 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 590020 639074 590620 639076
rect -4816 636076 -4216 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588140 636076 588740 636078
rect -4816 636054 588740 636076
rect -4816 635818 -4634 636054
rect -4398 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588322 636054
rect 588558 635818 588740 636054
rect -4816 635734 588740 635818
rect -4816 635498 -4634 635734
rect -4398 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588322 635734
rect 588558 635498 588740 635734
rect -4816 635476 588740 635498
rect -4816 635474 -4216 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588140 635474 588740 635476
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -7636 625276 -7036 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590960 625276 591560 625278
rect -8576 625254 592500 625276
rect -8576 625018 -7454 625254
rect -7218 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591142 625254
rect 591378 625018 592500 625254
rect -8576 624934 592500 625018
rect -8576 624698 -7454 624934
rect -7218 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591142 624934
rect 591378 624698 592500 624934
rect -8576 624676 592500 624698
rect -7636 624674 -7036 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590960 624674 591560 624676
rect -5756 621676 -5156 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589080 621676 589680 621678
rect -6696 621654 590620 621676
rect -6696 621418 -5574 621654
rect -5338 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589262 621654
rect 589498 621418 590620 621654
rect -6696 621334 590620 621418
rect -6696 621098 -5574 621334
rect -5338 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589262 621334
rect 589498 621098 590620 621334
rect -6696 621076 590620 621098
rect -5756 621074 -5156 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589080 621074 589680 621076
rect -3876 618076 -3276 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587200 618076 587800 618078
rect -4816 618054 588740 618076
rect -4816 617818 -3694 618054
rect -3458 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587382 618054
rect 587618 617818 588740 618054
rect -4816 617734 588740 617818
rect -4816 617498 -3694 617734
rect -3458 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587382 617734
rect 587618 617498 588740 617734
rect -4816 617476 588740 617498
rect -3876 617474 -3276 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587200 617474 587800 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8576 607276 -7976 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591900 607276 592500 607278
rect -8576 607254 592500 607276
rect -8576 607018 -8394 607254
rect -8158 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 592082 607254
rect 592318 607018 592500 607254
rect -8576 606934 592500 607018
rect -8576 606698 -8394 606934
rect -8158 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 592082 606934
rect 592318 606698 592500 606934
rect -8576 606676 592500 606698
rect -8576 606674 -7976 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591900 606674 592500 606676
rect -6696 603676 -6096 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 590020 603676 590620 603678
rect -6696 603654 590620 603676
rect -6696 603418 -6514 603654
rect -6278 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590202 603654
rect 590438 603418 590620 603654
rect -6696 603334 590620 603418
rect -6696 603098 -6514 603334
rect -6278 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590202 603334
rect 590438 603098 590620 603334
rect -6696 603076 590620 603098
rect -6696 603074 -6096 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 590020 603074 590620 603076
rect -4816 600076 -4216 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588140 600076 588740 600078
rect -4816 600054 588740 600076
rect -4816 599818 -4634 600054
rect -4398 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588322 600054
rect 588558 599818 588740 600054
rect -4816 599734 588740 599818
rect -4816 599498 -4634 599734
rect -4398 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588322 599734
rect 588558 599498 588740 599734
rect -4816 599476 588740 599498
rect -4816 599474 -4216 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588140 599474 588740 599476
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -7636 589276 -7036 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590960 589276 591560 589278
rect -8576 589254 592500 589276
rect -8576 589018 -7454 589254
rect -7218 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591142 589254
rect 591378 589018 592500 589254
rect -8576 588934 592500 589018
rect -8576 588698 -7454 588934
rect -7218 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591142 588934
rect 591378 588698 592500 588934
rect -8576 588676 592500 588698
rect -7636 588674 -7036 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590960 588674 591560 588676
rect -5756 585676 -5156 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589080 585676 589680 585678
rect -6696 585654 590620 585676
rect -6696 585418 -5574 585654
rect -5338 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589262 585654
rect 589498 585418 590620 585654
rect -6696 585334 590620 585418
rect -6696 585098 -5574 585334
rect -5338 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589262 585334
rect 589498 585098 590620 585334
rect -6696 585076 590620 585098
rect -5756 585074 -5156 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589080 585074 589680 585076
rect -3876 582076 -3276 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587200 582076 587800 582078
rect -4816 582054 588740 582076
rect -4816 581818 -3694 582054
rect -3458 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587382 582054
rect 587618 581818 588740 582054
rect -4816 581734 588740 581818
rect -4816 581498 -3694 581734
rect -3458 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587382 581734
rect 587618 581498 588740 581734
rect -4816 581476 588740 581498
rect -3876 581474 -3276 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587200 581474 587800 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8576 571276 -7976 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591900 571276 592500 571278
rect -8576 571254 592500 571276
rect -8576 571018 -8394 571254
rect -8158 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 592082 571254
rect 592318 571018 592500 571254
rect -8576 570934 592500 571018
rect -8576 570698 -8394 570934
rect -8158 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 592082 570934
rect 592318 570698 592500 570934
rect -8576 570676 592500 570698
rect -8576 570674 -7976 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591900 570674 592500 570676
rect -6696 567676 -6096 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 590020 567676 590620 567678
rect -6696 567654 590620 567676
rect -6696 567418 -6514 567654
rect -6278 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590202 567654
rect 590438 567418 590620 567654
rect -6696 567334 590620 567418
rect -6696 567098 -6514 567334
rect -6278 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590202 567334
rect 590438 567098 590620 567334
rect -6696 567076 590620 567098
rect -6696 567074 -6096 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 590020 567074 590620 567076
rect -4816 564076 -4216 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588140 564076 588740 564078
rect -4816 564054 588740 564076
rect -4816 563818 -4634 564054
rect -4398 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588322 564054
rect 588558 563818 588740 564054
rect -4816 563734 588740 563818
rect -4816 563498 -4634 563734
rect -4398 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588322 563734
rect 588558 563498 588740 563734
rect -4816 563476 588740 563498
rect -4816 563474 -4216 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588140 563474 588740 563476
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 319568 560476 319888 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 319610 560454
rect 319846 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 319610 560134
rect 319846 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 319568 559874 319888 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -7636 553276 -7036 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590960 553276 591560 553278
rect -8576 553254 592500 553276
rect -8576 553018 -7454 553254
rect -7218 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591142 553254
rect 591378 553018 592500 553254
rect -8576 552934 592500 553018
rect -8576 552698 -7454 552934
rect -7218 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591142 552934
rect 591378 552698 592500 552934
rect -8576 552676 592500 552698
rect -7636 552674 -7036 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590960 552674 591560 552676
rect -5756 549676 -5156 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589080 549676 589680 549678
rect -6696 549654 590620 549676
rect -6696 549418 -5574 549654
rect -5338 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589262 549654
rect 589498 549418 590620 549654
rect -6696 549334 590620 549418
rect -6696 549098 -5574 549334
rect -5338 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589262 549334
rect 589498 549098 590620 549334
rect -6696 549076 590620 549098
rect -5756 549074 -5156 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589080 549074 589680 549076
rect -3876 546076 -3276 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587200 546076 587800 546078
rect -4816 546054 588740 546076
rect -4816 545818 -3694 546054
rect -3458 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587382 546054
rect 587618 545818 588740 546054
rect -4816 545734 588740 545818
rect -4816 545498 -3694 545734
rect -3458 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587382 545734
rect 587618 545498 588740 545734
rect -4816 545476 588740 545498
rect -3876 545474 -3276 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587200 545474 587800 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 91529 542476 91849 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 203909 542476 204229 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 304208 542476 304528 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 485438 542476 485758 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 91571 542454
rect 91807 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 203951 542454
rect 204187 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 304250 542454
rect 304486 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 485480 542454
rect 485716 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 91571 542134
rect 91807 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 203951 542134
rect 204187 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 304250 542134
rect 304486 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 485480 542134
rect 485716 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 91529 541874 91849 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 203909 541874 204229 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 304208 541874 304528 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 485438 541874 485758 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8576 535276 -7976 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591900 535276 592500 535278
rect -8576 535254 592500 535276
rect -8576 535018 -8394 535254
rect -8158 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 592082 535254
rect 592318 535018 592500 535254
rect -8576 534934 592500 535018
rect -8576 534698 -8394 534934
rect -8158 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 592082 534934
rect 592318 534698 592500 534934
rect -8576 534676 592500 534698
rect -8576 534674 -7976 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591900 534674 592500 534676
rect -6696 531676 -6096 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 590020 531676 590620 531678
rect -6696 531654 590620 531676
rect -6696 531418 -6514 531654
rect -6278 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590202 531654
rect 590438 531418 590620 531654
rect -6696 531334 590620 531418
rect -6696 531098 -6514 531334
rect -6278 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590202 531334
rect 590438 531098 590620 531334
rect -6696 531076 590620 531098
rect -6696 531074 -6096 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 590020 531074 590620 531076
rect -4816 528076 -4216 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588140 528076 588740 528078
rect -4816 528054 588740 528076
rect -4816 527818 -4634 528054
rect -4398 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588322 528054
rect 588558 527818 588740 528054
rect -4816 527734 588740 527818
rect -4816 527498 -4634 527734
rect -4398 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588322 527734
rect 588558 527498 588740 527734
rect -4816 527476 588740 527498
rect -4816 527474 -4216 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588140 527474 588740 527476
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 96113 524476 96433 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 206875 524476 207195 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 319568 524476 319888 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 490498 524476 490818 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 96155 524454
rect 96391 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 206917 524454
rect 207153 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 319610 524454
rect 319846 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 490540 524454
rect 490776 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 96155 524134
rect 96391 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 206917 524134
rect 207153 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 319610 524134
rect 319846 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 490540 524134
rect 490776 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 96113 523874 96433 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 206875 523874 207195 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 319568 523874 319888 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 490498 523874 490818 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586260 523874 586860 523876
rect -7636 517276 -7036 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590960 517276 591560 517278
rect -8576 517254 592500 517276
rect -8576 517018 -7454 517254
rect -7218 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591142 517254
rect 591378 517018 592500 517254
rect -8576 516934 592500 517018
rect -8576 516698 -7454 516934
rect -7218 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591142 516934
rect 591378 516698 592500 516934
rect -8576 516676 592500 516698
rect -7636 516674 -7036 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590960 516674 591560 516676
rect -5756 513676 -5156 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589080 513676 589680 513678
rect -6696 513654 590620 513676
rect -6696 513418 -5574 513654
rect -5338 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589262 513654
rect 589498 513418 590620 513654
rect -6696 513334 590620 513418
rect -6696 513098 -5574 513334
rect -5338 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589262 513334
rect 589498 513098 590620 513334
rect -6696 513076 590620 513098
rect -5756 513074 -5156 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589080 513074 589680 513076
rect -3876 510076 -3276 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587200 510076 587800 510078
rect -4816 510054 588740 510076
rect -4816 509818 -3694 510054
rect -3458 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587382 510054
rect 587618 509818 588740 510054
rect -4816 509734 588740 509818
rect -4816 509498 -3694 509734
rect -3458 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587382 509734
rect 587618 509498 588740 509734
rect -4816 509476 588740 509498
rect -3876 509474 -3276 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587200 509474 587800 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 304208 506476 304528 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 304250 506454
rect 304486 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 304250 506134
rect 304486 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 304208 505874 304528 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8576 499276 -7976 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591900 499276 592500 499278
rect -8576 499254 592500 499276
rect -8576 499018 -8394 499254
rect -8158 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 592082 499254
rect 592318 499018 592500 499254
rect -8576 498934 592500 499018
rect -8576 498698 -8394 498934
rect -8158 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 592082 498934
rect 592318 498698 592500 498934
rect -8576 498676 592500 498698
rect -8576 498674 -7976 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591900 498674 592500 498676
rect -6696 495676 -6096 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 590020 495676 590620 495678
rect -6696 495654 590620 495676
rect -6696 495418 -6514 495654
rect -6278 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590202 495654
rect 590438 495418 590620 495654
rect -6696 495334 590620 495418
rect -6696 495098 -6514 495334
rect -6278 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590202 495334
rect 590438 495098 590620 495334
rect -6696 495076 590620 495098
rect -6696 495074 -6096 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 590020 495074 590620 495076
rect -4816 492076 -4216 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588140 492076 588740 492078
rect -4816 492054 588740 492076
rect -4816 491818 -4634 492054
rect -4398 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588322 492054
rect 588558 491818 588740 492054
rect -4816 491734 588740 491818
rect -4816 491498 -4634 491734
rect -4398 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588322 491734
rect 588558 491498 588740 491734
rect -4816 491476 588740 491498
rect -4816 491474 -4216 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588140 491474 588740 491476
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -7636 481276 -7036 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 263604 481276 264204 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590960 481276 591560 481278
rect -8576 481254 592500 481276
rect -8576 481018 -7454 481254
rect -7218 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 263786 481254
rect 264022 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591142 481254
rect 591378 481018 592500 481254
rect -8576 480934 592500 481018
rect -8576 480698 -7454 480934
rect -7218 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 263786 480934
rect 264022 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591142 480934
rect 591378 480698 592500 480934
rect -8576 480676 592500 480698
rect -7636 480674 -7036 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 263604 480674 264204 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590960 480674 591560 480676
rect -5756 477676 -5156 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 260004 477676 260604 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589080 477676 589680 477678
rect -6696 477654 590620 477676
rect -6696 477418 -5574 477654
rect -5338 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 260186 477654
rect 260422 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589262 477654
rect 589498 477418 590620 477654
rect -6696 477334 590620 477418
rect -6696 477098 -5574 477334
rect -5338 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 260186 477334
rect 260422 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589262 477334
rect 589498 477098 590620 477334
rect -6696 477076 590620 477098
rect -5756 477074 -5156 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 260004 477074 260604 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589080 477074 589680 477076
rect -3876 474076 -3276 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587200 474076 587800 474078
rect -4816 474054 588740 474076
rect -4816 473818 -3694 474054
rect -3458 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587382 474054
rect 587618 473818 588740 474054
rect -4816 473734 588740 473818
rect -4816 473498 -3694 473734
rect -3458 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587382 473734
rect 587618 473498 588740 473734
rect -4816 473476 588740 473498
rect -3876 473474 -3276 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587200 473474 587800 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8576 463276 -7976 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 281604 463276 282204 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591900 463276 592500 463278
rect -8576 463254 592500 463276
rect -8576 463018 -8394 463254
rect -8158 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 281786 463254
rect 282022 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 592082 463254
rect 592318 463018 592500 463254
rect -8576 462934 592500 463018
rect -8576 462698 -8394 462934
rect -8158 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 281786 462934
rect 282022 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 592082 462934
rect 592318 462698 592500 462934
rect -8576 462676 592500 462698
rect -8576 462674 -7976 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 281604 462674 282204 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591900 462674 592500 462676
rect -6696 459676 -6096 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 278004 459676 278604 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 590020 459676 590620 459678
rect -6696 459654 590620 459676
rect -6696 459418 -6514 459654
rect -6278 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 278186 459654
rect 278422 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590202 459654
rect 590438 459418 590620 459654
rect -6696 459334 590620 459418
rect -6696 459098 -6514 459334
rect -6278 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 278186 459334
rect 278422 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590202 459334
rect 590438 459098 590620 459334
rect -6696 459076 590620 459098
rect -6696 459074 -6096 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 278004 459074 278604 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 590020 459074 590620 459076
rect -4816 456076 -4216 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588140 456076 588740 456078
rect -4816 456054 588740 456076
rect -4816 455818 -4634 456054
rect -4398 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588322 456054
rect 588558 455818 588740 456054
rect -4816 455734 588740 455818
rect -4816 455498 -4634 455734
rect -4398 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588322 455734
rect 588558 455498 588740 455734
rect -4816 455476 588740 455498
rect -4816 455474 -4216 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588140 455474 588740 455476
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -7636 445276 -7036 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590960 445276 591560 445278
rect -8576 445254 592500 445276
rect -8576 445018 -7454 445254
rect -7218 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591142 445254
rect 591378 445018 592500 445254
rect -8576 444934 592500 445018
rect -8576 444698 -7454 444934
rect -7218 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591142 444934
rect 591378 444698 592500 444934
rect -8576 444676 592500 444698
rect -7636 444674 -7036 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590960 444674 591560 444676
rect -5756 441676 -5156 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 260004 441676 260604 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589080 441676 589680 441678
rect -6696 441654 590620 441676
rect -6696 441418 -5574 441654
rect -5338 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 260186 441654
rect 260422 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589262 441654
rect 589498 441418 590620 441654
rect -6696 441334 590620 441418
rect -6696 441098 -5574 441334
rect -5338 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 260186 441334
rect 260422 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589262 441334
rect 589498 441098 590620 441334
rect -6696 441076 590620 441098
rect -5756 441074 -5156 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 260004 441074 260604 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589080 441074 589680 441076
rect -3876 438076 -3276 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587200 438076 587800 438078
rect -4816 438054 588740 438076
rect -4816 437818 -3694 438054
rect -3458 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587382 438054
rect 587618 437818 588740 438054
rect -4816 437734 588740 437818
rect -4816 437498 -3694 437734
rect -3458 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587382 437734
rect 587618 437498 588740 437734
rect -4816 437476 588740 437498
rect -3876 437474 -3276 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587200 437474 587800 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8576 427276 -7976 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 281604 427276 282204 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591900 427276 592500 427278
rect -8576 427254 592500 427276
rect -8576 427018 -8394 427254
rect -8158 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 281786 427254
rect 282022 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 592082 427254
rect 592318 427018 592500 427254
rect -8576 426934 592500 427018
rect -8576 426698 -8394 426934
rect -8158 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 281786 426934
rect 282022 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 592082 426934
rect 592318 426698 592500 426934
rect -8576 426676 592500 426698
rect -8576 426674 -7976 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 281604 426674 282204 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591900 426674 592500 426676
rect -6696 423676 -6096 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 278004 423676 278604 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 590020 423676 590620 423678
rect -6696 423654 590620 423676
rect -6696 423418 -6514 423654
rect -6278 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 278186 423654
rect 278422 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590202 423654
rect 590438 423418 590620 423654
rect -6696 423334 590620 423418
rect -6696 423098 -6514 423334
rect -6278 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 278186 423334
rect 278422 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590202 423334
rect 590438 423098 590620 423334
rect -6696 423076 590620 423098
rect -6696 423074 -6096 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 278004 423074 278604 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 590020 423074 590620 423076
rect -4816 420076 -4216 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 238404 420076 239004 420078
rect 274404 420076 275004 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588140 420076 588740 420078
rect -4816 420054 588740 420076
rect -4816 419818 -4634 420054
rect -4398 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 238586 420054
rect 238822 419818 274586 420054
rect 274822 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588322 420054
rect 588558 419818 588740 420054
rect -4816 419734 588740 419818
rect -4816 419498 -4634 419734
rect -4398 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 238586 419734
rect 238822 419498 274586 419734
rect 274822 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588322 419734
rect 588558 419498 588740 419734
rect -4816 419476 588740 419498
rect -4816 419474 -4216 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 238404 419474 239004 419476
rect 274404 419474 275004 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588140 419474 588740 419476
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect -7636 409276 -7036 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 155604 409276 156204 409278
rect 191604 409276 192204 409278
rect 299604 409276 300204 409278
rect 335604 409276 336204 409278
rect 371604 409276 372204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590960 409276 591560 409278
rect -8576 409254 592500 409276
rect -8576 409018 -7454 409254
rect -7218 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 155786 409254
rect 156022 409018 191786 409254
rect 192022 409018 299786 409254
rect 300022 409018 335786 409254
rect 336022 409018 371786 409254
rect 372022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591142 409254
rect 591378 409018 592500 409254
rect -8576 408934 592500 409018
rect -8576 408698 -7454 408934
rect -7218 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 155786 408934
rect 156022 408698 191786 408934
rect 192022 408698 299786 408934
rect 300022 408698 335786 408934
rect 336022 408698 371786 408934
rect 372022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591142 408934
rect 591378 408698 592500 408934
rect -8576 408676 592500 408698
rect -7636 408674 -7036 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 155604 408674 156204 408676
rect 191604 408674 192204 408676
rect 299604 408674 300204 408676
rect 335604 408674 336204 408676
rect 371604 408674 372204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590960 408674 591560 408676
rect -5756 405676 -5156 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 188004 405676 188604 405678
rect 296004 405676 296604 405678
rect 332004 405676 332604 405678
rect 368004 405676 368604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589080 405676 589680 405678
rect -6696 405654 590620 405676
rect -6696 405418 -5574 405654
rect -5338 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 188186 405654
rect 188422 405418 296186 405654
rect 296422 405418 332186 405654
rect 332422 405418 368186 405654
rect 368422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589262 405654
rect 589498 405418 590620 405654
rect -6696 405334 590620 405418
rect -6696 405098 -5574 405334
rect -5338 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 188186 405334
rect 188422 405098 296186 405334
rect 296422 405098 332186 405334
rect 332422 405098 368186 405334
rect 368422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589262 405334
rect 589498 405098 590620 405334
rect -6696 405076 590620 405098
rect -5756 405074 -5156 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 188004 405074 188604 405076
rect 296004 405074 296604 405076
rect 332004 405074 332604 405076
rect 368004 405074 368604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589080 405074 589680 405076
rect -3876 402076 -3276 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 184404 402076 185004 402078
rect 292404 402076 293004 402078
rect 328404 402076 329004 402078
rect 364404 402076 365004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587200 402076 587800 402078
rect -4816 402054 588740 402076
rect -4816 401818 -3694 402054
rect -3458 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 184586 402054
rect 184822 401818 292586 402054
rect 292822 401818 328586 402054
rect 328822 401818 364586 402054
rect 364822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587382 402054
rect 587618 401818 588740 402054
rect -4816 401734 588740 401818
rect -4816 401498 -3694 401734
rect -3458 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 184586 401734
rect 184822 401498 292586 401734
rect 292822 401498 328586 401734
rect 328822 401498 364586 401734
rect 364822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587382 401734
rect 587618 401498 588740 401734
rect -4816 401476 588740 401498
rect -3876 401474 -3276 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 184404 401474 185004 401476
rect 292404 401474 293004 401476
rect 328404 401474 329004 401476
rect 364404 401474 365004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587200 401474 587800 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 204208 398476 204528 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 204250 398454
rect 204486 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 204250 398134
rect 204486 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 204208 397874 204528 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8576 391276 -7976 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 137604 391276 138204 391278
rect 173604 391276 174204 391278
rect 281604 391276 282204 391278
rect 317604 391276 318204 391278
rect 353604 391276 354204 391278
rect 389604 391276 390204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591900 391276 592500 391278
rect -8576 391254 592500 391276
rect -8576 391018 -8394 391254
rect -8158 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 137786 391254
rect 138022 391018 173786 391254
rect 174022 391018 281786 391254
rect 282022 391018 317786 391254
rect 318022 391018 353786 391254
rect 354022 391018 389786 391254
rect 390022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 592082 391254
rect 592318 391018 592500 391254
rect -8576 390934 592500 391018
rect -8576 390698 -8394 390934
rect -8158 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 137786 390934
rect 138022 390698 173786 390934
rect 174022 390698 281786 390934
rect 282022 390698 317786 390934
rect 318022 390698 353786 390934
rect 354022 390698 389786 390934
rect 390022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 592082 390934
rect 592318 390698 592500 390934
rect -8576 390676 592500 390698
rect -8576 390674 -7976 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 137604 390674 138204 390676
rect 173604 390674 174204 390676
rect 281604 390674 282204 390676
rect 317604 390674 318204 390676
rect 353604 390674 354204 390676
rect 389604 390674 390204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591900 390674 592500 390676
rect -6696 387676 -6096 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 134004 387676 134604 387678
rect 170004 387676 170604 387678
rect 278004 387676 278604 387678
rect 314004 387676 314604 387678
rect 350004 387676 350604 387678
rect 386004 387676 386604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 590020 387676 590620 387678
rect -6696 387654 590620 387676
rect -6696 387418 -6514 387654
rect -6278 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 134186 387654
rect 134422 387418 170186 387654
rect 170422 387418 278186 387654
rect 278422 387418 314186 387654
rect 314422 387418 350186 387654
rect 350422 387418 386186 387654
rect 386422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590202 387654
rect 590438 387418 590620 387654
rect -6696 387334 590620 387418
rect -6696 387098 -6514 387334
rect -6278 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 134186 387334
rect 134422 387098 170186 387334
rect 170422 387098 278186 387334
rect 278422 387098 314186 387334
rect 314422 387098 350186 387334
rect 350422 387098 386186 387334
rect 386422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590202 387334
rect 590438 387098 590620 387334
rect -6696 387076 590620 387098
rect -6696 387074 -6096 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 134004 387074 134604 387076
rect 170004 387074 170604 387076
rect 278004 387074 278604 387076
rect 314004 387074 314604 387076
rect 350004 387074 350604 387076
rect 386004 387074 386604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 590020 387074 590620 387076
rect -4816 384076 -4216 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 130404 384076 131004 384078
rect 166404 384076 167004 384078
rect 274404 384076 275004 384078
rect 310404 384076 311004 384078
rect 346404 384076 347004 384078
rect 382404 384076 383004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588140 384076 588740 384078
rect -4816 384054 588740 384076
rect -4816 383818 -4634 384054
rect -4398 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 130586 384054
rect 130822 383818 166586 384054
rect 166822 383818 274586 384054
rect 274822 383818 310586 384054
rect 310822 383818 346586 384054
rect 346822 383818 382586 384054
rect 382822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588322 384054
rect 588558 383818 588740 384054
rect -4816 383734 588740 383818
rect -4816 383498 -4634 383734
rect -4398 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 130586 383734
rect 130822 383498 166586 383734
rect 166822 383498 274586 383734
rect 274822 383498 310586 383734
rect 310822 383498 346586 383734
rect 346822 383498 382586 383734
rect 382822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588322 383734
rect 588558 383498 588740 383734
rect -4816 383476 588740 383498
rect -4816 383474 -4216 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 130404 383474 131004 383476
rect 166404 383474 167004 383476
rect 274404 383474 275004 383476
rect 310404 383474 311004 383476
rect 346404 383474 347004 383476
rect 382404 383474 383004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588140 383474 588740 383476
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 91568 380476 91888 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 219568 380476 219888 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 394604 380476 394924 380478
rect 450804 380476 451404 380478
rect 479568 380476 479888 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 91610 380454
rect 91846 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 219610 380454
rect 219846 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 394646 380454
rect 394882 380218 450986 380454
rect 451222 380218 479610 380454
rect 479846 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 91610 380134
rect 91846 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 219610 380134
rect 219846 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 394646 380134
rect 394882 379898 450986 380134
rect 451222 379898 479610 380134
rect 479846 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 91568 379874 91888 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 219568 379874 219888 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 394604 379874 394924 379876
rect 450804 379874 451404 379876
rect 479568 379874 479888 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -7636 373276 -7036 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 155604 373276 156204 373278
rect 191604 373276 192204 373278
rect 299604 373276 300204 373278
rect 335604 373276 336204 373278
rect 371604 373276 372204 373278
rect 443604 373276 444204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590960 373276 591560 373278
rect -8576 373254 592500 373276
rect -8576 373018 -7454 373254
rect -7218 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 155786 373254
rect 156022 373018 191786 373254
rect 192022 373018 299786 373254
rect 300022 373018 335786 373254
rect 336022 373018 371786 373254
rect 372022 373018 443786 373254
rect 444022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591142 373254
rect 591378 373018 592500 373254
rect -8576 372934 592500 373018
rect -8576 372698 -7454 372934
rect -7218 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 155786 372934
rect 156022 372698 191786 372934
rect 192022 372698 299786 372934
rect 300022 372698 335786 372934
rect 336022 372698 371786 372934
rect 372022 372698 443786 372934
rect 444022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591142 372934
rect 591378 372698 592500 372934
rect -8576 372676 592500 372698
rect -7636 372674 -7036 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 155604 372674 156204 372676
rect 191604 372674 192204 372676
rect 299604 372674 300204 372676
rect 335604 372674 336204 372676
rect 371604 372674 372204 372676
rect 443604 372674 444204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590960 372674 591560 372676
rect -5756 369676 -5156 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 152004 369676 152604 369678
rect 188004 369676 188604 369678
rect 296004 369676 296604 369678
rect 332004 369676 332604 369678
rect 368004 369676 368604 369678
rect 440004 369676 440604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589080 369676 589680 369678
rect -6696 369654 590620 369676
rect -6696 369418 -5574 369654
rect -5338 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 152186 369654
rect 152422 369418 188186 369654
rect 188422 369418 296186 369654
rect 296422 369418 332186 369654
rect 332422 369418 368186 369654
rect 368422 369418 440186 369654
rect 440422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589262 369654
rect 589498 369418 590620 369654
rect -6696 369334 590620 369418
rect -6696 369098 -5574 369334
rect -5338 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 152186 369334
rect 152422 369098 188186 369334
rect 188422 369098 296186 369334
rect 296422 369098 332186 369334
rect 332422 369098 368186 369334
rect 368422 369098 440186 369334
rect 440422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589262 369334
rect 589498 369098 590620 369334
rect -6696 369076 590620 369098
rect -5756 369074 -5156 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 152004 369074 152604 369076
rect 188004 369074 188604 369076
rect 296004 369074 296604 369076
rect 332004 369074 332604 369076
rect 368004 369074 368604 369076
rect 440004 369074 440604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589080 369074 589680 369076
rect -3876 366076 -3276 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 148404 366076 149004 366078
rect 184404 366076 185004 366078
rect 292404 366076 293004 366078
rect 328404 366076 329004 366078
rect 364404 366076 365004 366078
rect 436404 366076 437004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587200 366076 587800 366078
rect -4816 366054 588740 366076
rect -4816 365818 -3694 366054
rect -3458 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 148586 366054
rect 148822 365818 184586 366054
rect 184822 365818 292586 366054
rect 292822 365818 328586 366054
rect 328822 365818 364586 366054
rect 364822 365818 436586 366054
rect 436822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587382 366054
rect 587618 365818 588740 366054
rect -4816 365734 588740 365818
rect -4816 365498 -3694 365734
rect -3458 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 148586 365734
rect 148822 365498 184586 365734
rect 184822 365498 292586 365734
rect 292822 365498 328586 365734
rect 328822 365498 364586 365734
rect 364822 365498 436586 365734
rect 436822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587382 365734
rect 587618 365498 588740 365734
rect -4816 365476 588740 365498
rect -3876 365474 -3276 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 148404 365474 149004 365476
rect 184404 365474 185004 365476
rect 292404 365474 293004 365476
rect 328404 365474 329004 365476
rect 364404 365474 365004 365476
rect 436404 365474 437004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587200 365474 587800 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 76208 362476 76528 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 204208 362476 204528 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 389774 362476 390094 362478
rect 432804 362476 433404 362478
rect 464208 362476 464528 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 76250 362454
rect 76486 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 204250 362454
rect 204486 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 389816 362454
rect 390052 362218 432986 362454
rect 433222 362218 464250 362454
rect 464486 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 76250 362134
rect 76486 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 204250 362134
rect 204486 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 389816 362134
rect 390052 361898 432986 362134
rect 433222 361898 464250 362134
rect 464486 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 76208 361874 76528 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 204208 361874 204528 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 389774 361874 390094 361876
rect 432804 361874 433404 361876
rect 464208 361874 464528 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8576 355276 -7976 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 137604 355276 138204 355278
rect 173604 355276 174204 355278
rect 281604 355276 282204 355278
rect 317604 355276 318204 355278
rect 353604 355276 354204 355278
rect 425604 355276 426204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591900 355276 592500 355278
rect -8576 355254 592500 355276
rect -8576 355018 -8394 355254
rect -8158 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 137786 355254
rect 138022 355018 173786 355254
rect 174022 355018 281786 355254
rect 282022 355018 317786 355254
rect 318022 355018 353786 355254
rect 354022 355018 425786 355254
rect 426022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 592082 355254
rect 592318 355018 592500 355254
rect -8576 354934 592500 355018
rect -8576 354698 -8394 354934
rect -8158 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 137786 354934
rect 138022 354698 173786 354934
rect 174022 354698 281786 354934
rect 282022 354698 317786 354934
rect 318022 354698 353786 354934
rect 354022 354698 425786 354934
rect 426022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 592082 354934
rect 592318 354698 592500 354934
rect -8576 354676 592500 354698
rect -8576 354674 -7976 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 137604 354674 138204 354676
rect 173604 354674 174204 354676
rect 281604 354674 282204 354676
rect 317604 354674 318204 354676
rect 353604 354674 354204 354676
rect 425604 354674 426204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591900 354674 592500 354676
rect -6696 351676 -6096 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 134004 351676 134604 351678
rect 170004 351676 170604 351678
rect 278004 351676 278604 351678
rect 314004 351676 314604 351678
rect 350004 351676 350604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 590020 351676 590620 351678
rect -6696 351654 590620 351676
rect -6696 351418 -6514 351654
rect -6278 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 134186 351654
rect 134422 351418 170186 351654
rect 170422 351418 278186 351654
rect 278422 351418 314186 351654
rect 314422 351418 350186 351654
rect 350422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590202 351654
rect 590438 351418 590620 351654
rect -6696 351334 590620 351418
rect -6696 351098 -6514 351334
rect -6278 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 134186 351334
rect 134422 351098 170186 351334
rect 170422 351098 278186 351334
rect 278422 351098 314186 351334
rect 314422 351098 350186 351334
rect 350422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590202 351334
rect 590438 351098 590620 351334
rect -6696 351076 590620 351098
rect -6696 351074 -6096 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 134004 351074 134604 351076
rect 170004 351074 170604 351076
rect 278004 351074 278604 351076
rect 314004 351074 314604 351076
rect 350004 351074 350604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 590020 351074 590620 351076
rect -4816 348076 -4216 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 130404 348076 131004 348078
rect 166404 348076 167004 348078
rect 274404 348076 275004 348078
rect 310404 348076 311004 348078
rect 346404 348076 347004 348078
rect 382404 348076 383004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588140 348076 588740 348078
rect -4816 348054 588740 348076
rect -4816 347818 -4634 348054
rect -4398 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 130586 348054
rect 130822 347818 166586 348054
rect 166822 347818 274586 348054
rect 274822 347818 310586 348054
rect 310822 347818 346586 348054
rect 346822 347818 382586 348054
rect 382822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588322 348054
rect 588558 347818 588740 348054
rect -4816 347734 588740 347818
rect -4816 347498 -4634 347734
rect -4398 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 130586 347734
rect 130822 347498 166586 347734
rect 166822 347498 274586 347734
rect 274822 347498 310586 347734
rect 310822 347498 346586 347734
rect 346822 347498 382586 347734
rect 382822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588322 347734
rect 588558 347498 588740 347734
rect -4816 347476 588740 347498
rect -4816 347474 -4216 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 130404 347474 131004 347476
rect 166404 347474 167004 347476
rect 274404 347474 275004 347476
rect 310404 347474 311004 347476
rect 346404 347474 347004 347476
rect 382404 347474 383004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588140 347474 588740 347476
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 91568 344476 91888 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 219568 344476 219888 344478
rect 270804 344476 271404 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 479568 344476 479888 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 91610 344454
rect 91846 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 219610 344454
rect 219846 344218 270986 344454
rect 271222 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 479610 344454
rect 479846 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 91610 344134
rect 91846 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 219610 344134
rect 219846 343898 270986 344134
rect 271222 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 479610 344134
rect 479846 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 91568 343874 91888 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 219568 343874 219888 343876
rect 270804 343874 271404 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 479568 343874 479888 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -7636 337276 -7036 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 155604 337276 156204 337278
rect 191604 337276 192204 337278
rect 227604 337276 228204 337278
rect 263604 337276 264204 337278
rect 299604 337276 300204 337278
rect 335604 337276 336204 337278
rect 371604 337276 372204 337278
rect 407604 337276 408204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590960 337276 591560 337278
rect -8576 337254 592500 337276
rect -8576 337018 -7454 337254
rect -7218 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 155786 337254
rect 156022 337018 191786 337254
rect 192022 337018 227786 337254
rect 228022 337018 263786 337254
rect 264022 337018 299786 337254
rect 300022 337018 335786 337254
rect 336022 337018 371786 337254
rect 372022 337018 407786 337254
rect 408022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591142 337254
rect 591378 337018 592500 337254
rect -8576 336934 592500 337018
rect -8576 336698 -7454 336934
rect -7218 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 155786 336934
rect 156022 336698 191786 336934
rect 192022 336698 227786 336934
rect 228022 336698 263786 336934
rect 264022 336698 299786 336934
rect 300022 336698 335786 336934
rect 336022 336698 371786 336934
rect 372022 336698 407786 336934
rect 408022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591142 336934
rect 591378 336698 592500 336934
rect -8576 336676 592500 336698
rect -7636 336674 -7036 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 155604 336674 156204 336676
rect 191604 336674 192204 336676
rect 227604 336674 228204 336676
rect 263604 336674 264204 336676
rect 299604 336674 300204 336676
rect 335604 336674 336204 336676
rect 371604 336674 372204 336676
rect 407604 336674 408204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590960 336674 591560 336676
rect -5756 333676 -5156 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 188004 333676 188604 333678
rect 224004 333676 224604 333678
rect 260004 333676 260604 333678
rect 296004 333676 296604 333678
rect 332004 333676 332604 333678
rect 368004 333676 368604 333678
rect 404004 333676 404604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589080 333676 589680 333678
rect -6696 333654 590620 333676
rect -6696 333418 -5574 333654
rect -5338 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 188186 333654
rect 188422 333418 224186 333654
rect 224422 333418 260186 333654
rect 260422 333418 296186 333654
rect 296422 333418 332186 333654
rect 332422 333418 368186 333654
rect 368422 333418 404186 333654
rect 404422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589262 333654
rect 589498 333418 590620 333654
rect -6696 333334 590620 333418
rect -6696 333098 -5574 333334
rect -5338 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 188186 333334
rect 188422 333098 224186 333334
rect 224422 333098 260186 333334
rect 260422 333098 296186 333334
rect 296422 333098 332186 333334
rect 332422 333098 368186 333334
rect 368422 333098 404186 333334
rect 404422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589262 333334
rect 589498 333098 590620 333334
rect -6696 333076 590620 333098
rect -5756 333074 -5156 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 188004 333074 188604 333076
rect 224004 333074 224604 333076
rect 260004 333074 260604 333076
rect 296004 333074 296604 333076
rect 332004 333074 332604 333076
rect 368004 333074 368604 333076
rect 404004 333074 404604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589080 333074 589680 333076
rect -3876 330076 -3276 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 184404 330076 185004 330078
rect 220404 330076 221004 330078
rect 256404 330076 257004 330078
rect 292404 330076 293004 330078
rect 328404 330076 329004 330078
rect 364404 330076 365004 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587200 330076 587800 330078
rect -4816 330054 588740 330076
rect -4816 329818 -3694 330054
rect -3458 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 184586 330054
rect 184822 329818 220586 330054
rect 220822 329818 256586 330054
rect 256822 329818 292586 330054
rect 292822 329818 328586 330054
rect 328822 329818 364586 330054
rect 364822 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587382 330054
rect 587618 329818 588740 330054
rect -4816 329734 588740 329818
rect -4816 329498 -3694 329734
rect -3458 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 184586 329734
rect 184822 329498 220586 329734
rect 220822 329498 256586 329734
rect 256822 329498 292586 329734
rect 292822 329498 328586 329734
rect 328822 329498 364586 329734
rect 364822 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587382 329734
rect 587618 329498 588740 329734
rect -4816 329476 588740 329498
rect -3876 329474 -3276 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 184404 329474 185004 329476
rect 220404 329474 221004 329476
rect 256404 329474 257004 329476
rect 292404 329474 293004 329476
rect 328404 329474 329004 329476
rect 364404 329474 365004 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587200 329474 587800 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8576 319276 -7976 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 173604 319276 174204 319278
rect 209604 319276 210204 319278
rect 245604 319276 246204 319278
rect 281604 319276 282204 319278
rect 317604 319276 318204 319278
rect 353604 319276 354204 319278
rect 389604 319276 390204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591900 319276 592500 319278
rect -8576 319254 592500 319276
rect -8576 319018 -8394 319254
rect -8158 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 173786 319254
rect 174022 319018 209786 319254
rect 210022 319018 245786 319254
rect 246022 319018 281786 319254
rect 282022 319018 317786 319254
rect 318022 319018 353786 319254
rect 354022 319018 389786 319254
rect 390022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 592082 319254
rect 592318 319018 592500 319254
rect -8576 318934 592500 319018
rect -8576 318698 -8394 318934
rect -8158 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 173786 318934
rect 174022 318698 209786 318934
rect 210022 318698 245786 318934
rect 246022 318698 281786 318934
rect 282022 318698 317786 318934
rect 318022 318698 353786 318934
rect 354022 318698 389786 318934
rect 390022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 592082 318934
rect 592318 318698 592500 318934
rect -8576 318676 592500 318698
rect -8576 318674 -7976 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 173604 318674 174204 318676
rect 209604 318674 210204 318676
rect 245604 318674 246204 318676
rect 281604 318674 282204 318676
rect 317604 318674 318204 318676
rect 353604 318674 354204 318676
rect 389604 318674 390204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591900 318674 592500 318676
rect -6696 315676 -6096 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 590020 315676 590620 315678
rect -6696 315654 590620 315676
rect -6696 315418 -6514 315654
rect -6278 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590202 315654
rect 590438 315418 590620 315654
rect -6696 315334 590620 315418
rect -6696 315098 -6514 315334
rect -6278 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590202 315334
rect 590438 315098 590620 315334
rect -6696 315076 590620 315098
rect -6696 315074 -6096 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 590020 315074 590620 315076
rect -4816 312076 -4216 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588140 312076 588740 312078
rect -4816 312054 588740 312076
rect -4816 311818 -4634 312054
rect -4398 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588322 312054
rect 588558 311818 588740 312054
rect -4816 311734 588740 311818
rect -4816 311498 -4634 311734
rect -4398 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588322 311734
rect 588558 311498 588740 311734
rect -4816 311476 588740 311498
rect -4816 311474 -4216 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588140 311474 588740 311476
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -7636 301276 -7036 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590960 301276 591560 301278
rect -8576 301254 592500 301276
rect -8576 301018 -7454 301254
rect -7218 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591142 301254
rect 591378 301018 592500 301254
rect -8576 300934 592500 301018
rect -8576 300698 -7454 300934
rect -7218 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591142 300934
rect 591378 300698 592500 300934
rect -8576 300676 592500 300698
rect -7636 300674 -7036 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590960 300674 591560 300676
rect -5756 297676 -5156 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589080 297676 589680 297678
rect -6696 297654 590620 297676
rect -6696 297418 -5574 297654
rect -5338 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589262 297654
rect 589498 297418 590620 297654
rect -6696 297334 590620 297418
rect -6696 297098 -5574 297334
rect -5338 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589262 297334
rect 589498 297098 590620 297334
rect -6696 297076 590620 297098
rect -5756 297074 -5156 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589080 297074 589680 297076
rect -3876 294076 -3276 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587200 294076 587800 294078
rect -4816 294054 588740 294076
rect -4816 293818 -3694 294054
rect -3458 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587382 294054
rect 587618 293818 588740 294054
rect -4816 293734 588740 293818
rect -4816 293498 -3694 293734
rect -3458 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587382 293734
rect 587618 293498 588740 293734
rect -4816 293476 588740 293498
rect -3876 293474 -3276 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587200 293474 587800 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8576 283276 -7976 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591900 283276 592500 283278
rect -8576 283254 592500 283276
rect -8576 283018 -8394 283254
rect -8158 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 592082 283254
rect 592318 283018 592500 283254
rect -8576 282934 592500 283018
rect -8576 282698 -8394 282934
rect -8158 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 592082 282934
rect 592318 282698 592500 282934
rect -8576 282676 592500 282698
rect -8576 282674 -7976 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591900 282674 592500 282676
rect -6696 279676 -6096 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 590020 279676 590620 279678
rect -6696 279654 590620 279676
rect -6696 279418 -6514 279654
rect -6278 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590202 279654
rect 590438 279418 590620 279654
rect -6696 279334 590620 279418
rect -6696 279098 -6514 279334
rect -6278 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590202 279334
rect 590438 279098 590620 279334
rect -6696 279076 590620 279098
rect -6696 279074 -6096 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 590020 279074 590620 279076
rect -4816 276076 -4216 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588140 276076 588740 276078
rect -4816 276054 588740 276076
rect -4816 275818 -4634 276054
rect -4398 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588322 276054
rect 588558 275818 588740 276054
rect -4816 275734 588740 275818
rect -4816 275498 -4634 275734
rect -4398 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588322 275734
rect 588558 275498 588740 275734
rect -4816 275476 588740 275498
rect -4816 275474 -4216 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588140 275474 588740 275476
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -7636 265276 -7036 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590960 265276 591560 265278
rect -8576 265254 592500 265276
rect -8576 265018 -7454 265254
rect -7218 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591142 265254
rect 591378 265018 592500 265254
rect -8576 264934 592500 265018
rect -8576 264698 -7454 264934
rect -7218 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591142 264934
rect 591378 264698 592500 264934
rect -8576 264676 592500 264698
rect -7636 264674 -7036 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590960 264674 591560 264676
rect -5756 261676 -5156 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589080 261676 589680 261678
rect -6696 261654 590620 261676
rect -6696 261418 -5574 261654
rect -5338 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589262 261654
rect 589498 261418 590620 261654
rect -6696 261334 590620 261418
rect -6696 261098 -5574 261334
rect -5338 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589262 261334
rect 589498 261098 590620 261334
rect -6696 261076 590620 261098
rect -5756 261074 -5156 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589080 261074 589680 261076
rect -3876 258076 -3276 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587200 258076 587800 258078
rect -4816 258054 588740 258076
rect -4816 257818 -3694 258054
rect -3458 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587382 258054
rect 587618 257818 588740 258054
rect -4816 257734 588740 257818
rect -4816 257498 -3694 257734
rect -3458 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587382 257734
rect 587618 257498 588740 257734
rect -4816 257476 588740 257498
rect -3876 257474 -3276 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587200 257474 587800 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8576 247276 -7976 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591900 247276 592500 247278
rect -8576 247254 592500 247276
rect -8576 247018 -8394 247254
rect -8158 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 592082 247254
rect 592318 247018 592500 247254
rect -8576 246934 592500 247018
rect -8576 246698 -8394 246934
rect -8158 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 592082 246934
rect 592318 246698 592500 246934
rect -8576 246676 592500 246698
rect -8576 246674 -7976 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591900 246674 592500 246676
rect -6696 243676 -6096 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 590020 243676 590620 243678
rect -6696 243654 590620 243676
rect -6696 243418 -6514 243654
rect -6278 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590202 243654
rect 590438 243418 590620 243654
rect -6696 243334 590620 243418
rect -6696 243098 -6514 243334
rect -6278 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590202 243334
rect 590438 243098 590620 243334
rect -6696 243076 590620 243098
rect -6696 243074 -6096 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 590020 243074 590620 243076
rect -4816 240076 -4216 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588140 240076 588740 240078
rect -4816 240054 588740 240076
rect -4816 239818 -4634 240054
rect -4398 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588322 240054
rect 588558 239818 588740 240054
rect -4816 239734 588740 239818
rect -4816 239498 -4634 239734
rect -4398 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588322 239734
rect 588558 239498 588740 239734
rect -4816 239476 588740 239498
rect -4816 239474 -4216 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588140 239474 588740 239476
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -7636 229276 -7036 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590960 229276 591560 229278
rect -8576 229254 592500 229276
rect -8576 229018 -7454 229254
rect -7218 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591142 229254
rect 591378 229018 592500 229254
rect -8576 228934 592500 229018
rect -8576 228698 -7454 228934
rect -7218 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591142 228934
rect 591378 228698 592500 228934
rect -8576 228676 592500 228698
rect -7636 228674 -7036 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590960 228674 591560 228676
rect -5756 225676 -5156 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589080 225676 589680 225678
rect -6696 225654 590620 225676
rect -6696 225418 -5574 225654
rect -5338 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589262 225654
rect 589498 225418 590620 225654
rect -6696 225334 590620 225418
rect -6696 225098 -5574 225334
rect -5338 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589262 225334
rect 589498 225098 590620 225334
rect -6696 225076 590620 225098
rect -5756 225074 -5156 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589080 225074 589680 225076
rect -3876 222076 -3276 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587200 222076 587800 222078
rect -4816 222054 588740 222076
rect -4816 221818 -3694 222054
rect -3458 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587382 222054
rect 587618 221818 588740 222054
rect -4816 221734 588740 221818
rect -4816 221498 -3694 221734
rect -3458 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587382 221734
rect 587618 221498 588740 221734
rect -4816 221476 588740 221498
rect -3876 221474 -3276 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587200 221474 587800 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8576 211276 -7976 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591900 211276 592500 211278
rect -8576 211254 592500 211276
rect -8576 211018 -8394 211254
rect -8158 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 592082 211254
rect 592318 211018 592500 211254
rect -8576 210934 592500 211018
rect -8576 210698 -8394 210934
rect -8158 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 592082 210934
rect 592318 210698 592500 210934
rect -8576 210676 592500 210698
rect -8576 210674 -7976 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591900 210674 592500 210676
rect -6696 207676 -6096 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 590020 207676 590620 207678
rect -6696 207654 590620 207676
rect -6696 207418 -6514 207654
rect -6278 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590202 207654
rect 590438 207418 590620 207654
rect -6696 207334 590620 207418
rect -6696 207098 -6514 207334
rect -6278 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590202 207334
rect 590438 207098 590620 207334
rect -6696 207076 590620 207098
rect -6696 207074 -6096 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 590020 207074 590620 207076
rect -4816 204076 -4216 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588140 204076 588740 204078
rect -4816 204054 588740 204076
rect -4816 203818 -4634 204054
rect -4398 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588322 204054
rect 588558 203818 588740 204054
rect -4816 203734 588740 203818
rect -4816 203498 -4634 203734
rect -4398 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588322 203734
rect 588558 203498 588740 203734
rect -4816 203476 588740 203498
rect -4816 203474 -4216 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588140 203474 588740 203476
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -7636 193276 -7036 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590960 193276 591560 193278
rect -8576 193254 592500 193276
rect -8576 193018 -7454 193254
rect -7218 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591142 193254
rect 591378 193018 592500 193254
rect -8576 192934 592500 193018
rect -8576 192698 -7454 192934
rect -7218 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591142 192934
rect 591378 192698 592500 192934
rect -8576 192676 592500 192698
rect -7636 192674 -7036 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590960 192674 591560 192676
rect -5756 189676 -5156 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589080 189676 589680 189678
rect -6696 189654 590620 189676
rect -6696 189418 -5574 189654
rect -5338 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589262 189654
rect 589498 189418 590620 189654
rect -6696 189334 590620 189418
rect -6696 189098 -5574 189334
rect -5338 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589262 189334
rect 589498 189098 590620 189334
rect -6696 189076 590620 189098
rect -5756 189074 -5156 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589080 189074 589680 189076
rect -3876 186076 -3276 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587200 186076 587800 186078
rect -4816 186054 588740 186076
rect -4816 185818 -3694 186054
rect -3458 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587382 186054
rect 587618 185818 588740 186054
rect -4816 185734 588740 185818
rect -4816 185498 -3694 185734
rect -3458 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587382 185734
rect 587618 185498 588740 185734
rect -4816 185476 588740 185498
rect -3876 185474 -3276 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587200 185474 587800 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 138208 182476 138528 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 138250 182454
rect 138486 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 138250 182134
rect 138486 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 138208 181874 138528 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8576 175276 -7976 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591900 175276 592500 175278
rect -8576 175254 592500 175276
rect -8576 175018 -8394 175254
rect -8158 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 592082 175254
rect 592318 175018 592500 175254
rect -8576 174934 592500 175018
rect -8576 174698 -8394 174934
rect -8158 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 592082 174934
rect 592318 174698 592500 174934
rect -8576 174676 592500 174698
rect -8576 174674 -7976 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591900 174674 592500 174676
rect -6696 171676 -6096 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 590020 171676 590620 171678
rect -6696 171654 590620 171676
rect -6696 171418 -6514 171654
rect -6278 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590202 171654
rect 590438 171418 590620 171654
rect -6696 171334 590620 171418
rect -6696 171098 -6514 171334
rect -6278 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590202 171334
rect 590438 171098 590620 171334
rect -6696 171076 590620 171098
rect -6696 171074 -6096 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 590020 171074 590620 171076
rect -4816 168076 -4216 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588140 168076 588740 168078
rect -4816 168054 588740 168076
rect -4816 167818 -4634 168054
rect -4398 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588322 168054
rect 588558 167818 588740 168054
rect -4816 167734 588740 167818
rect -4816 167498 -4634 167734
rect -4398 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588322 167734
rect 588558 167498 588740 167734
rect -4816 167476 588740 167498
rect -4816 167474 -4216 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588140 167474 588740 167476
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 153568 164476 153888 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 153610 164454
rect 153846 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 153610 164134
rect 153846 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 153568 163874 153888 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -7636 157276 -7036 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590960 157276 591560 157278
rect -8576 157254 592500 157276
rect -8576 157018 -7454 157254
rect -7218 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591142 157254
rect 591378 157018 592500 157254
rect -8576 156934 592500 157018
rect -8576 156698 -7454 156934
rect -7218 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591142 156934
rect 591378 156698 592500 156934
rect -8576 156676 592500 156698
rect -7636 156674 -7036 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590960 156674 591560 156676
rect -5756 153676 -5156 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589080 153676 589680 153678
rect -6696 153654 590620 153676
rect -6696 153418 -5574 153654
rect -5338 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589262 153654
rect 589498 153418 590620 153654
rect -6696 153334 590620 153418
rect -6696 153098 -5574 153334
rect -5338 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589262 153334
rect 589498 153098 590620 153334
rect -6696 153076 590620 153098
rect -5756 153074 -5156 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589080 153074 589680 153076
rect -3876 150076 -3276 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587200 150076 587800 150078
rect -4816 150054 588740 150076
rect -4816 149818 -3694 150054
rect -3458 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587382 150054
rect 587618 149818 588740 150054
rect -4816 149734 588740 149818
rect -4816 149498 -3694 149734
rect -3458 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587382 149734
rect 587618 149498 588740 149734
rect -4816 149476 588740 149498
rect -3876 149474 -3276 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587200 149474 587800 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 138208 146476 138528 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 138250 146454
rect 138486 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 138250 146134
rect 138486 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 138208 145874 138528 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8576 139276 -7976 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591900 139276 592500 139278
rect -8576 139254 592500 139276
rect -8576 139018 -8394 139254
rect -8158 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 592082 139254
rect 592318 139018 592500 139254
rect -8576 138934 592500 139018
rect -8576 138698 -8394 138934
rect -8158 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 592082 138934
rect 592318 138698 592500 138934
rect -8576 138676 592500 138698
rect -8576 138674 -7976 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591900 138674 592500 138676
rect -6696 135676 -6096 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 590020 135676 590620 135678
rect -6696 135654 590620 135676
rect -6696 135418 -6514 135654
rect -6278 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590202 135654
rect 590438 135418 590620 135654
rect -6696 135334 590620 135418
rect -6696 135098 -6514 135334
rect -6278 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590202 135334
rect 590438 135098 590620 135334
rect -6696 135076 590620 135098
rect -6696 135074 -6096 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 590020 135074 590620 135076
rect -4816 132076 -4216 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588140 132076 588740 132078
rect -4816 132054 588740 132076
rect -4816 131818 -4634 132054
rect -4398 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588322 132054
rect 588558 131818 588740 132054
rect -4816 131734 588740 131818
rect -4816 131498 -4634 131734
rect -4398 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588322 131734
rect 588558 131498 588740 131734
rect -4816 131476 588740 131498
rect -4816 131474 -4216 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588140 131474 588740 131476
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 153568 128476 153888 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 153610 128454
rect 153846 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 153610 128134
rect 153846 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 153568 127874 153888 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -7636 121276 -7036 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590960 121276 591560 121278
rect -8576 121254 592500 121276
rect -8576 121018 -7454 121254
rect -7218 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591142 121254
rect 591378 121018 592500 121254
rect -8576 120934 592500 121018
rect -8576 120698 -7454 120934
rect -7218 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591142 120934
rect 591378 120698 592500 120934
rect -8576 120676 592500 120698
rect -7636 120674 -7036 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590960 120674 591560 120676
rect -5756 117676 -5156 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589080 117676 589680 117678
rect -6696 117654 590620 117676
rect -6696 117418 -5574 117654
rect -5338 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589262 117654
rect 589498 117418 590620 117654
rect -6696 117334 590620 117418
rect -6696 117098 -5574 117334
rect -5338 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589262 117334
rect 589498 117098 590620 117334
rect -6696 117076 590620 117098
rect -5756 117074 -5156 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589080 117074 589680 117076
rect -3876 114076 -3276 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587200 114076 587800 114078
rect -4816 114054 588740 114076
rect -4816 113818 -3694 114054
rect -3458 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587382 114054
rect 587618 113818 588740 114054
rect -4816 113734 588740 113818
rect -4816 113498 -3694 113734
rect -3458 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587382 113734
rect 587618 113498 588740 113734
rect -4816 113476 588740 113498
rect -3876 113474 -3276 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587200 113474 587800 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8576 103276 -7976 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591900 103276 592500 103278
rect -8576 103254 592500 103276
rect -8576 103018 -8394 103254
rect -8158 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 592082 103254
rect 592318 103018 592500 103254
rect -8576 102934 592500 103018
rect -8576 102698 -8394 102934
rect -8158 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 592082 102934
rect 592318 102698 592500 102934
rect -8576 102676 592500 102698
rect -8576 102674 -7976 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591900 102674 592500 102676
rect -6696 99676 -6096 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 590020 99676 590620 99678
rect -6696 99654 590620 99676
rect -6696 99418 -6514 99654
rect -6278 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590202 99654
rect 590438 99418 590620 99654
rect -6696 99334 590620 99418
rect -6696 99098 -6514 99334
rect -6278 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590202 99334
rect 590438 99098 590620 99334
rect -6696 99076 590620 99098
rect -6696 99074 -6096 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 590020 99074 590620 99076
rect -4816 96076 -4216 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588140 96076 588740 96078
rect -4816 96054 588740 96076
rect -4816 95818 -4634 96054
rect -4398 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588322 96054
rect 588558 95818 588740 96054
rect -4816 95734 588740 95818
rect -4816 95498 -4634 95734
rect -4398 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588322 95734
rect 588558 95498 588740 95734
rect -4816 95476 588740 95498
rect -4816 95474 -4216 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588140 95474 588740 95476
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -7636 85276 -7036 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590960 85276 591560 85278
rect -8576 85254 592500 85276
rect -8576 85018 -7454 85254
rect -7218 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591142 85254
rect 591378 85018 592500 85254
rect -8576 84934 592500 85018
rect -8576 84698 -7454 84934
rect -7218 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591142 84934
rect 591378 84698 592500 84934
rect -8576 84676 592500 84698
rect -7636 84674 -7036 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590960 84674 591560 84676
rect -5756 81676 -5156 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589080 81676 589680 81678
rect -6696 81654 590620 81676
rect -6696 81418 -5574 81654
rect -5338 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589262 81654
rect 589498 81418 590620 81654
rect -6696 81334 590620 81418
rect -6696 81098 -5574 81334
rect -5338 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589262 81334
rect 589498 81098 590620 81334
rect -6696 81076 590620 81098
rect -5756 81074 -5156 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589080 81074 589680 81076
rect -3876 78076 -3276 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587200 78076 587800 78078
rect -4816 78054 588740 78076
rect -4816 77818 -3694 78054
rect -3458 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587382 78054
rect 587618 77818 588740 78054
rect -4816 77734 588740 77818
rect -4816 77498 -3694 77734
rect -3458 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587382 77734
rect 587618 77498 588740 77734
rect -4816 77476 588740 77498
rect -3876 77474 -3276 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587200 77474 587800 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8576 67276 -7976 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591900 67276 592500 67278
rect -8576 67254 592500 67276
rect -8576 67018 -8394 67254
rect -8158 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 592082 67254
rect 592318 67018 592500 67254
rect -8576 66934 592500 67018
rect -8576 66698 -8394 66934
rect -8158 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 592082 66934
rect 592318 66698 592500 66934
rect -8576 66676 592500 66698
rect -8576 66674 -7976 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591900 66674 592500 66676
rect -6696 63676 -6096 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 590020 63676 590620 63678
rect -6696 63654 590620 63676
rect -6696 63418 -6514 63654
rect -6278 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590202 63654
rect 590438 63418 590620 63654
rect -6696 63334 590620 63418
rect -6696 63098 -6514 63334
rect -6278 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590202 63334
rect 590438 63098 590620 63334
rect -6696 63076 590620 63098
rect -6696 63074 -6096 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 590020 63074 590620 63076
rect -4816 60076 -4216 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588140 60076 588740 60078
rect -4816 60054 588740 60076
rect -4816 59818 -4634 60054
rect -4398 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588322 60054
rect 588558 59818 588740 60054
rect -4816 59734 588740 59818
rect -4816 59498 -4634 59734
rect -4398 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588322 59734
rect 588558 59498 588740 59734
rect -4816 59476 588740 59498
rect -4816 59474 -4216 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588140 59474 588740 59476
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -7636 49276 -7036 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590960 49276 591560 49278
rect -8576 49254 592500 49276
rect -8576 49018 -7454 49254
rect -7218 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591142 49254
rect 591378 49018 592500 49254
rect -8576 48934 592500 49018
rect -8576 48698 -7454 48934
rect -7218 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591142 48934
rect 591378 48698 592500 48934
rect -8576 48676 592500 48698
rect -7636 48674 -7036 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590960 48674 591560 48676
rect -5756 45676 -5156 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589080 45676 589680 45678
rect -6696 45654 590620 45676
rect -6696 45418 -5574 45654
rect -5338 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589262 45654
rect 589498 45418 590620 45654
rect -6696 45334 590620 45418
rect -6696 45098 -5574 45334
rect -5338 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589262 45334
rect 589498 45098 590620 45334
rect -6696 45076 590620 45098
rect -5756 45074 -5156 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589080 45074 589680 45076
rect -3876 42076 -3276 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587200 42076 587800 42078
rect -4816 42054 588740 42076
rect -4816 41818 -3694 42054
rect -3458 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587382 42054
rect 587618 41818 588740 42054
rect -4816 41734 588740 41818
rect -4816 41498 -3694 41734
rect -3458 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587382 41734
rect 587618 41498 588740 41734
rect -4816 41476 588740 41498
rect -3876 41474 -3276 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587200 41474 587800 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8576 31276 -7976 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591900 31276 592500 31278
rect -8576 31254 592500 31276
rect -8576 31018 -8394 31254
rect -8158 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 592082 31254
rect 592318 31018 592500 31254
rect -8576 30934 592500 31018
rect -8576 30698 -8394 30934
rect -8158 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 592082 30934
rect 592318 30698 592500 30934
rect -8576 30676 592500 30698
rect -8576 30674 -7976 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591900 30674 592500 30676
rect -6696 27676 -6096 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 590020 27676 590620 27678
rect -6696 27654 590620 27676
rect -6696 27418 -6514 27654
rect -6278 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590202 27654
rect 590438 27418 590620 27654
rect -6696 27334 590620 27418
rect -6696 27098 -6514 27334
rect -6278 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590202 27334
rect 590438 27098 590620 27334
rect -6696 27076 590620 27098
rect -6696 27074 -6096 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 590020 27074 590620 27076
rect -4816 24076 -4216 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588140 24076 588740 24078
rect -4816 24054 588740 24076
rect -4816 23818 -4634 24054
rect -4398 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588322 24054
rect 588558 23818 588740 24054
rect -4816 23734 588740 23818
rect -4816 23498 -4634 23734
rect -4398 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588322 23734
rect 588558 23498 588740 23734
rect -4816 23476 588740 23498
rect -4816 23474 -4216 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588140 23474 588740 23476
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -7636 13276 -7036 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590960 13276 591560 13278
rect -8576 13254 592500 13276
rect -8576 13018 -7454 13254
rect -7218 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591142 13254
rect 591378 13018 592500 13254
rect -8576 12934 592500 13018
rect -8576 12698 -7454 12934
rect -7218 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591142 12934
rect 591378 12698 592500 12934
rect -8576 12676 592500 12698
rect -7636 12674 -7036 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590960 12674 591560 12676
rect -5756 9676 -5156 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589080 9676 589680 9678
rect -6696 9654 590620 9676
rect -6696 9418 -5574 9654
rect -5338 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589262 9654
rect 589498 9418 590620 9654
rect -6696 9334 590620 9418
rect -6696 9098 -5574 9334
rect -5338 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589262 9334
rect 589498 9098 590620 9334
rect -6696 9076 590620 9098
rect -5756 9074 -5156 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589080 9074 589680 9076
rect -3876 6076 -3276 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587200 6076 587800 6078
rect -4816 6054 588740 6076
rect -4816 5818 -3694 6054
rect -3458 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587382 6054
rect 587618 5818 588740 6054
rect -4816 5734 588740 5818
rect -4816 5498 -3694 5734
rect -3458 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587382 5734
rect 587618 5498 588740 5734
rect -4816 5476 588740 5498
rect -3876 5474 -3276 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587200 5474 587800 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 4586 -2226
rect 4822 -2462 40586 -2226
rect 40822 -2462 76586 -2226
rect 76822 -2462 112586 -2226
rect 112822 -2462 148586 -2226
rect 148822 -2462 184586 -2226
rect 184822 -2462 220586 -2226
rect 220822 -2462 256586 -2226
rect 256822 -2462 292586 -2226
rect 292822 -2462 328586 -2226
rect 328822 -2462 364586 -2226
rect 364822 -2462 400586 -2226
rect 400822 -2462 436586 -2226
rect 436822 -2462 472586 -2226
rect 472822 -2462 508586 -2226
rect 508822 -2462 544586 -2226
rect 544822 -2462 580586 -2226
rect 580822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 4586 -2546
rect 4822 -2782 40586 -2546
rect 40822 -2782 76586 -2546
rect 76822 -2782 112586 -2546
rect 112822 -2782 148586 -2546
rect 148822 -2782 184586 -2546
rect 184822 -2782 220586 -2546
rect 220822 -2782 256586 -2546
rect 256822 -2782 292586 -2546
rect 292822 -2782 328586 -2546
rect 328822 -2782 364586 -2546
rect 364822 -2782 400586 -2546
rect 400822 -2782 436586 -2546
rect 436822 -2782 472586 -2546
rect 472822 -2782 508586 -2546
rect 508822 -2782 544586 -2546
rect 544822 -2782 580586 -2546
rect 580822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 22586 -3166
rect 22822 -3402 58586 -3166
rect 58822 -3402 94586 -3166
rect 94822 -3402 130586 -3166
rect 130822 -3402 166586 -3166
rect 166822 -3402 202586 -3166
rect 202822 -3402 238586 -3166
rect 238822 -3402 274586 -3166
rect 274822 -3402 310586 -3166
rect 310822 -3402 346586 -3166
rect 346822 -3402 382586 -3166
rect 382822 -3402 418586 -3166
rect 418822 -3402 454586 -3166
rect 454822 -3402 490586 -3166
rect 490822 -3402 526586 -3166
rect 526822 -3402 562586 -3166
rect 562822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 22586 -3486
rect 22822 -3722 58586 -3486
rect 58822 -3722 94586 -3486
rect 94822 -3722 130586 -3486
rect 130822 -3722 166586 -3486
rect 166822 -3722 202586 -3486
rect 202822 -3722 238586 -3486
rect 238822 -3722 274586 -3486
rect 274822 -3722 310586 -3486
rect 310822 -3722 346586 -3486
rect 346822 -3722 382586 -3486
rect 382822 -3722 418586 -3486
rect 418822 -3722 454586 -3486
rect 454822 -3722 490586 -3486
rect 490822 -3722 526586 -3486
rect 526822 -3722 562586 -3486
rect 562822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 8186 -4106
rect 8422 -4342 44186 -4106
rect 44422 -4342 80186 -4106
rect 80422 -4342 116186 -4106
rect 116422 -4342 152186 -4106
rect 152422 -4342 188186 -4106
rect 188422 -4342 224186 -4106
rect 224422 -4342 260186 -4106
rect 260422 -4342 296186 -4106
rect 296422 -4342 332186 -4106
rect 332422 -4342 368186 -4106
rect 368422 -4342 404186 -4106
rect 404422 -4342 440186 -4106
rect 440422 -4342 476186 -4106
rect 476422 -4342 512186 -4106
rect 512422 -4342 548186 -4106
rect 548422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 8186 -4426
rect 8422 -4662 44186 -4426
rect 44422 -4662 80186 -4426
rect 80422 -4662 116186 -4426
rect 116422 -4662 152186 -4426
rect 152422 -4662 188186 -4426
rect 188422 -4662 224186 -4426
rect 224422 -4662 260186 -4426
rect 260422 -4662 296186 -4426
rect 296422 -4662 332186 -4426
rect 332422 -4662 368186 -4426
rect 368422 -4662 404186 -4426
rect 404422 -4662 440186 -4426
rect 440422 -4662 476186 -4426
rect 476422 -4662 512186 -4426
rect 512422 -4662 548186 -4426
rect 548422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 26186 -5046
rect 26422 -5282 62186 -5046
rect 62422 -5282 98186 -5046
rect 98422 -5282 134186 -5046
rect 134422 -5282 170186 -5046
rect 170422 -5282 206186 -5046
rect 206422 -5282 242186 -5046
rect 242422 -5282 278186 -5046
rect 278422 -5282 314186 -5046
rect 314422 -5282 350186 -5046
rect 350422 -5282 386186 -5046
rect 386422 -5282 422186 -5046
rect 422422 -5282 458186 -5046
rect 458422 -5282 494186 -5046
rect 494422 -5282 530186 -5046
rect 530422 -5282 566186 -5046
rect 566422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 26186 -5366
rect 26422 -5602 62186 -5366
rect 62422 -5602 98186 -5366
rect 98422 -5602 134186 -5366
rect 134422 -5602 170186 -5366
rect 170422 -5602 206186 -5366
rect 206422 -5602 242186 -5366
rect 242422 -5602 278186 -5366
rect 278422 -5602 314186 -5366
rect 314422 -5602 350186 -5366
rect 350422 -5602 386186 -5366
rect 386422 -5602 422186 -5366
rect 422422 -5602 458186 -5366
rect 458422 -5602 494186 -5366
rect 494422 -5602 530186 -5366
rect 530422 -5602 566186 -5366
rect 566422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 11786 -5986
rect 12022 -6222 47786 -5986
rect 48022 -6222 83786 -5986
rect 84022 -6222 119786 -5986
rect 120022 -6222 155786 -5986
rect 156022 -6222 191786 -5986
rect 192022 -6222 227786 -5986
rect 228022 -6222 263786 -5986
rect 264022 -6222 299786 -5986
rect 300022 -6222 335786 -5986
rect 336022 -6222 371786 -5986
rect 372022 -6222 407786 -5986
rect 408022 -6222 443786 -5986
rect 444022 -6222 479786 -5986
rect 480022 -6222 515786 -5986
rect 516022 -6222 551786 -5986
rect 552022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 11786 -6306
rect 12022 -6542 47786 -6306
rect 48022 -6542 83786 -6306
rect 84022 -6542 119786 -6306
rect 120022 -6542 155786 -6306
rect 156022 -6542 191786 -6306
rect 192022 -6542 227786 -6306
rect 228022 -6542 263786 -6306
rect 264022 -6542 299786 -6306
rect 300022 -6542 335786 -6306
rect 336022 -6542 371786 -6306
rect 372022 -6542 407786 -6306
rect 408022 -6542 443786 -6306
rect 444022 -6542 479786 -6306
rect 480022 -6542 515786 -6306
rect 516022 -6542 551786 -6306
rect 552022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 29786 -6926
rect 30022 -7162 65786 -6926
rect 66022 -7162 101786 -6926
rect 102022 -7162 137786 -6926
rect 138022 -7162 173786 -6926
rect 174022 -7162 209786 -6926
rect 210022 -7162 245786 -6926
rect 246022 -7162 281786 -6926
rect 282022 -7162 317786 -6926
rect 318022 -7162 353786 -6926
rect 354022 -7162 389786 -6926
rect 390022 -7162 425786 -6926
rect 426022 -7162 461786 -6926
rect 462022 -7162 497786 -6926
rect 498022 -7162 533786 -6926
rect 534022 -7162 569786 -6926
rect 570022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 29786 -7246
rect 30022 -7482 65786 -7246
rect 66022 -7482 101786 -7246
rect 102022 -7482 137786 -7246
rect 138022 -7482 173786 -7246
rect 174022 -7482 209786 -7246
rect 210022 -7482 245786 -7246
rect 246022 -7482 281786 -7246
rect 282022 -7482 317786 -7246
rect 318022 -7482 353786 -7246
rect 354022 -7482 389786 -7246
rect 390022 -7482 425786 -7246
rect 426022 -7482 461786 -7246
rect 462022 -7482 497786 -7246
rect 498022 -7482 533786 -7246
rect 534022 -7482 569786 -7246
rect 570022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
use MM2hdmi  proj_7
timestamp 1608124775
transform 1 0 200000 0 1 520000
box 0 0 20000 40000
use challenge  proj_6
timestamp 1608124775
transform 1 0 480000 0 1 520000
box 0 0 31344 34764
use watch_hhmm  proj_5
timestamp 1608124775
transform 1 0 384000 0 1 350000
box 0 0 31275 33419
use asic_freq  proj_4
timestamp 1608124775
transform 1 0 300000 0 1 500000
box 0 0 77867 80011
use spinet5  proj_3
timestamp 1608124775
transform 1 0 200000 0 1 340000
box 0 0 66678 68822
use vga_clock  proj_2
timestamp 1608124775
transform 1 0 460000 0 1 340000
box 0 0 45405 47549
use ws2812  proj_1
timestamp 1608124775
transform 1 0 72000 0 1 340000
box 0 0 54206 56350
use seven_segment_seconds  proj_0
timestamp 1608124775
transform 1 0 86000 0 1 520000
box 0 0 29760 31904
use multi_project_harness  mprj
timestamp 1608124775
transform 1 0 134000 0 1 120000
box 0 0 300000 80000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
