magic
tech sky130A
magscale 1 2
timestamp 1608040051
<< locali >>
rect 153577 666587 153611 684437
rect 153485 647275 153519 656829
rect 153301 636259 153335 645813
rect 153301 589339 153335 598893
rect 315221 578459 315255 579309
rect 317429 578391 317463 579309
rect 343005 578323 343039 579309
rect 364257 578255 364291 579309
rect 99331 518721 99423 518755
rect 99389 518687 99423 518721
rect 118709 518687 118743 518721
rect 118559 518653 118743 518687
rect 106289 518483 106323 518585
rect 115857 518483 115891 518653
rect 284033 485775 284067 491249
rect 153393 466395 153427 473297
rect 284033 463811 284067 481593
rect 299673 466395 299707 473297
rect 126069 443819 126103 452557
rect 284033 444499 284067 453985
rect 299673 447083 299707 453985
rect 153393 437427 153427 444329
rect 125885 427771 125919 434673
rect 284033 425187 284067 434673
rect 299673 427771 299707 434673
rect 126069 405739 126103 415361
rect 128553 405739 128587 415361
rect 284033 405739 284067 415361
rect 299673 405739 299707 415361
rect 128553 398735 128587 405569
rect 153393 396083 153427 398905
rect 84025 395607 84059 395709
rect 84117 395607 84151 395845
rect 133981 386427 134015 395981
rect 153301 389147 153335 395913
rect 133981 376771 134015 386257
rect 284033 383707 284067 393261
rect 297465 386427 297499 393057
rect 299581 386427 299615 395981
rect 357357 386563 357391 394961
rect 375941 392751 375975 392853
rect 375849 392547 375883 392717
rect 375757 392343 375791 392513
rect 376033 392479 376067 392853
rect 377229 392411 377263 392785
rect 375665 392207 375699 392309
rect 379437 392275 379471 392853
rect 379621 392615 379655 392853
rect 379713 392683 379747 392785
rect 380725 392207 380759 392717
rect 297465 375411 297499 383469
rect 357357 376771 357391 386325
rect 128829 365755 128863 375309
rect 153577 357459 153611 367013
rect 284033 357459 284067 367013
rect 297557 357459 297591 370481
rect 357357 367115 357391 376601
rect 299673 357459 299707 362253
rect 134257 347803 134291 357357
rect 128829 340527 128863 347701
rect 284033 338215 284067 347701
rect 297557 346443 297591 355997
rect 390937 346443 390971 355997
rect 283975 338045 284217 338079
rect 96537 337739 96571 337909
rect 99389 337535 99423 337637
rect 106289 337535 106323 337637
rect 128921 332367 128955 337977
rect 241345 337331 241379 337773
rect 128737 328491 128771 331245
rect 213929 328491 213963 331313
rect 128645 309179 128679 317373
rect 134165 309179 134199 318733
rect 209789 309179 209823 318733
rect 257721 317475 257755 335257
rect 284125 328559 284159 337977
rect 284033 318835 284067 328389
rect 390937 327131 390971 336685
rect 297649 318903 297683 323629
rect 390845 321555 390879 321657
rect 503913 321555 503947 321725
rect 504005 318835 504039 321657
rect 503729 309179 503763 318733
rect 128737 302175 128771 307717
rect 128737 292451 128771 298061
rect 134257 288439 134291 298061
rect 209789 289867 209823 299421
rect 257813 298163 257847 307717
rect 284033 299591 284067 309077
rect 284033 289935 284067 299421
rect 297557 298163 297591 307717
rect 390845 299523 390879 309077
rect 504373 299523 504407 309077
rect 128645 278783 128679 282897
rect 128645 270487 128679 273309
rect 134257 269127 134291 278681
rect 153393 273275 153427 280109
rect 209789 270555 209823 280109
rect 257813 278783 257847 288269
rect 284033 280279 284067 289765
rect 284033 270555 284067 280109
rect 297557 270555 297591 288337
rect 390845 280211 390879 289765
rect 504281 280279 504315 288405
rect 357265 270555 357299 280109
rect 153577 260899 153611 270453
rect 257813 263551 257847 270453
rect 284033 260967 284067 263653
rect 297557 260899 297591 263653
rect 390937 263483 390971 270453
rect 504465 269127 504499 278681
rect 128645 241587 128679 259369
rect 134257 250631 134291 260797
rect 209789 251311 209823 260797
rect 257813 253827 257847 260797
rect 390937 253827 390971 260797
rect 504281 253827 504315 260797
rect 284159 251209 284401 251243
rect 257721 241519 257755 251141
rect 390937 241519 390971 251141
rect 504281 241519 504315 251141
rect 134257 222207 134291 235297
rect 153209 222207 153243 224961
rect 257721 222207 257755 224961
rect 504373 222207 504407 231761
rect 364533 212551 364567 222105
rect 153301 202895 153335 212449
rect 257721 202895 257755 205649
rect 504189 202895 504223 205649
rect 214331 201909 214573 201943
rect 215217 201399 215251 202045
rect 215861 201467 215895 201841
rect 216229 201535 216263 201841
rect 219265 201603 219299 202045
rect 216965 201399 216999 201569
rect 219357 201535 219391 201977
rect 223129 201535 223163 201705
rect 232421 201603 232455 201977
rect 233893 201671 233927 202045
rect 238953 201535 238987 202657
rect 240057 201603 240091 202521
rect 258641 202283 258675 202657
rect 257077 202215 257111 202249
rect 257077 202181 257261 202215
rect 257537 201603 257571 201977
rect 258825 201807 258859 202657
rect 258917 202011 258951 202385
rect 259009 201807 259043 202385
rect 306941 202011 306975 202385
rect 307033 201943 307067 202317
rect 258917 201773 259043 201807
rect 307769 201807 307803 202521
rect 311357 201875 311391 202385
rect 359565 202079 359599 202453
rect 258549 201739 258583 201773
rect 258917 201739 258951 201773
rect 258549 201705 258951 201739
rect 259561 201535 259595 201705
rect 260941 201603 260975 201705
rect 131497 196027 131531 198305
rect 131773 195959 131807 196061
rect 132877 195959 132911 196061
rect 134073 195959 134107 200073
rect 128645 186235 128679 191709
rect 129013 183923 129047 191709
rect 131129 183379 131163 186269
rect 128645 172567 128679 182053
rect 133981 172567 134015 180353
rect 99331 154513 99515 154547
rect 9689 154207 9723 154309
rect 19257 154207 19291 154377
rect 57989 154343 58023 154513
rect 99481 154479 99515 154513
rect 118651 154513 118835 154547
rect 67557 154343 67591 154445
rect 109049 154411 109083 154513
rect 118801 154479 118835 154513
rect 80103 154377 80161 154411
rect 128645 153255 128679 162809
rect 17969 152779 18003 152881
rect 22753 152779 22787 153017
rect 27629 152915 27663 153017
rect 32413 152915 32447 153085
rect 77309 152847 77343 152949
rect 86877 152847 86911 153017
rect 108957 152915 108991 153085
rect 115857 152915 115891 153017
rect 115949 152915 115983 153085
rect 125517 152915 125551 153017
rect 131313 151895 131347 153085
rect 128645 147543 128679 147713
rect 80011 144857 80195 144891
rect 41371 144721 41429 144755
rect 60691 144721 60749 144755
rect 29009 144551 29043 144653
rect 38577 144551 38611 144721
rect 48329 144551 48363 144653
rect 57897 144551 57931 144721
rect 67649 144687 67683 144857
rect 80161 144755 80195 144857
rect 99331 144857 99515 144891
rect 86969 144619 87003 144721
rect 96537 144619 96571 144857
rect 99481 144823 99515 144857
rect 118651 144857 118835 144891
rect 109049 144755 109083 144857
rect 118801 144755 118835 144857
rect 131221 132515 131255 147577
rect 133889 143599 133923 162809
rect 132693 135235 132727 142069
rect 75837 118507 75871 119085
rect 81357 118031 81391 118473
rect 89729 118303 89763 118609
rect 99297 118371 99331 118609
rect 104173 118439 104207 118609
rect 112545 117963 112579 118337
rect 113833 118303 113867 118609
rect 122665 118099 122699 118405
rect 122757 118303 122791 118609
rect 75929 117759 75963 117929
rect 85497 117759 85531 117861
rect 89729 117827 89763 117929
rect 96629 117827 96663 117929
rect 106289 117623 106323 117725
rect 115857 117623 115891 117793
rect 117329 117351 117363 117793
rect 122757 117759 122791 118065
rect 129565 117691 129599 118065
rect 73905 108987 73939 115889
rect 131129 114563 131163 124117
rect 132417 117351 132451 117929
rect 132693 117351 132727 132413
rect 133889 125647 133923 138669
rect 133095 118065 133187 118099
rect 133153 117691 133187 118065
rect 133245 117759 133279 118133
rect 133337 117691 133371 117725
rect 133153 117657 133371 117691
rect 133061 115923 133095 117317
rect 138857 117147 138891 120921
rect 248245 118643 248279 118677
rect 141985 117487 142019 117929
rect 157257 117487 157291 117929
rect 210433 117555 210467 118133
rect 225797 117827 225831 118201
rect 231501 117351 231535 118405
rect 238401 117963 238435 118541
rect 239321 118541 239539 118575
rect 239321 118235 239355 118541
rect 239505 118507 239539 118541
rect 239413 118235 239447 118473
rect 240885 118439 240919 118473
rect 240885 118405 241069 118439
rect 238493 117963 238527 118133
rect 161305 117181 161397 117215
rect 161305 117147 161339 117181
rect 143549 117011 143583 117113
rect 186145 117147 186179 117249
rect 235089 117215 235123 117589
rect 235181 117419 235215 117589
rect 238769 117487 238803 117521
rect 238769 117453 238953 117487
rect 239505 117351 239539 118065
rect 239597 117351 239631 117521
rect 240517 117351 240551 117725
rect 242449 117555 242483 118541
rect 244933 118303 244967 118609
rect 248187 118609 248279 118643
rect 244749 117963 244783 118201
rect 244565 117419 244599 117861
rect 245853 117555 245887 118609
rect 248889 118541 249165 118575
rect 248889 118235 248923 118541
rect 248981 117895 249015 118473
rect 248981 117861 249165 117895
rect 249257 117555 249291 118133
rect 246037 117283 246071 117453
rect 249901 117351 249935 118269
rect 250177 118099 250211 118133
rect 250177 118065 250453 118099
rect 252845 118031 252879 118541
rect 334575 118473 334909 118507
rect 396825 118439 396859 118609
rect 315497 117623 315531 117861
rect 315589 117487 315623 117861
rect 320741 117623 320775 118133
rect 324881 117487 324915 118065
rect 151829 117011 151863 117113
rect 131313 99331 131347 106233
rect 133153 95251 133187 104805
rect 180993 104771 181027 113101
rect 194701 104907 194735 109701
rect 212641 100759 212675 110381
rect 243737 104907 243771 114461
rect 248337 106335 248371 115889
rect 325709 114563 325743 117725
rect 336749 117691 336783 117861
rect 350457 117827 350491 117861
rect 354413 117827 354447 118065
rect 350457 117793 350549 117827
rect 355333 117827 355367 118133
rect 384313 118031 384347 118269
rect 389925 118235 389959 118405
rect 398757 118303 398791 118609
rect 433349 118575 433383 118677
rect 433349 118541 433567 118575
rect 389867 118201 389959 118235
rect 340831 117725 340889 117759
rect 413385 117555 413419 117725
rect 420745 117555 420779 117793
rect 422769 117419 422803 117793
rect 426449 117419 426483 117793
rect 426541 117555 426575 117793
rect 427829 117555 427863 117725
rect 432613 117555 432647 117861
rect 432705 117487 432739 117861
rect 433533 117759 433567 118541
rect 444389 117487 444423 118541
rect 456717 117487 456751 118541
rect 463801 117487 463835 118065
rect 463743 117453 463835 117487
rect 476037 117487 476071 118065
rect 492597 117487 492631 117657
rect 425069 117147 425103 117249
rect 434637 117147 434671 117453
rect 492689 116943 492723 117589
rect 495391 117521 495449 117555
rect 73721 87023 73755 89845
rect 144929 85595 144963 90389
rect 156061 84235 156095 93789
rect 179521 84235 179555 88961
rect 157441 66283 157475 75837
rect 162869 74579 162903 84133
rect 181177 82875 181211 92429
rect 216689 91103 216723 99365
rect 221105 95251 221139 100045
rect 184857 77163 184891 77333
rect 190745 77299 190779 86921
rect 194885 75939 194919 85493
rect 200313 75939 200347 85493
rect 207121 81447 207155 91001
rect 227729 89675 227763 96577
rect 233433 95251 233467 104805
rect 238861 89675 238895 96577
rect 243737 95251 243771 99365
rect 248245 95251 248279 104805
rect 272257 103547 272291 114461
rect 403909 106335 403943 115889
rect 420469 108987 420503 115821
rect 301973 99331 302007 106233
rect 322673 99331 322707 106233
rect 325709 95251 325743 104805
rect 394433 99331 394467 106233
rect 128921 57851 128955 66181
rect 174001 64923 174035 74477
rect 133153 48331 133187 57885
rect 145113 56559 145147 64821
rect 147965 55267 147999 64821
rect 150725 48331 150759 57885
rect 159097 55267 159131 64821
rect 181085 63563 181119 73117
rect 183753 66351 183787 75837
rect 205925 74103 205959 80121
rect 207213 76619 207247 80121
rect 221013 79951 221047 80121
rect 227913 77299 227947 82093
rect 233433 77299 233467 86853
rect 238953 77299 238987 81413
rect 243737 77299 243771 86921
rect 245761 77299 245795 86921
rect 248337 75939 248371 85493
rect 274833 77299 274867 86921
rect 279709 84303 279743 93789
rect 383117 87023 383151 96577
rect 388637 87023 388671 96577
rect 403909 87023 403943 96577
rect 415041 95251 415075 104805
rect 420653 95251 420687 104805
rect 431693 99331 431727 106233
rect 209881 67643 209915 70465
rect 211261 66283 211295 75837
rect 181177 50643 181211 61013
rect 183753 56627 183787 66181
rect 184949 57919 184983 60809
rect 195161 56627 195195 66181
rect 205833 57987 205867 60809
rect 184949 48331 184983 51085
rect 200313 48331 200347 57885
rect 207121 56627 207155 66181
rect 212733 57919 212767 68357
rect 233433 62815 233467 67541
rect 234721 66283 234755 67677
rect 240241 67643 240275 70465
rect 244289 66283 244323 75837
rect 245761 66283 245795 75837
rect 271889 70295 271923 75837
rect 279709 74579 279743 84133
rect 322673 77299 322707 86921
rect 301973 67643 302007 77129
rect 325709 75939 325743 85493
rect 358001 79951 358035 80121
rect 394433 77299 394467 86921
rect 426173 85595 426207 95149
rect 341349 67643 341383 77129
rect 383209 67643 383243 77129
rect 388729 67643 388763 77129
rect 404001 67643 404035 77129
rect 426081 69683 426115 84133
rect 431601 66283 431635 75837
rect 73813 35343 73847 48229
rect 209881 46971 209915 51153
rect 212549 51119 212583 57885
rect 216873 48331 216907 57885
rect 240149 56627 240183 58021
rect 248337 56627 248371 66181
rect 227913 48331 227947 53125
rect 234721 46971 234755 56525
rect 279893 48331 279927 57885
rect 301789 48331 301823 57885
rect 322673 48331 322707 57885
rect 325525 56627 325559 66181
rect 248337 46971 248371 48297
rect 150817 38607 150851 41429
rect 128921 29019 128955 38573
rect 133153 31059 133187 38573
rect 157349 37315 157383 46869
rect 150725 27659 150759 37213
rect 181177 31671 181211 44081
rect 190745 29019 190779 46869
rect 194701 37315 194735 46869
rect 211261 45611 211295 46937
rect 200405 29019 200439 38573
rect 207213 35955 207247 45509
rect 238861 41327 238895 45849
rect 276121 37315 276155 46869
rect 229201 29019 229235 31841
rect 74273 12359 74307 20009
rect 143641 9707 143675 19261
rect 157349 9707 157383 27557
rect 175565 24871 175599 26265
rect 178049 24735 178083 25041
rect 168389 9707 168423 12461
rect 168331 9605 168481 9639
rect 168205 9435 168239 9537
rect 125793 7055 125827 7157
rect 174001 6919 174035 20009
rect 178141 9639 178175 12325
rect 179429 6919 179463 24769
rect 184949 19363 184983 28917
rect 234721 27659 234755 37213
rect 238861 27659 238895 37213
rect 244289 31671 244323 37213
rect 245761 31739 245795 37213
rect 248337 27659 248371 37213
rect 271889 27659 271923 37213
rect 322673 29019 322707 38573
rect 325709 29087 325743 46869
rect 341533 45611 341567 51153
rect 383209 48331 383243 57885
rect 388729 48331 388763 57885
rect 404001 48331 404035 57885
rect 415041 56627 415075 66181
rect 341441 38267 341475 45441
rect 358001 38675 358035 48229
rect 243737 26299 243771 27625
rect 190653 18003 190687 19397
rect 205741 19363 205775 22185
rect 233341 19295 233375 22117
rect 200405 12291 200439 19261
rect 234629 18003 234663 22797
rect 244565 11883 244599 19261
rect 274833 9707 274867 18105
rect 276121 18003 276155 27557
rect 279985 19363 280019 28917
rect 183569 6851 183603 9469
rect 183661 6103 183695 9605
rect 301881 8347 301915 26197
rect 325709 9707 325743 27557
rect 357725 26367 357759 29053
rect 383209 29019 383243 38573
rect 404001 29019 404035 38573
rect 414949 35955 414983 45509
rect 425989 37315 426023 46869
rect 431601 37315 431635 46869
rect 431601 31671 431635 37145
rect 357909 22015 357943 26197
rect 383393 19363 383427 25245
rect 383301 9707 383335 12529
rect 394341 9707 394375 19261
rect 415041 16643 415075 26197
rect 420469 18003 420503 27557
rect 431509 16643 431543 26197
rect 414799 8245 415041 8279
rect 412649 7055 412683 7565
rect 169677 4199 169711 4369
rect 205649 4267 205683 4369
rect 57989 3043 58023 3145
rect 62773 3043 62807 3281
rect 67189 595 67223 4165
rect 507041 4063 507075 4097
rect 513941 4097 514159 4131
rect 220093 3791 220127 3961
rect 147689 3315 147723 3417
rect 103529 3043 103563 3281
rect 110613 3043 110647 3281
rect 122849 2839 122883 3281
rect 137937 2839 137971 3281
rect 154589 3247 154623 3485
rect 164157 3247 164191 3485
rect 196725 3383 196759 3621
rect 195621 2907 195655 3145
rect 196633 2839 196667 3213
rect 207673 3043 207707 3349
rect 202797 1343 202831 3009
rect 204453 2839 204487 3009
rect 208869 2907 208903 3417
rect 210341 2975 210375 3417
rect 210433 2975 210467 3553
rect 211169 3451 211203 3621
rect 217977 2907 218011 3757
rect 219725 3519 219759 3757
rect 225061 3723 225095 4029
rect 507041 4029 507317 4063
rect 326445 595 326479 3757
rect 340153 3587 340187 3757
rect 361037 3587 361071 4029
rect 398849 3655 398883 3825
rect 407405 3519 407439 3757
rect 417985 3519 418019 3621
rect 418203 3485 418295 3519
rect 418261 2975 418295 3485
rect 422309 2771 422343 2941
rect 432521 2771 432555 3417
rect 437397 2975 437431 3417
rect 442273 2907 442307 3485
rect 513941 3383 513975 4097
rect 514125 4063 514159 4097
rect 482293 3281 482385 3315
rect 477911 3077 478061 3111
rect 482293 2975 482327 3281
rect 485145 2975 485179 3145
rect 484961 2771 484995 2873
rect 485053 2839 485087 2941
rect 485697 2907 485731 3281
rect 489561 3043 489595 3281
rect 496001 3247 496035 3349
rect 496001 3213 496645 3247
rect 504373 3179 504407 3349
rect 489653 3145 489837 3179
rect 514033 3383 514067 4029
rect 489101 2975 489135 3009
rect 489653 2975 489687 3145
rect 489101 2941 489687 2975
rect 504465 2975 504499 3349
<< viali >>
rect 153577 684437 153611 684471
rect 153577 666553 153611 666587
rect 153485 656829 153519 656863
rect 153485 647241 153519 647275
rect 153301 645813 153335 645847
rect 153301 636225 153335 636259
rect 153301 598893 153335 598927
rect 153301 589305 153335 589339
rect 315221 579309 315255 579343
rect 315221 578425 315255 578459
rect 317429 579309 317463 579343
rect 317429 578357 317463 578391
rect 343005 579309 343039 579343
rect 343005 578289 343039 578323
rect 364257 579309 364291 579343
rect 364257 578221 364291 578255
rect 99297 518721 99331 518755
rect 118709 518721 118743 518755
rect 99389 518653 99423 518687
rect 115857 518653 115891 518687
rect 118525 518653 118559 518687
rect 106289 518585 106323 518619
rect 106289 518449 106323 518483
rect 115857 518449 115891 518483
rect 284033 491249 284067 491283
rect 284033 485741 284067 485775
rect 284033 481593 284067 481627
rect 153393 473297 153427 473331
rect 153393 466361 153427 466395
rect 299673 473297 299707 473331
rect 299673 466361 299707 466395
rect 284033 463777 284067 463811
rect 284033 453985 284067 454019
rect 126069 452557 126103 452591
rect 299673 453985 299707 454019
rect 299673 447049 299707 447083
rect 284033 444465 284067 444499
rect 126069 443785 126103 443819
rect 153393 444329 153427 444363
rect 153393 437393 153427 437427
rect 125885 434673 125919 434707
rect 125885 427737 125919 427771
rect 284033 434673 284067 434707
rect 299673 434673 299707 434707
rect 299673 427737 299707 427771
rect 284033 425153 284067 425187
rect 126069 415361 126103 415395
rect 126069 405705 126103 405739
rect 128553 415361 128587 415395
rect 128553 405705 128587 405739
rect 284033 415361 284067 415395
rect 284033 405705 284067 405739
rect 299673 415361 299707 415395
rect 299673 405705 299707 405739
rect 128553 405569 128587 405603
rect 128553 398701 128587 398735
rect 153393 398905 153427 398939
rect 153393 396049 153427 396083
rect 133981 395981 134015 396015
rect 84117 395845 84151 395879
rect 84025 395709 84059 395743
rect 84025 395573 84059 395607
rect 84117 395573 84151 395607
rect 299581 395981 299615 396015
rect 153301 395913 153335 395947
rect 153301 389113 153335 389147
rect 284033 393261 284067 393295
rect 133981 386393 134015 386427
rect 133981 386257 134015 386291
rect 297465 393057 297499 393091
rect 297465 386393 297499 386427
rect 357357 394961 357391 394995
rect 375941 392853 375975 392887
rect 375849 392717 375883 392751
rect 375941 392717 375975 392751
rect 376033 392853 376067 392887
rect 375757 392513 375791 392547
rect 375849 392513 375883 392547
rect 379437 392853 379471 392887
rect 376033 392445 376067 392479
rect 377229 392785 377263 392819
rect 377229 392377 377263 392411
rect 375665 392309 375699 392343
rect 375757 392309 375791 392343
rect 379621 392853 379655 392887
rect 379713 392785 379747 392819
rect 379713 392649 379747 392683
rect 380725 392717 380759 392751
rect 379621 392581 379655 392615
rect 379437 392241 379471 392275
rect 375665 392173 375699 392207
rect 380725 392173 380759 392207
rect 357357 386529 357391 386563
rect 299581 386393 299615 386427
rect 284033 383673 284067 383707
rect 357357 386325 357391 386359
rect 133981 376737 134015 376771
rect 297465 383469 297499 383503
rect 357357 376737 357391 376771
rect 297465 375377 297499 375411
rect 357357 376601 357391 376635
rect 128829 375309 128863 375343
rect 297557 370481 297591 370515
rect 128829 365721 128863 365755
rect 153577 367013 153611 367047
rect 153577 357425 153611 357459
rect 284033 367013 284067 367047
rect 284033 357425 284067 357459
rect 357357 367081 357391 367115
rect 297557 357425 297591 357459
rect 299673 362253 299707 362287
rect 299673 357425 299707 357459
rect 134257 357357 134291 357391
rect 134257 347769 134291 347803
rect 297557 355997 297591 356031
rect 128829 347701 128863 347735
rect 128829 340493 128863 340527
rect 284033 347701 284067 347735
rect 297557 346409 297591 346443
rect 390937 355997 390971 356031
rect 390937 346409 390971 346443
rect 284033 338181 284067 338215
rect 283941 338045 283975 338079
rect 284217 338045 284251 338079
rect 128921 337977 128955 338011
rect 96537 337909 96571 337943
rect 96537 337705 96571 337739
rect 99389 337637 99423 337671
rect 99389 337501 99423 337535
rect 106289 337637 106323 337671
rect 106289 337501 106323 337535
rect 284125 337977 284159 338011
rect 241345 337773 241379 337807
rect 241345 337297 241379 337331
rect 128921 332333 128955 332367
rect 257721 335257 257755 335291
rect 213929 331313 213963 331347
rect 128737 331245 128771 331279
rect 128737 328457 128771 328491
rect 213929 328457 213963 328491
rect 134165 318733 134199 318767
rect 128645 317373 128679 317407
rect 128645 309145 128679 309179
rect 134165 309145 134199 309179
rect 209789 318733 209823 318767
rect 284125 328525 284159 328559
rect 390937 336685 390971 336719
rect 284033 328389 284067 328423
rect 390937 327097 390971 327131
rect 297649 323629 297683 323663
rect 503913 321725 503947 321759
rect 390845 321657 390879 321691
rect 390845 321521 390879 321555
rect 503913 321521 503947 321555
rect 504005 321657 504039 321691
rect 297649 318869 297683 318903
rect 284033 318801 284067 318835
rect 504005 318801 504039 318835
rect 257721 317441 257755 317475
rect 503729 318733 503763 318767
rect 209789 309145 209823 309179
rect 503729 309145 503763 309179
rect 284033 309077 284067 309111
rect 128737 307717 128771 307751
rect 128737 302141 128771 302175
rect 257813 307717 257847 307751
rect 209789 299421 209823 299455
rect 128737 298061 128771 298095
rect 128737 292417 128771 292451
rect 134257 298061 134291 298095
rect 390845 309077 390879 309111
rect 284033 299557 284067 299591
rect 297557 307717 297591 307751
rect 257813 298129 257847 298163
rect 284033 299421 284067 299455
rect 390845 299489 390879 299523
rect 504373 309077 504407 309111
rect 504373 299489 504407 299523
rect 297557 298129 297591 298163
rect 284033 289901 284067 289935
rect 209789 289833 209823 289867
rect 134257 288405 134291 288439
rect 284033 289765 284067 289799
rect 257813 288269 257847 288303
rect 128645 282897 128679 282931
rect 128645 278749 128679 278783
rect 153393 280109 153427 280143
rect 134257 278681 134291 278715
rect 128645 273309 128679 273343
rect 128645 270453 128679 270487
rect 153393 273241 153427 273275
rect 209789 280109 209823 280143
rect 390845 289765 390879 289799
rect 284033 280245 284067 280279
rect 297557 288337 297591 288371
rect 257813 278749 257847 278783
rect 284033 280109 284067 280143
rect 209789 270521 209823 270555
rect 284033 270521 284067 270555
rect 504281 288405 504315 288439
rect 504281 280245 504315 280279
rect 390845 280177 390879 280211
rect 297557 270521 297591 270555
rect 357265 280109 357299 280143
rect 357265 270521 357299 270555
rect 504465 278681 504499 278715
rect 134257 269093 134291 269127
rect 153577 270453 153611 270487
rect 257813 270453 257847 270487
rect 390937 270453 390971 270487
rect 257813 263517 257847 263551
rect 284033 263653 284067 263687
rect 284033 260933 284067 260967
rect 297557 263653 297591 263687
rect 153577 260865 153611 260899
rect 504465 269093 504499 269127
rect 390937 263449 390971 263483
rect 297557 260865 297591 260899
rect 134257 260797 134291 260831
rect 128645 259369 128679 259403
rect 209789 260797 209823 260831
rect 257813 260797 257847 260831
rect 257813 253793 257847 253827
rect 390937 260797 390971 260831
rect 390937 253793 390971 253827
rect 504281 260797 504315 260831
rect 504281 253793 504315 253827
rect 209789 251277 209823 251311
rect 284125 251209 284159 251243
rect 284401 251209 284435 251243
rect 134257 250597 134291 250631
rect 257721 251141 257755 251175
rect 128645 241553 128679 241587
rect 257721 241485 257755 241519
rect 390937 251141 390971 251175
rect 390937 241485 390971 241519
rect 504281 251141 504315 251175
rect 504281 241485 504315 241519
rect 134257 235297 134291 235331
rect 504373 231761 504407 231795
rect 134257 222173 134291 222207
rect 153209 224961 153243 224995
rect 153209 222173 153243 222207
rect 257721 224961 257755 224995
rect 257721 222173 257755 222207
rect 504373 222173 504407 222207
rect 364533 222105 364567 222139
rect 364533 212517 364567 212551
rect 153301 212449 153335 212483
rect 153301 202861 153335 202895
rect 257721 205649 257755 205683
rect 257721 202861 257755 202895
rect 504189 205649 504223 205683
rect 504189 202861 504223 202895
rect 238953 202657 238987 202691
rect 215217 202045 215251 202079
rect 214297 201909 214331 201943
rect 214573 201909 214607 201943
rect 219265 202045 219299 202079
rect 215861 201841 215895 201875
rect 216229 201841 216263 201875
rect 233893 202045 233927 202079
rect 216229 201501 216263 201535
rect 216965 201569 216999 201603
rect 219265 201569 219299 201603
rect 219357 201977 219391 202011
rect 215861 201433 215895 201467
rect 215217 201365 215251 201399
rect 232421 201977 232455 202011
rect 219357 201501 219391 201535
rect 223129 201705 223163 201739
rect 233893 201637 233927 201671
rect 232421 201569 232455 201603
rect 223129 201501 223163 201535
rect 258641 202657 258675 202691
rect 240057 202521 240091 202555
rect 257077 202249 257111 202283
rect 258641 202249 258675 202283
rect 258825 202657 258859 202691
rect 257261 202181 257295 202215
rect 240057 201569 240091 201603
rect 257537 201977 257571 202011
rect 307769 202521 307803 202555
rect 258917 202385 258951 202419
rect 258917 201977 258951 202011
rect 259009 202385 259043 202419
rect 306941 202385 306975 202419
rect 306941 201977 306975 202011
rect 307033 202317 307067 202351
rect 307033 201909 307067 201943
rect 258549 201773 258583 201807
rect 258825 201773 258859 201807
rect 359565 202453 359599 202487
rect 311357 202385 311391 202419
rect 359565 202045 359599 202079
rect 311357 201841 311391 201875
rect 307769 201773 307803 201807
rect 259561 201705 259595 201739
rect 257537 201569 257571 201603
rect 238953 201501 238987 201535
rect 260941 201705 260975 201739
rect 260941 201569 260975 201603
rect 259561 201501 259595 201535
rect 216965 201365 216999 201399
rect 134073 200073 134107 200107
rect 131497 198305 131531 198339
rect 131497 195993 131531 196027
rect 131773 196061 131807 196095
rect 131773 195925 131807 195959
rect 132877 196061 132911 196095
rect 132877 195925 132911 195959
rect 134073 195925 134107 195959
rect 128645 191709 128679 191743
rect 128645 186201 128679 186235
rect 129013 191709 129047 191743
rect 129013 183889 129047 183923
rect 131129 186269 131163 186303
rect 131129 183345 131163 183379
rect 128645 182053 128679 182087
rect 128645 172533 128679 172567
rect 133981 180353 134015 180387
rect 133981 172533 134015 172567
rect 128645 162809 128679 162843
rect 57989 154513 58023 154547
rect 99297 154513 99331 154547
rect 19257 154377 19291 154411
rect 9689 154309 9723 154343
rect 9689 154173 9723 154207
rect 57989 154309 58023 154343
rect 67557 154445 67591 154479
rect 99481 154445 99515 154479
rect 109049 154513 109083 154547
rect 118617 154513 118651 154547
rect 118801 154445 118835 154479
rect 80069 154377 80103 154411
rect 80161 154377 80195 154411
rect 109049 154377 109083 154411
rect 67557 154309 67591 154343
rect 19257 154173 19291 154207
rect 128645 153221 128679 153255
rect 133889 162809 133923 162843
rect 32413 153085 32447 153119
rect 22753 153017 22787 153051
rect 17969 152881 18003 152915
rect 17969 152745 18003 152779
rect 27629 153017 27663 153051
rect 27629 152881 27663 152915
rect 108957 153085 108991 153119
rect 86877 153017 86911 153051
rect 32413 152881 32447 152915
rect 77309 152949 77343 152983
rect 77309 152813 77343 152847
rect 115949 153085 115983 153119
rect 108957 152881 108991 152915
rect 115857 153017 115891 153051
rect 115857 152881 115891 152915
rect 131313 153085 131347 153119
rect 115949 152881 115983 152915
rect 125517 153017 125551 153051
rect 125517 152881 125551 152915
rect 86877 152813 86911 152847
rect 22753 152745 22787 152779
rect 131313 151861 131347 151895
rect 128645 147713 128679 147747
rect 128645 147509 128679 147543
rect 131221 147577 131255 147611
rect 67649 144857 67683 144891
rect 79977 144857 80011 144891
rect 38577 144721 38611 144755
rect 41337 144721 41371 144755
rect 41429 144721 41463 144755
rect 57897 144721 57931 144755
rect 60657 144721 60691 144755
rect 60749 144721 60783 144755
rect 29009 144653 29043 144687
rect 29009 144517 29043 144551
rect 38577 144517 38611 144551
rect 48329 144653 48363 144687
rect 48329 144517 48363 144551
rect 96537 144857 96571 144891
rect 99297 144857 99331 144891
rect 80161 144721 80195 144755
rect 86969 144721 87003 144755
rect 67649 144653 67683 144687
rect 86969 144585 87003 144619
rect 99481 144789 99515 144823
rect 109049 144857 109083 144891
rect 118617 144857 118651 144891
rect 109049 144721 109083 144755
rect 118801 144721 118835 144755
rect 96537 144585 96571 144619
rect 57897 144517 57931 144551
rect 133889 143565 133923 143599
rect 132693 142069 132727 142103
rect 132693 135201 132727 135235
rect 133889 138669 133923 138703
rect 131221 132481 131255 132515
rect 132693 132413 132727 132447
rect 131129 124117 131163 124151
rect 75837 119085 75871 119119
rect 89729 118609 89763 118643
rect 75837 118473 75871 118507
rect 81357 118473 81391 118507
rect 99297 118609 99331 118643
rect 104173 118609 104207 118643
rect 104173 118405 104207 118439
rect 113833 118609 113867 118643
rect 99297 118337 99331 118371
rect 112545 118337 112579 118371
rect 89729 118269 89763 118303
rect 81357 117997 81391 118031
rect 122757 118609 122791 118643
rect 113833 118269 113867 118303
rect 122665 118405 122699 118439
rect 122757 118269 122791 118303
rect 122665 118065 122699 118099
rect 122757 118065 122791 118099
rect 75929 117929 75963 117963
rect 89729 117929 89763 117963
rect 75929 117725 75963 117759
rect 85497 117861 85531 117895
rect 89729 117793 89763 117827
rect 96629 117929 96663 117963
rect 112545 117929 112579 117963
rect 96629 117793 96663 117827
rect 115857 117793 115891 117827
rect 85497 117725 85531 117759
rect 106289 117725 106323 117759
rect 106289 117589 106323 117623
rect 115857 117589 115891 117623
rect 117329 117793 117363 117827
rect 122757 117725 122791 117759
rect 129565 118065 129599 118099
rect 129565 117657 129599 117691
rect 117329 117317 117363 117351
rect 73905 115889 73939 115923
rect 132417 117929 132451 117963
rect 132417 117317 132451 117351
rect 133889 125613 133923 125647
rect 138857 120921 138891 120955
rect 133245 118133 133279 118167
rect 133061 118065 133095 118099
rect 133245 117725 133279 117759
rect 133337 117725 133371 117759
rect 132693 117317 132727 117351
rect 133061 117317 133095 117351
rect 248245 118677 248279 118711
rect 433349 118677 433383 118711
rect 244933 118609 244967 118643
rect 238401 118541 238435 118575
rect 231501 118405 231535 118439
rect 225797 118201 225831 118235
rect 210433 118133 210467 118167
rect 141985 117929 142019 117963
rect 141985 117453 142019 117487
rect 157257 117929 157291 117963
rect 225797 117793 225831 117827
rect 210433 117521 210467 117555
rect 157257 117453 157291 117487
rect 242449 118541 242483 118575
rect 239321 118201 239355 118235
rect 239413 118473 239447 118507
rect 239505 118473 239539 118507
rect 240885 118473 240919 118507
rect 241069 118405 241103 118439
rect 239413 118201 239447 118235
rect 238401 117929 238435 117963
rect 238493 118133 238527 118167
rect 238493 117929 238527 117963
rect 239505 118065 239539 118099
rect 231501 117317 231535 117351
rect 235089 117589 235123 117623
rect 186145 117249 186179 117283
rect 161397 117181 161431 117215
rect 138857 117113 138891 117147
rect 143549 117113 143583 117147
rect 143549 116977 143583 117011
rect 151829 117113 151863 117147
rect 161305 117113 161339 117147
rect 235181 117589 235215 117623
rect 238769 117521 238803 117555
rect 238953 117453 238987 117487
rect 235181 117385 235215 117419
rect 240517 117725 240551 117759
rect 239505 117317 239539 117351
rect 239597 117521 239631 117555
rect 239597 117317 239631 117351
rect 244933 118269 244967 118303
rect 245853 118609 245887 118643
rect 248153 118609 248187 118643
rect 396825 118609 396859 118643
rect 244749 118201 244783 118235
rect 244749 117929 244783 117963
rect 242449 117521 242483 117555
rect 244565 117861 244599 117895
rect 249165 118541 249199 118575
rect 252845 118541 252879 118575
rect 248889 118201 248923 118235
rect 248981 118473 249015 118507
rect 249901 118269 249935 118303
rect 249257 118133 249291 118167
rect 249165 117861 249199 117895
rect 245853 117521 245887 117555
rect 249257 117521 249291 117555
rect 244565 117385 244599 117419
rect 246037 117453 246071 117487
rect 240517 117317 240551 117351
rect 250177 118133 250211 118167
rect 250453 118065 250487 118099
rect 334541 118473 334575 118507
rect 334909 118473 334943 118507
rect 389925 118405 389959 118439
rect 396825 118405 396859 118439
rect 398757 118609 398791 118643
rect 384313 118269 384347 118303
rect 252845 117997 252879 118031
rect 320741 118133 320775 118167
rect 315497 117861 315531 117895
rect 315497 117589 315531 117623
rect 315589 117861 315623 117895
rect 355333 118133 355367 118167
rect 320741 117589 320775 117623
rect 324881 118065 324915 118099
rect 315589 117453 315623 117487
rect 354413 118065 354447 118099
rect 336749 117861 336783 117895
rect 324881 117453 324915 117487
rect 325709 117725 325743 117759
rect 249901 117317 249935 117351
rect 246037 117249 246071 117283
rect 235089 117181 235123 117215
rect 186145 117113 186179 117147
rect 151829 116977 151863 117011
rect 133061 115889 133095 115923
rect 248337 115889 248371 115923
rect 131129 114529 131163 114563
rect 243737 114461 243771 114495
rect 73905 108953 73939 108987
rect 180993 113101 181027 113135
rect 131313 106233 131347 106267
rect 131313 99297 131347 99331
rect 133153 104805 133187 104839
rect 212641 110381 212675 110415
rect 194701 109701 194735 109735
rect 194701 104873 194735 104907
rect 180993 104737 181027 104771
rect 350457 117861 350491 117895
rect 350549 117793 350583 117827
rect 354413 117793 354447 117827
rect 398757 118269 398791 118303
rect 389833 118201 389867 118235
rect 384313 117997 384347 118031
rect 432613 117861 432647 117895
rect 355333 117793 355367 117827
rect 420745 117793 420779 117827
rect 340797 117725 340831 117759
rect 340889 117725 340923 117759
rect 413385 117725 413419 117759
rect 336749 117657 336783 117691
rect 413385 117521 413419 117555
rect 420745 117521 420779 117555
rect 422769 117793 422803 117827
rect 422769 117385 422803 117419
rect 426449 117793 426483 117827
rect 426541 117793 426575 117827
rect 426541 117521 426575 117555
rect 427829 117725 427863 117759
rect 427829 117521 427863 117555
rect 432613 117521 432647 117555
rect 432705 117861 432739 117895
rect 433533 117725 433567 117759
rect 444389 118541 444423 118575
rect 432705 117453 432739 117487
rect 434637 117453 434671 117487
rect 444389 117453 444423 117487
rect 456717 118541 456751 118575
rect 463801 118065 463835 118099
rect 456717 117453 456751 117487
rect 463709 117453 463743 117487
rect 476037 118065 476071 118099
rect 476037 117453 476071 117487
rect 492597 117657 492631 117691
rect 492597 117453 492631 117487
rect 492689 117589 492723 117623
rect 426449 117385 426483 117419
rect 425069 117249 425103 117283
rect 425069 117113 425103 117147
rect 434637 117113 434671 117147
rect 495357 117521 495391 117555
rect 495449 117521 495483 117555
rect 492689 116909 492723 116943
rect 325709 114529 325743 114563
rect 403909 115889 403943 115923
rect 248337 106301 248371 106335
rect 272257 114461 272291 114495
rect 243737 104873 243771 104907
rect 212641 100725 212675 100759
rect 233433 104805 233467 104839
rect 221105 100045 221139 100079
rect 133153 95217 133187 95251
rect 216689 99365 216723 99399
rect 156061 93789 156095 93823
rect 144929 90389 144963 90423
rect 73721 89845 73755 89879
rect 73721 86989 73755 87023
rect 144929 85561 144963 85595
rect 181177 92429 181211 92463
rect 156061 84201 156095 84235
rect 179521 88961 179555 88995
rect 179521 84201 179555 84235
rect 162869 84133 162903 84167
rect 157441 75837 157475 75871
rect 221105 95217 221139 95251
rect 227729 96577 227763 96611
rect 216689 91069 216723 91103
rect 207121 91001 207155 91035
rect 181177 82841 181211 82875
rect 190745 86921 190779 86955
rect 184857 77333 184891 77367
rect 190745 77265 190779 77299
rect 194885 85493 194919 85527
rect 184857 77129 184891 77163
rect 194885 75905 194919 75939
rect 200313 85493 200347 85527
rect 248245 104805 248279 104839
rect 243737 99365 243771 99399
rect 233433 95217 233467 95251
rect 238861 96577 238895 96611
rect 227729 89641 227763 89675
rect 243737 95217 243771 95251
rect 420469 115821 420503 115855
rect 420469 108953 420503 108987
rect 403909 106301 403943 106335
rect 272257 103513 272291 103547
rect 301973 106233 302007 106267
rect 301973 99297 302007 99331
rect 322673 106233 322707 106267
rect 394433 106233 394467 106267
rect 322673 99297 322707 99331
rect 325709 104805 325743 104839
rect 248245 95217 248279 95251
rect 431693 106233 431727 106267
rect 394433 99297 394467 99331
rect 415041 104805 415075 104839
rect 325709 95217 325743 95251
rect 383117 96577 383151 96611
rect 238861 89641 238895 89675
rect 279709 93789 279743 93823
rect 243737 86921 243771 86955
rect 233433 86853 233467 86887
rect 207121 81413 207155 81447
rect 227913 82093 227947 82127
rect 200313 75905 200347 75939
rect 205925 80121 205959 80155
rect 162869 74545 162903 74579
rect 183753 75837 183787 75871
rect 157441 66249 157475 66283
rect 174001 74477 174035 74511
rect 128921 66181 128955 66215
rect 174001 64889 174035 64923
rect 181085 73117 181119 73151
rect 145113 64821 145147 64855
rect 128921 57817 128955 57851
rect 133153 57885 133187 57919
rect 145113 56525 145147 56559
rect 147965 64821 147999 64855
rect 159097 64821 159131 64855
rect 147965 55233 147999 55267
rect 150725 57885 150759 57919
rect 133153 48297 133187 48331
rect 207213 80121 207247 80155
rect 221013 80121 221047 80155
rect 221013 79917 221047 79951
rect 227913 77265 227947 77299
rect 233433 77265 233467 77299
rect 238953 81413 238987 81447
rect 238953 77265 238987 77299
rect 243737 77265 243771 77299
rect 245761 86921 245795 86955
rect 274833 86921 274867 86955
rect 245761 77265 245795 77299
rect 248337 85493 248371 85527
rect 207213 76585 207247 76619
rect 383117 86989 383151 87023
rect 388637 96577 388671 96611
rect 388637 86989 388671 87023
rect 403909 96577 403943 96611
rect 415041 95217 415075 95251
rect 420653 104805 420687 104839
rect 431693 99297 431727 99331
rect 420653 95217 420687 95251
rect 403909 86989 403943 87023
rect 426173 95149 426207 95183
rect 279709 84269 279743 84303
rect 322673 86921 322707 86955
rect 274833 77265 274867 77299
rect 279709 84133 279743 84167
rect 248337 75905 248371 75939
rect 205925 74069 205959 74103
rect 211261 75837 211295 75871
rect 209881 70465 209915 70499
rect 209881 67609 209915 67643
rect 183753 66317 183787 66351
rect 244289 75837 244323 75871
rect 240241 70465 240275 70499
rect 211261 66249 211295 66283
rect 212733 68357 212767 68391
rect 181085 63529 181119 63563
rect 183753 66181 183787 66215
rect 159097 55233 159131 55267
rect 181177 61013 181211 61047
rect 195161 66181 195195 66215
rect 184949 60809 184983 60843
rect 184949 57885 184983 57919
rect 183753 56593 183787 56627
rect 207121 66181 207155 66215
rect 205833 60809 205867 60843
rect 205833 57953 205867 57987
rect 195161 56593 195195 56627
rect 200313 57885 200347 57919
rect 181177 50609 181211 50643
rect 184949 51085 184983 51119
rect 150725 48297 150759 48331
rect 184949 48297 184983 48331
rect 234721 67677 234755 67711
rect 233433 67541 233467 67575
rect 240241 67609 240275 67643
rect 234721 66249 234755 66283
rect 244289 66249 244323 66283
rect 245761 75837 245795 75871
rect 271889 75837 271923 75871
rect 394433 86921 394467 86955
rect 322673 77265 322707 77299
rect 325709 85493 325743 85527
rect 279709 74545 279743 74579
rect 301973 77129 302007 77163
rect 271889 70261 271923 70295
rect 358001 80121 358035 80155
rect 358001 79917 358035 79951
rect 426173 85561 426207 85595
rect 394433 77265 394467 77299
rect 426081 84133 426115 84167
rect 325709 75905 325743 75939
rect 341349 77129 341383 77163
rect 301973 67609 302007 67643
rect 341349 67609 341383 67643
rect 383209 77129 383243 77163
rect 383209 67609 383243 67643
rect 388729 77129 388763 77163
rect 388729 67609 388763 67643
rect 404001 77129 404035 77163
rect 426081 69649 426115 69683
rect 431601 75837 431635 75871
rect 404001 67609 404035 67643
rect 245761 66249 245795 66283
rect 431601 66249 431635 66283
rect 233433 62781 233467 62815
rect 248337 66181 248371 66215
rect 240149 58021 240183 58055
rect 207121 56593 207155 56627
rect 212549 57885 212583 57919
rect 212733 57885 212767 57919
rect 216873 57885 216907 57919
rect 200313 48297 200347 48331
rect 209881 51153 209915 51187
rect 73813 48229 73847 48263
rect 212549 51085 212583 51119
rect 240149 56593 240183 56627
rect 325525 66181 325559 66215
rect 248337 56593 248371 56627
rect 279893 57885 279927 57919
rect 234721 56525 234755 56559
rect 216873 48297 216907 48331
rect 227913 53125 227947 53159
rect 227913 48297 227947 48331
rect 209881 46937 209915 46971
rect 211261 46937 211295 46971
rect 234721 46937 234755 46971
rect 248337 48297 248371 48331
rect 279893 48297 279927 48331
rect 301789 57885 301823 57919
rect 301789 48297 301823 48331
rect 322673 57885 322707 57919
rect 415041 66181 415075 66215
rect 325525 56593 325559 56627
rect 383209 57885 383243 57919
rect 322673 48297 322707 48331
rect 341533 51153 341567 51187
rect 248337 46937 248371 46971
rect 157349 46869 157383 46903
rect 150817 41429 150851 41463
rect 73813 35309 73847 35343
rect 128921 38573 128955 38607
rect 133153 38573 133187 38607
rect 150817 38573 150851 38607
rect 190745 46869 190779 46903
rect 157349 37281 157383 37315
rect 181177 44081 181211 44115
rect 133153 31025 133187 31059
rect 150725 37213 150759 37247
rect 128921 28985 128955 29019
rect 181177 31637 181211 31671
rect 194701 46869 194735 46903
rect 276121 46869 276155 46903
rect 211261 45577 211295 45611
rect 238861 45849 238895 45883
rect 207213 45509 207247 45543
rect 194701 37281 194735 37315
rect 200405 38573 200439 38607
rect 190745 28985 190779 29019
rect 238861 41293 238895 41327
rect 325709 46869 325743 46903
rect 276121 37281 276155 37315
rect 322673 38573 322707 38607
rect 207213 35921 207247 35955
rect 234721 37213 234755 37247
rect 200405 28985 200439 29019
rect 229201 31841 229235 31875
rect 229201 28985 229235 29019
rect 150725 27625 150759 27659
rect 184949 28917 184983 28951
rect 157349 27557 157383 27591
rect 74273 20009 74307 20043
rect 74273 12325 74307 12359
rect 143641 19261 143675 19295
rect 143641 9673 143675 9707
rect 175565 26265 175599 26299
rect 175565 24837 175599 24871
rect 178049 25041 178083 25075
rect 178049 24701 178083 24735
rect 179429 24769 179463 24803
rect 174001 20009 174035 20043
rect 157349 9673 157383 9707
rect 168389 12461 168423 12495
rect 168389 9673 168423 9707
rect 168297 9605 168331 9639
rect 168481 9605 168515 9639
rect 168205 9537 168239 9571
rect 168205 9401 168239 9435
rect 125793 7157 125827 7191
rect 125793 7021 125827 7055
rect 178141 12325 178175 12359
rect 178141 9605 178175 9639
rect 174001 6885 174035 6919
rect 234721 27625 234755 27659
rect 238861 37213 238895 37247
rect 244289 37213 244323 37247
rect 245761 37213 245795 37247
rect 245761 31705 245795 31739
rect 248337 37213 248371 37247
rect 244289 31637 244323 31671
rect 238861 27625 238895 27659
rect 243737 27625 243771 27659
rect 248337 27625 248371 27659
rect 271889 37213 271923 37247
rect 383209 48297 383243 48331
rect 388729 57885 388763 57919
rect 388729 48297 388763 48331
rect 404001 57885 404035 57919
rect 415041 56593 415075 56627
rect 404001 48297 404035 48331
rect 341533 45577 341567 45611
rect 358001 48229 358035 48263
rect 341441 45441 341475 45475
rect 425989 46869 426023 46903
rect 358001 38641 358035 38675
rect 414949 45509 414983 45543
rect 341441 38233 341475 38267
rect 383209 38573 383243 38607
rect 325709 29053 325743 29087
rect 357725 29053 357759 29087
rect 322673 28985 322707 29019
rect 271889 27625 271923 27659
rect 279985 28917 280019 28951
rect 243737 26265 243771 26299
rect 276121 27557 276155 27591
rect 234629 22797 234663 22831
rect 205741 22185 205775 22219
rect 184949 19329 184983 19363
rect 190653 19397 190687 19431
rect 205741 19329 205775 19363
rect 233341 22117 233375 22151
rect 190653 17969 190687 18003
rect 200405 19261 200439 19295
rect 233341 19261 233375 19295
rect 234629 17969 234663 18003
rect 244565 19261 244599 19295
rect 200405 12257 200439 12291
rect 244565 11849 244599 11883
rect 274833 18105 274867 18139
rect 325709 27557 325743 27591
rect 279985 19329 280019 19363
rect 301881 26197 301915 26231
rect 276121 17969 276155 18003
rect 274833 9673 274867 9707
rect 183661 9605 183695 9639
rect 179429 6885 179463 6919
rect 183569 9469 183603 9503
rect 183569 6817 183603 6851
rect 383209 28985 383243 29019
rect 404001 38573 404035 38607
rect 425989 37281 426023 37315
rect 431601 46869 431635 46903
rect 431601 37281 431635 37315
rect 414949 35921 414983 35955
rect 431601 37145 431635 37179
rect 431601 31637 431635 31671
rect 404001 28985 404035 29019
rect 357725 26333 357759 26367
rect 420469 27557 420503 27591
rect 357909 26197 357943 26231
rect 415041 26197 415075 26231
rect 357909 21981 357943 22015
rect 383393 25245 383427 25279
rect 383393 19329 383427 19363
rect 394341 19261 394375 19295
rect 325709 9673 325743 9707
rect 383301 12529 383335 12563
rect 383301 9673 383335 9707
rect 420469 17969 420503 18003
rect 431509 26197 431543 26231
rect 415041 16609 415075 16643
rect 431509 16609 431543 16643
rect 394341 9673 394375 9707
rect 301881 8313 301915 8347
rect 414765 8245 414799 8279
rect 415041 8245 415075 8279
rect 412649 7565 412683 7599
rect 412649 7021 412683 7055
rect 183661 6069 183695 6103
rect 169677 4369 169711 4403
rect 205649 4369 205683 4403
rect 205649 4233 205683 4267
rect 67189 4165 67223 4199
rect 169677 4165 169711 4199
rect 62773 3281 62807 3315
rect 57989 3145 58023 3179
rect 57989 3009 58023 3043
rect 62773 3009 62807 3043
rect 507041 4097 507075 4131
rect 225061 4029 225095 4063
rect 220093 3961 220127 3995
rect 217977 3757 218011 3791
rect 196725 3621 196759 3655
rect 154589 3485 154623 3519
rect 147689 3417 147723 3451
rect 103529 3281 103563 3315
rect 103529 3009 103563 3043
rect 110613 3281 110647 3315
rect 110613 3009 110647 3043
rect 122849 3281 122883 3315
rect 122849 2805 122883 2839
rect 137937 3281 137971 3315
rect 147689 3281 147723 3315
rect 154589 3213 154623 3247
rect 164157 3485 164191 3519
rect 211169 3621 211203 3655
rect 210433 3553 210467 3587
rect 208869 3417 208903 3451
rect 196725 3349 196759 3383
rect 207673 3349 207707 3383
rect 164157 3213 164191 3247
rect 196633 3213 196667 3247
rect 195621 3145 195655 3179
rect 195621 2873 195655 2907
rect 137937 2805 137971 2839
rect 196633 2805 196667 2839
rect 202797 3009 202831 3043
rect 204453 3009 204487 3043
rect 207673 3009 207707 3043
rect 210341 3417 210375 3451
rect 210341 2941 210375 2975
rect 211169 3417 211203 3451
rect 210433 2941 210467 2975
rect 208869 2873 208903 2907
rect 219725 3757 219759 3791
rect 220093 3757 220127 3791
rect 361037 4029 361071 4063
rect 507317 4029 507351 4063
rect 225061 3689 225095 3723
rect 326445 3757 326479 3791
rect 219725 3485 219759 3519
rect 217977 2873 218011 2907
rect 204453 2805 204487 2839
rect 202797 1309 202831 1343
rect 67189 561 67223 595
rect 340153 3757 340187 3791
rect 340153 3553 340187 3587
rect 398849 3825 398883 3859
rect 398849 3621 398883 3655
rect 407405 3757 407439 3791
rect 361037 3553 361071 3587
rect 407405 3485 407439 3519
rect 417985 3621 418019 3655
rect 417985 3485 418019 3519
rect 418169 3485 418203 3519
rect 442273 3485 442307 3519
rect 432521 3417 432555 3451
rect 418261 2941 418295 2975
rect 422309 2941 422343 2975
rect 422309 2737 422343 2771
rect 437397 3417 437431 3451
rect 437397 2941 437431 2975
rect 496001 3349 496035 3383
rect 482385 3281 482419 3315
rect 485697 3281 485731 3315
rect 477877 3077 477911 3111
rect 478061 3077 478095 3111
rect 485145 3145 485179 3179
rect 482293 2941 482327 2975
rect 485053 2941 485087 2975
rect 485145 2941 485179 2975
rect 442273 2873 442307 2907
rect 484961 2873 484995 2907
rect 432521 2737 432555 2771
rect 489561 3281 489595 3315
rect 504373 3349 504407 3383
rect 496645 3213 496679 3247
rect 489101 3009 489135 3043
rect 489561 3009 489595 3043
rect 489837 3145 489871 3179
rect 504373 3145 504407 3179
rect 504465 3349 504499 3383
rect 513941 3349 513975 3383
rect 514033 4029 514067 4063
rect 514125 4029 514159 4063
rect 514033 3349 514067 3383
rect 504465 2941 504499 2975
rect 485697 2873 485731 2907
rect 485053 2805 485087 2839
rect 484961 2737 484995 2771
rect 326445 561 326479 595
<< metal1 >>
rect 133874 700952 133880 701004
rect 133932 700992 133938 701004
rect 267642 700992 267648 701004
rect 133932 700964 267648 700992
rect 133932 700952 133938 700964
rect 267642 700952 267648 700964
rect 267700 700952 267706 701004
rect 133782 700884 133788 700936
rect 133840 700924 133846 700936
rect 283834 700924 283840 700936
rect 133840 700896 283840 700924
rect 133840 700884 133846 700896
rect 283834 700884 283840 700896
rect 283892 700884 283898 700936
rect 300118 700884 300124 700936
rect 300176 700924 300182 700936
rect 434070 700924 434076 700936
rect 300176 700896 434076 700924
rect 300176 700884 300182 700896
rect 434070 700884 434076 700896
rect 434128 700884 434134 700936
rect 132494 700816 132500 700868
rect 132552 700856 132558 700868
rect 332502 700856 332508 700868
rect 132552 700828 332508 700856
rect 132552 700816 132558 700828
rect 332502 700816 332508 700828
rect 332560 700816 332566 700868
rect 133690 700748 133696 700800
rect 133748 700788 133754 700800
rect 218974 700788 218980 700800
rect 133748 700760 218980 700788
rect 133748 700748 133754 700760
rect 218974 700748 218980 700760
rect 219032 700748 219038 700800
rect 235166 700748 235172 700800
rect 235224 700788 235230 700800
rect 434162 700788 434168 700800
rect 235224 700760 434168 700788
rect 235224 700748 235230 700760
rect 434162 700748 434168 700760
rect 434220 700748 434226 700800
rect 131114 700680 131120 700732
rect 131172 700720 131178 700732
rect 348786 700720 348792 700732
rect 131172 700692 348792 700720
rect 131172 700680 131178 700692
rect 348786 700680 348792 700692
rect 348844 700680 348850 700732
rect 364978 700680 364984 700732
rect 365036 700720 365042 700732
rect 433978 700720 433984 700732
rect 365036 700692 433984 700720
rect 365036 700680 365042 700692
rect 433978 700680 433984 700692
rect 434036 700680 434042 700732
rect 170306 700612 170312 700664
rect 170364 700652 170370 700664
rect 434346 700652 434352 700664
rect 170364 700624 434352 700652
rect 170364 700612 170370 700624
rect 434346 700612 434352 700624
rect 434404 700612 434410 700664
rect 131206 700544 131212 700596
rect 131264 700584 131270 700596
rect 397454 700584 397460 700596
rect 131264 700556 397460 700584
rect 131264 700544 131270 700556
rect 397454 700544 397460 700556
rect 397512 700544 397518 700596
rect 132310 700476 132316 700528
rect 132368 700516 132374 700528
rect 413646 700516 413652 700528
rect 132368 700488 413652 700516
rect 132368 700476 132374 700488
rect 413646 700476 413652 700488
rect 413704 700476 413710 700528
rect 105446 700408 105452 700460
rect 105504 700448 105510 700460
rect 434438 700448 434444 700460
rect 105504 700420 434444 700448
rect 105504 700408 105510 700420
rect 434438 700408 434444 700420
rect 434496 700408 434502 700460
rect 438118 700408 438124 700460
rect 438176 700448 438182 700460
rect 494790 700448 494796 700460
rect 438176 700420 494796 700448
rect 438176 700408 438182 700420
rect 494790 700408 494796 700420
rect 494848 700408 494854 700460
rect 8110 700340 8116 700392
rect 8168 700380 8174 700392
rect 13078 700380 13084 700392
rect 8168 700352 13084 700380
rect 8168 700340 8174 700352
rect 13078 700340 13084 700352
rect 13136 700340 13142 700392
rect 89162 700340 89168 700392
rect 89220 700380 89226 700392
rect 126238 700380 126244 700392
rect 89220 700352 126244 700380
rect 89220 700340 89226 700352
rect 126238 700340 126244 700352
rect 126296 700340 126302 700392
rect 132586 700340 132592 700392
rect 132644 700380 132650 700392
rect 462314 700380 462320 700392
rect 132644 700352 462320 700380
rect 132644 700340 132650 700352
rect 462314 700340 462320 700352
rect 462372 700340 462378 700392
rect 40494 700272 40500 700324
rect 40552 700312 40558 700324
rect 434254 700312 434260 700324
rect 40552 700284 434260 700312
rect 40552 700272 40558 700284
rect 434254 700272 434260 700284
rect 434312 700272 434318 700324
rect 447778 700272 447784 700324
rect 447836 700312 447842 700324
rect 559650 700312 559656 700324
rect 447836 700284 559656 700312
rect 447836 700272 447842 700284
rect 559650 700272 559656 700284
rect 559708 700272 559714 700324
rect 133414 700204 133420 700256
rect 133472 700244 133478 700256
rect 202782 700244 202788 700256
rect 133472 700216 202788 700244
rect 133472 700204 133478 700216
rect 202782 700204 202788 700216
rect 202840 700204 202846 700256
rect 24302 699660 24308 699712
rect 24360 699700 24366 699712
rect 24762 699700 24768 699712
rect 24360 699672 24768 699700
rect 24360 699660 24366 699672
rect 24762 699660 24768 699672
rect 24820 699660 24826 699712
rect 72418 699660 72424 699712
rect 72476 699700 72482 699712
rect 72970 699700 72976 699712
rect 72476 699672 72976 699700
rect 72476 699660 72482 699672
rect 72970 699660 72976 699672
rect 73028 699660 73034 699712
rect 133322 699660 133328 699712
rect 133380 699700 133386 699712
rect 137830 699700 137836 699712
rect 133380 699672 137836 699700
rect 133380 699660 133386 699672
rect 137830 699660 137836 699672
rect 137888 699660 137894 699712
rect 429838 699660 429844 699712
rect 429896 699700 429902 699712
rect 433886 699700 433892 699712
rect 429896 699672 433892 699700
rect 429896 699660 429902 699672
rect 433886 699660 433892 699672
rect 433944 699660 433950 699712
rect 153562 698232 153568 698284
rect 153620 698272 153626 698284
rect 154206 698272 154212 698284
rect 153620 698244 154212 698272
rect 153620 698232 153626 698244
rect 154206 698232 154212 698244
rect 154264 698232 154270 698284
rect 147582 697076 147588 697128
rect 147640 697116 147646 697128
rect 154482 697116 154488 697128
rect 147640 697088 154488 697116
rect 147640 697076 147646 697088
rect 154482 697076 154488 697088
rect 154540 697076 154546 697128
rect 166902 697076 166908 697128
rect 166960 697116 166966 697128
rect 173802 697116 173808 697128
rect 166960 697088 173808 697116
rect 166960 697076 166966 697088
rect 173802 697076 173808 697088
rect 173860 697076 173866 697128
rect 186222 697076 186228 697128
rect 186280 697116 186286 697128
rect 193122 697116 193128 697128
rect 186280 697088 193128 697116
rect 186280 697076 186286 697088
rect 193122 697076 193128 697088
rect 193180 697076 193186 697128
rect 205542 697076 205548 697128
rect 205600 697116 205606 697128
rect 212442 697116 212448 697128
rect 205600 697088 212448 697116
rect 205600 697076 205606 697088
rect 212442 697076 212448 697088
rect 212500 697076 212506 697128
rect 224862 697076 224868 697128
rect 224920 697116 224926 697128
rect 231762 697116 231768 697128
rect 224920 697088 231768 697116
rect 224920 697076 224926 697088
rect 231762 697076 231768 697088
rect 231820 697076 231826 697128
rect 244182 697076 244188 697128
rect 244240 697116 244246 697128
rect 251082 697116 251088 697128
rect 244240 697088 251088 697116
rect 244240 697076 244246 697088
rect 251082 697076 251088 697088
rect 251140 697076 251146 697128
rect 263502 697076 263508 697128
rect 263560 697116 263566 697128
rect 270402 697116 270408 697128
rect 263560 697088 270408 697116
rect 263560 697076 263566 697088
rect 270402 697076 270408 697088
rect 270460 697076 270466 697128
rect 282822 697076 282828 697128
rect 282880 697116 282886 697128
rect 289722 697116 289728 697128
rect 282880 697088 289728 697116
rect 282880 697076 282886 697088
rect 289722 697076 289728 697088
rect 289780 697076 289786 697128
rect 302142 697076 302148 697128
rect 302200 697116 302206 697128
rect 309042 697116 309048 697128
rect 302200 697088 309048 697116
rect 302200 697076 302206 697088
rect 309042 697076 309048 697088
rect 309100 697076 309106 697128
rect 321462 697076 321468 697128
rect 321520 697116 321526 697128
rect 328362 697116 328368 697128
rect 321520 697088 328368 697116
rect 321520 697076 321526 697088
rect 328362 697076 328368 697088
rect 328420 697076 328426 697128
rect 154574 686264 154580 686316
rect 154632 686304 154638 686316
rect 159450 686304 159456 686316
rect 154632 686276 159456 686304
rect 154632 686264 154638 686276
rect 159450 686264 159456 686276
rect 159508 686264 159514 686316
rect 135254 686128 135260 686180
rect 135312 686168 135318 686180
rect 142890 686168 142896 686180
rect 135312 686140 142896 686168
rect 135312 686128 135318 686140
rect 142890 686128 142896 686140
rect 142948 686128 142954 686180
rect 153286 685924 153292 685976
rect 153344 685964 153350 685976
rect 153654 685964 153660 685976
rect 153344 685936 153660 685964
rect 153344 685924 153350 685936
rect 153654 685924 153660 685936
rect 153712 685924 153718 685976
rect 153286 684428 153292 684480
rect 153344 684468 153350 684480
rect 153565 684471 153623 684477
rect 153565 684468 153577 684471
rect 153344 684440 153577 684468
rect 153344 684428 153350 684440
rect 153565 684437 153577 684440
rect 153611 684437 153623 684471
rect 153565 684431 153623 684437
rect 3510 681708 3516 681760
rect 3568 681748 3574 681760
rect 434714 681748 434720 681760
rect 3568 681720 434720 681748
rect 3568 681708 3574 681720
rect 434714 681708 434720 681720
rect 434772 681708 434778 681760
rect 446398 673480 446404 673532
rect 446456 673520 446462 673532
rect 580166 673520 580172 673532
rect 446456 673492 580172 673520
rect 446456 673480 446462 673492
rect 580166 673480 580172 673492
rect 580224 673480 580230 673532
rect 3418 667904 3424 667956
rect 3476 667944 3482 667956
rect 19978 667944 19984 667956
rect 3476 667916 19984 667944
rect 3476 667904 3482 667916
rect 19978 667904 19984 667916
rect 20036 667904 20042 667956
rect 153565 666587 153623 666593
rect 153565 666553 153577 666587
rect 153611 666584 153623 666587
rect 153654 666584 153660 666596
rect 153611 666556 153660 666584
rect 153611 666553 153623 666556
rect 153565 666547 153623 666553
rect 153654 666544 153660 666556
rect 153712 666544 153718 666596
rect 153470 656860 153476 656872
rect 153431 656832 153476 656860
rect 153470 656820 153476 656832
rect 153528 656820 153534 656872
rect 154574 650360 154580 650412
rect 154632 650400 154638 650412
rect 159450 650400 159456 650412
rect 154632 650372 159456 650400
rect 154632 650360 154638 650372
rect 159450 650360 159456 650372
rect 159508 650360 159514 650412
rect 135254 650224 135260 650276
rect 135312 650264 135318 650276
rect 142890 650264 142896 650276
rect 135312 650236 142896 650264
rect 135312 650224 135318 650236
rect 142890 650224 142896 650236
rect 142948 650224 142954 650276
rect 153473 647275 153531 647281
rect 153473 647241 153485 647275
rect 153519 647272 153531 647275
rect 153562 647272 153568 647284
rect 153519 647244 153568 647272
rect 153519 647241 153531 647244
rect 153473 647235 153531 647241
rect 153562 647232 153568 647244
rect 153620 647232 153626 647284
rect 153289 645847 153347 645853
rect 153289 645813 153301 645847
rect 153335 645844 153347 645847
rect 153562 645844 153568 645856
rect 153335 645816 153568 645844
rect 153335 645813 153347 645816
rect 153289 645807 153347 645813
rect 153562 645804 153568 645816
rect 153620 645804 153626 645856
rect 153286 636256 153292 636268
rect 153247 636228 153292 636256
rect 153286 636216 153292 636228
rect 153344 636216 153350 636268
rect 153286 630504 153292 630556
rect 153344 630544 153350 630556
rect 153562 630544 153568 630556
rect 153344 630516 153568 630544
rect 153344 630504 153350 630516
rect 153562 630504 153568 630516
rect 153620 630504 153626 630556
rect 445018 626560 445024 626612
rect 445076 626600 445082 626612
rect 580166 626600 580172 626612
rect 445076 626572 580172 626600
rect 445076 626560 445082 626572
rect 580166 626560 580172 626572
rect 580224 626560 580230 626612
rect 3418 623772 3424 623824
rect 3476 623812 3482 623824
rect 434806 623812 434812 623824
rect 3476 623784 434812 623812
rect 3476 623772 3482 623784
rect 434806 623772 434812 623784
rect 434864 623772 434870 623824
rect 153562 621092 153568 621104
rect 153488 621064 153568 621092
rect 153488 620968 153516 621064
rect 153562 621052 153568 621064
rect 153620 621052 153626 621104
rect 153470 620916 153476 620968
rect 153528 620916 153534 620968
rect 3418 609968 3424 610020
rect 3476 610008 3482 610020
rect 21358 610008 21364 610020
rect 3476 609980 21364 610008
rect 3476 609968 3482 609980
rect 21358 609968 21364 609980
rect 21416 609968 21422 610020
rect 153286 598924 153292 598936
rect 153247 598896 153292 598924
rect 153286 598884 153292 598896
rect 153344 598884 153350 598936
rect 4062 594804 4068 594856
rect 4120 594844 4126 594856
rect 4890 594844 4896 594856
rect 4120 594816 4896 594844
rect 4120 594804 4126 594816
rect 4890 594804 4896 594816
rect 4948 594804 4954 594856
rect 154574 592424 154580 592476
rect 154632 592464 154638 592476
rect 159450 592464 159456 592476
rect 154632 592436 159456 592464
rect 154632 592424 154638 592436
rect 159450 592424 159456 592436
rect 159508 592424 159514 592476
rect 135254 592288 135260 592340
rect 135312 592328 135318 592340
rect 142890 592328 142896 592340
rect 135312 592300 142896 592328
rect 135312 592288 135318 592300
rect 142890 592288 142896 592300
rect 142948 592288 142954 592340
rect 153289 589339 153347 589345
rect 153289 589305 153301 589339
rect 153335 589336 153347 589339
rect 153470 589336 153476 589348
rect 153335 589308 153476 589336
rect 153335 589305 153347 589308
rect 153289 589299 153347 589305
rect 153470 589296 153476 589308
rect 153528 589296 153534 589348
rect 270402 583652 270408 583704
rect 270460 583692 270466 583704
rect 307018 583692 307024 583704
rect 270460 583664 307024 583692
rect 270460 583652 270466 583664
rect 307018 583652 307024 583664
rect 307076 583652 307082 583704
rect 287698 583584 287704 583636
rect 287756 583624 287762 583636
rect 319714 583624 319720 583636
rect 287756 583596 319720 583624
rect 287756 583584 287762 583596
rect 319714 583584 319720 583596
rect 319772 583584 319778 583636
rect 130378 583516 130384 583568
rect 130436 583556 130442 583568
rect 311250 583556 311256 583568
rect 130436 583528 311256 583556
rect 130436 583516 130442 583528
rect 311250 583516 311256 583528
rect 311308 583516 311314 583568
rect 128998 583448 129004 583500
rect 129056 583488 129062 583500
rect 330386 583488 330392 583500
rect 129056 583460 330392 583488
rect 129056 583448 129062 583460
rect 330386 583448 330392 583460
rect 330444 583448 330450 583500
rect 129274 583380 129280 583432
rect 129332 583420 129338 583432
rect 347498 583420 347504 583432
rect 129332 583392 347504 583420
rect 129332 583380 129338 583392
rect 347498 583380 347504 583392
rect 347556 583380 347562 583432
rect 119338 583312 119344 583364
rect 119396 583352 119402 583364
rect 336826 583352 336832 583364
rect 119396 583324 336832 583352
rect 119396 583312 119402 583324
rect 336826 583312 336832 583324
rect 336884 583312 336890 583364
rect 85390 583244 85396 583296
rect 85448 583284 85454 583296
rect 334618 583284 334624 583296
rect 85448 583256 334624 583284
rect 85448 583244 85454 583256
rect 334618 583244 334624 583256
rect 334676 583244 334682 583296
rect 298462 583176 298468 583228
rect 298520 583216 298526 583228
rect 332594 583216 332600 583228
rect 298520 583188 332600 583216
rect 298520 583176 298526 583188
rect 332594 583176 332600 583188
rect 332652 583176 332658 583228
rect 298370 583108 298376 583160
rect 298428 583148 298434 583160
rect 341058 583148 341064 583160
rect 298428 583120 341064 583148
rect 298428 583108 298434 583120
rect 341058 583108 341064 583120
rect 341116 583108 341122 583160
rect 293862 583040 293868 583092
rect 293920 583080 293926 583092
rect 338850 583080 338856 583092
rect 293920 583052 338856 583080
rect 293920 583040 293926 583052
rect 338850 583040 338856 583052
rect 338908 583040 338914 583092
rect 281442 582972 281448 583024
rect 281500 583012 281506 583024
rect 326154 583012 326160 583024
rect 281500 582984 326160 583012
rect 281500 582972 281506 582984
rect 326154 582972 326160 582984
rect 326212 582972 326218 583024
rect 298278 582904 298284 582956
rect 298336 582944 298342 582956
rect 353754 582944 353760 582956
rect 298336 582916 353760 582944
rect 298336 582904 298342 582916
rect 353754 582904 353760 582916
rect 353812 582904 353818 582956
rect 298554 582836 298560 582888
rect 298612 582876 298618 582888
rect 355962 582876 355968 582888
rect 298612 582848 355968 582876
rect 298612 582836 298618 582848
rect 355962 582836 355968 582848
rect 356020 582836 356026 582888
rect 291102 582768 291108 582820
rect 291160 582808 291166 582820
rect 351730 582808 351736 582820
rect 291160 582780 351736 582808
rect 291160 582768 291166 582780
rect 351730 582768 351736 582780
rect 351788 582768 351794 582820
rect 300486 582700 300492 582752
rect 300544 582740 300550 582752
rect 362402 582740 362408 582752
rect 300544 582712 362408 582740
rect 300544 582700 300550 582712
rect 362402 582700 362408 582712
rect 362460 582700 362466 582752
rect 298186 582632 298192 582684
rect 298244 582672 298250 582684
rect 345290 582672 345296 582684
rect 298244 582644 345296 582672
rect 298244 582632 298250 582644
rect 345290 582632 345296 582644
rect 345348 582632 345354 582684
rect 366634 582632 366640 582684
rect 366692 582672 366698 582684
rect 378226 582672 378232 582684
rect 366692 582644 378232 582672
rect 366692 582632 366698 582644
rect 378226 582632 378232 582644
rect 378284 582632 378290 582684
rect 294598 582564 294604 582616
rect 294656 582604 294662 582616
rect 313458 582604 313464 582616
rect 294656 582576 313464 582604
rect 294656 582564 294662 582576
rect 313458 582564 313464 582576
rect 313516 582564 313522 582616
rect 357986 582564 357992 582616
rect 358044 582604 358050 582616
rect 378410 582604 378416 582616
rect 358044 582576 378416 582604
rect 358044 582564 358050 582576
rect 378410 582564 378416 582576
rect 378468 582564 378474 582616
rect 298646 582496 298652 582548
rect 298704 582536 298710 582548
rect 321922 582536 321928 582548
rect 298704 582508 321928 582536
rect 298704 582496 298710 582508
rect 321922 582496 321928 582508
rect 321980 582496 321986 582548
rect 370866 582496 370872 582548
rect 370924 582536 370930 582548
rect 378594 582536 378600 582548
rect 370924 582508 378600 582536
rect 370924 582496 370930 582508
rect 378594 582496 378600 582508
rect 378652 582496 378658 582548
rect 298738 582428 298744 582480
rect 298796 582468 298802 582480
rect 328362 582468 328368 582480
rect 298796 582440 328368 582468
rect 298796 582428 298802 582440
rect 328362 582428 328368 582440
rect 328420 582428 328426 582480
rect 300394 582360 300400 582412
rect 300452 582400 300458 582412
rect 309226 582400 309232 582412
rect 300452 582372 309232 582400
rect 300452 582360 300458 582372
rect 309226 582360 309232 582372
rect 309284 582360 309290 582412
rect 372890 582360 372896 582412
rect 372948 582400 372954 582412
rect 378502 582400 378508 582412
rect 372948 582372 378508 582400
rect 372948 582360 372954 582372
rect 378502 582360 378508 582372
rect 378560 582360 378566 582412
rect 153378 579640 153384 579692
rect 153436 579680 153442 579692
rect 153470 579680 153476 579692
rect 153436 579652 153476 579680
rect 153436 579640 153442 579652
rect 153470 579640 153476 579652
rect 153528 579640 153534 579692
rect 299382 579640 299388 579692
rect 299440 579680 299446 579692
rect 304810 579680 304816 579692
rect 299440 579652 304816 579680
rect 299440 579640 299446 579652
rect 304810 579640 304816 579652
rect 304868 579640 304874 579692
rect 442258 579640 442264 579692
rect 442316 579680 442322 579692
rect 580166 579680 580172 579692
rect 442316 579652 580172 579680
rect 442316 579640 442322 579652
rect 580166 579640 580172 579652
rect 580224 579640 580230 579692
rect 299474 579300 299480 579352
rect 299532 579340 299538 579352
rect 300670 579340 300676 579352
rect 299532 579312 300676 579340
rect 299532 579300 299538 579312
rect 300670 579300 300676 579312
rect 300728 579300 300734 579352
rect 315206 579340 315212 579352
rect 315167 579312 315212 579340
rect 315206 579300 315212 579312
rect 315264 579300 315270 579352
rect 317414 579340 317420 579352
rect 317375 579312 317420 579340
rect 317414 579300 317420 579312
rect 317472 579300 317478 579352
rect 342990 579340 342996 579352
rect 342951 579312 342996 579340
rect 342990 579300 342996 579312
rect 343048 579300 343054 579352
rect 364242 579340 364248 579352
rect 364203 579312 364248 579340
rect 364242 579300 364248 579312
rect 364300 579300 364306 579352
rect 375374 579300 375380 579352
rect 375432 579340 375438 579352
rect 378318 579340 378324 579352
rect 375432 579312 378324 579340
rect 375432 579300 375438 579312
rect 378318 579300 378324 579312
rect 378376 579300 378382 579352
rect 122742 578416 122748 578468
rect 122800 578456 122806 578468
rect 315209 578459 315267 578465
rect 315209 578456 315221 578459
rect 122800 578428 315221 578456
rect 122800 578416 122806 578428
rect 315209 578425 315221 578428
rect 315255 578425 315267 578459
rect 315209 578419 315267 578425
rect 115382 578348 115388 578400
rect 115440 578388 115446 578400
rect 317417 578391 317475 578397
rect 317417 578388 317429 578391
rect 115440 578360 317429 578388
rect 115440 578348 115446 578360
rect 317417 578357 317429 578360
rect 317463 578357 317475 578391
rect 317417 578351 317475 578357
rect 115198 578280 115204 578332
rect 115256 578320 115262 578332
rect 342993 578323 343051 578329
rect 342993 578320 343005 578323
rect 115256 578292 343005 578320
rect 115256 578280 115262 578292
rect 342993 578289 343005 578292
rect 343039 578289 343051 578323
rect 342993 578283 343051 578289
rect 129182 578212 129188 578264
rect 129240 578252 129246 578264
rect 364245 578255 364303 578261
rect 364245 578252 364257 578255
rect 129240 578224 364257 578252
rect 129240 578212 129246 578224
rect 364245 578221 364257 578224
rect 364291 578221 364303 578255
rect 364245 578215 364303 578221
rect 110322 575492 110328 575544
rect 110380 575532 110386 575544
rect 298002 575532 298008 575544
rect 110380 575504 298008 575532
rect 110380 575492 110386 575504
rect 298002 575492 298008 575504
rect 298060 575492 298066 575544
rect 272518 569916 272524 569968
rect 272576 569956 272582 569968
rect 298002 569956 298008 569968
rect 272576 569928 298008 569956
rect 272576 569916 272582 569928
rect 298002 569916 298008 569928
rect 298060 569916 298066 569968
rect 129642 563048 129648 563100
rect 129700 563088 129706 563100
rect 296898 563088 296904 563100
rect 129700 563060 296904 563088
rect 129700 563048 129706 563060
rect 296898 563048 296904 563060
rect 296956 563048 296962 563100
rect 196176 562108 210464 562136
rect 196176 562068 196204 562108
rect 195992 562040 196204 562068
rect 195882 561960 195888 562012
rect 195940 562000 195946 562012
rect 195992 562000 196020 562040
rect 195940 561972 196020 562000
rect 195940 561960 195946 561972
rect 197078 561892 197084 561944
rect 197136 561932 197142 561944
rect 208670 561932 208676 561944
rect 197136 561904 208676 561932
rect 197136 561892 197142 561904
rect 208670 561892 208676 561904
rect 208728 561892 208734 561944
rect 210436 561932 210464 562108
rect 217870 561932 217876 561944
rect 210436 561904 217876 561932
rect 217870 561892 217876 561904
rect 217928 561892 217934 561944
rect 197262 561824 197268 561876
rect 197320 561864 197326 561876
rect 214742 561864 214748 561876
rect 197320 561836 214748 561864
rect 197320 561824 197326 561836
rect 214742 561824 214748 561836
rect 214800 561824 214806 561876
rect 196986 561756 196992 561808
rect 197044 561796 197050 561808
rect 202414 561796 202420 561808
rect 197044 561768 202420 561796
rect 197044 561756 197050 561768
rect 202414 561756 202420 561768
rect 202472 561756 202478 561808
rect 197170 561688 197176 561740
rect 197228 561728 197234 561740
rect 205542 561728 205548 561740
rect 197228 561700 205548 561728
rect 197228 561688 197234 561700
rect 205542 561688 205548 561700
rect 205600 561688 205606 561740
rect 153286 560260 153292 560312
rect 153344 560300 153350 560312
rect 153378 560300 153384 560312
rect 153344 560272 153384 560300
rect 153344 560260 153350 560272
rect 153378 560260 153384 560272
rect 153436 560260 153442 560312
rect 391198 556248 391204 556300
rect 391256 556288 391262 556300
rect 484394 556288 484400 556300
rect 391256 556260 484400 556288
rect 391256 556248 391262 556260
rect 484394 556248 484400 556260
rect 484452 556248 484458 556300
rect 273162 556180 273168 556232
rect 273220 556220 273226 556232
rect 297266 556220 297272 556232
rect 273220 556192 297272 556220
rect 273220 556180 273226 556192
rect 297266 556180 297272 556192
rect 297324 556180 297330 556232
rect 395338 556180 395344 556232
rect 395396 556220 395402 556232
rect 511258 556220 511264 556232
rect 395396 556192 511264 556220
rect 395396 556180 395402 556192
rect 511258 556180 511264 556192
rect 511316 556180 511322 556232
rect 109402 554752 109408 554804
rect 109460 554792 109466 554804
rect 110322 554792 110328 554804
rect 109460 554764 110328 554792
rect 109460 554752 109466 554764
rect 110322 554752 110328 554764
rect 110380 554792 110386 554804
rect 115934 554792 115940 554804
rect 110380 554764 115940 554792
rect 110380 554752 110386 554764
rect 115934 554752 115940 554764
rect 115992 554752 115998 554804
rect 92106 553936 92112 553988
rect 92164 553976 92170 553988
rect 115290 553976 115296 553988
rect 92164 553948 115296 553976
rect 92164 553936 92170 553948
rect 115290 553936 115296 553948
rect 115348 553936 115354 553988
rect 89162 553868 89168 553920
rect 89220 553908 89226 553920
rect 160738 553908 160744 553920
rect 89220 553880 160744 553908
rect 89220 553868 89226 553880
rect 160738 553868 160744 553880
rect 160796 553868 160802 553920
rect 115106 553800 115112 553852
rect 115164 553840 115170 553852
rect 128354 553840 128360 553852
rect 115164 553812 128360 553840
rect 115164 553800 115170 553812
rect 128354 553800 128360 553812
rect 128412 553840 128418 553852
rect 129274 553840 129280 553852
rect 128412 553812 129280 553840
rect 128412 553800 128418 553812
rect 129274 553800 129280 553812
rect 129332 553800 129338 553852
rect 95050 553732 95056 553784
rect 95108 553772 95114 553784
rect 120718 553772 120724 553784
rect 95108 553744 120724 553772
rect 95108 553732 95114 553744
rect 120718 553732 120724 553744
rect 120776 553732 120782 553784
rect 100754 553664 100760 553716
rect 100812 553704 100818 553716
rect 129090 553704 129096 553716
rect 100812 553676 129096 553704
rect 100812 553664 100818 553676
rect 129090 553664 129096 553676
rect 129148 553664 129154 553716
rect 106458 553596 106464 553648
rect 106516 553636 106522 553648
rect 140038 553636 140044 553648
rect 106516 553608 140044 553636
rect 106516 553596 106522 553608
rect 140038 553596 140044 553608
rect 140096 553596 140102 553648
rect 103698 553528 103704 553580
rect 103756 553568 103762 553580
rect 146938 553568 146944 553580
rect 103756 553540 146944 553568
rect 103756 553528 103762 553540
rect 146938 553528 146944 553540
rect 146996 553528 147002 553580
rect 97810 553460 97816 553512
rect 97868 553500 97874 553512
rect 153838 553500 153844 553512
rect 97868 553472 153844 553500
rect 97868 553460 97874 553472
rect 153838 553460 153844 553472
rect 153896 553460 153902 553512
rect 112346 553392 112352 553444
rect 112404 553432 112410 553444
rect 116026 553432 116032 553444
rect 112404 553404 116032 553432
rect 112404 553392 112410 553404
rect 116026 553392 116032 553404
rect 116084 553392 116090 553444
rect 3142 552032 3148 552084
rect 3200 552072 3206 552084
rect 28258 552072 28264 552084
rect 3200 552044 28264 552072
rect 3200 552032 3206 552044
rect 28258 552032 28264 552044
rect 28316 552032 28322 552084
rect 85482 549856 85488 549908
rect 85540 549896 85546 549908
rect 86402 549896 86408 549908
rect 85540 549868 86408 549896
rect 85540 549856 85546 549868
rect 86402 549856 86408 549868
rect 86460 549896 86466 549908
rect 115382 549896 115388 549908
rect 86460 549868 115388 549896
rect 86460 549856 86466 549868
rect 115382 549856 115388 549868
rect 115440 549856 115446 549908
rect 118602 542376 118608 542428
rect 118660 542416 118666 542428
rect 152458 542416 152464 542428
rect 118660 542388 152464 542416
rect 118660 542376 118666 542388
rect 152458 542376 152464 542388
rect 152516 542376 152522 542428
rect 286962 538228 286968 538280
rect 287020 538268 287026 538280
rect 297634 538268 297640 538280
rect 287020 538240 297640 538268
rect 287020 538228 287026 538240
rect 297634 538228 297640 538240
rect 297692 538228 297698 538280
rect 117774 536800 117780 536852
rect 117832 536840 117838 536852
rect 144178 536840 144184 536852
rect 117832 536812 144184 536840
rect 117832 536800 117838 536812
rect 144178 536800 144184 536812
rect 144236 536800 144242 536852
rect 296070 534012 296076 534064
rect 296128 534052 296134 534064
rect 297450 534052 297456 534064
rect 296128 534024 297456 534052
rect 296128 534012 296134 534024
rect 297450 534012 297456 534024
rect 297508 534012 297514 534064
rect 117774 532720 117780 532772
rect 117832 532760 117838 532772
rect 159358 532760 159364 532772
rect 117832 532732 159364 532760
rect 117832 532720 117838 532732
rect 159358 532720 159364 532732
rect 159416 532720 159422 532772
rect 514018 532720 514024 532772
rect 514076 532760 514082 532772
rect 580166 532760 580172 532772
rect 514076 532732 580172 532760
rect 514076 532720 514082 532732
rect 580166 532720 580172 532732
rect 580224 532720 580230 532772
rect 153378 531292 153384 531344
rect 153436 531332 153442 531344
rect 153470 531332 153476 531344
rect 153436 531304 153476 531332
rect 153436 531292 153442 531304
rect 153470 531292 153476 531304
rect 153528 531292 153534 531344
rect 117958 529864 117964 529916
rect 118016 529904 118022 529916
rect 119338 529904 119344 529916
rect 118016 529876 119344 529904
rect 118016 529864 118022 529876
rect 119338 529864 119344 529876
rect 119396 529864 119402 529916
rect 118602 525036 118608 525088
rect 118660 525076 118666 525088
rect 128722 525076 128728 525088
rect 118660 525048 128728 525076
rect 118660 525036 118666 525048
rect 128722 525036 128728 525048
rect 128780 525036 128786 525088
rect 128722 524764 128728 524816
rect 128780 524804 128786 524816
rect 129182 524804 129188 524816
rect 128780 524776 129188 524804
rect 128780 524764 128786 524776
rect 129182 524764 129188 524776
rect 129240 524764 129246 524816
rect 70118 524424 70124 524476
rect 70176 524464 70182 524476
rect 82814 524464 82820 524476
rect 70176 524436 82820 524464
rect 70176 524424 70182 524436
rect 82814 524424 82820 524436
rect 82872 524424 82878 524476
rect 153378 524424 153384 524476
rect 153436 524424 153442 524476
rect 153396 524396 153424 524424
rect 153470 524396 153476 524408
rect 153396 524368 153476 524396
rect 153470 524356 153476 524368
rect 153528 524356 153534 524408
rect 280062 521636 280068 521688
rect 280120 521676 280126 521688
rect 297174 521676 297180 521688
rect 280120 521648 297180 521676
rect 280120 521636 280126 521648
rect 297174 521636 297180 521648
rect 297232 521636 297238 521688
rect 128446 521568 128452 521620
rect 128504 521608 128510 521620
rect 128998 521608 129004 521620
rect 128504 521580 129004 521608
rect 128504 521568 128510 521580
rect 128998 521568 129004 521580
rect 129056 521568 129062 521620
rect 295334 521568 295340 521620
rect 295392 521608 295398 521620
rect 296070 521608 296076 521620
rect 295392 521580 296076 521608
rect 295392 521568 295398 521580
rect 296070 521568 296076 521580
rect 296128 521568 296134 521620
rect 85206 521228 85212 521280
rect 85264 521268 85270 521280
rect 295334 521268 295340 521280
rect 85264 521240 295340 521268
rect 85264 521228 85270 521240
rect 295334 521228 295340 521240
rect 295392 521228 295398 521280
rect 199378 521160 199384 521212
rect 199436 521200 199442 521212
rect 222378 521200 222384 521212
rect 199436 521172 222384 521200
rect 199436 521160 199442 521172
rect 222378 521160 222384 521172
rect 222436 521160 222442 521212
rect 199470 521092 199476 521144
rect 199528 521132 199534 521144
rect 222562 521132 222568 521144
rect 199528 521104 222568 521132
rect 199528 521092 199534 521104
rect 222562 521092 222568 521104
rect 222620 521092 222626 521144
rect 198182 521024 198188 521076
rect 198240 521064 198246 521076
rect 222654 521064 222660 521076
rect 198240 521036 222660 521064
rect 198240 521024 198246 521036
rect 222654 521024 222660 521036
rect 222712 521024 222718 521076
rect 117314 520956 117320 521008
rect 117372 520996 117378 521008
rect 128446 520996 128452 521008
rect 117372 520968 128452 520996
rect 117372 520956 117378 520968
rect 128446 520956 128452 520968
rect 128504 520956 128510 521008
rect 198274 520956 198280 521008
rect 198332 520996 198338 521008
rect 222470 520996 222476 521008
rect 198332 520968 222476 520996
rect 198332 520956 198338 520968
rect 222470 520956 222476 520968
rect 222528 520956 222534 521008
rect 85298 520888 85304 520940
rect 85356 520928 85362 520940
rect 295978 520928 295984 520940
rect 85356 520900 295984 520928
rect 85356 520888 85362 520900
rect 295978 520888 295984 520900
rect 296036 520928 296042 520940
rect 298186 520928 298192 520940
rect 296036 520900 298192 520928
rect 296036 520888 296042 520900
rect 298186 520888 298192 520900
rect 298244 520888 298250 520940
rect 279418 518916 279424 518968
rect 279476 518956 279482 518968
rect 297266 518956 297272 518968
rect 279476 518928 297272 518956
rect 279476 518916 279482 518928
rect 297266 518916 297272 518928
rect 297324 518916 297330 518968
rect 89346 518848 89352 518900
rect 89404 518888 89410 518900
rect 130378 518888 130384 518900
rect 89404 518860 130384 518888
rect 89404 518848 89410 518860
rect 130378 518848 130384 518860
rect 130436 518848 130442 518900
rect 109586 518780 109592 518832
rect 109644 518820 109650 518832
rect 113174 518820 113180 518832
rect 109644 518792 113180 518820
rect 109644 518780 109650 518792
rect 113174 518780 113180 518792
rect 113232 518820 113238 518832
rect 115198 518820 115204 518832
rect 113232 518792 115204 518820
rect 113232 518780 113238 518792
rect 115198 518780 115204 518792
rect 115256 518780 115262 518832
rect 127710 518820 127716 518832
rect 122852 518792 127716 518820
rect 86586 518712 86592 518764
rect 86644 518752 86650 518764
rect 99285 518755 99343 518761
rect 99285 518752 99297 518755
rect 86644 518724 99297 518752
rect 86644 518712 86650 518724
rect 99285 518721 99297 518724
rect 99331 518721 99343 518755
rect 99285 518715 99343 518721
rect 118697 518755 118755 518761
rect 118697 518721 118709 518755
rect 118743 518752 118755 518755
rect 122742 518752 122748 518764
rect 118743 518724 122748 518752
rect 118743 518721 118755 518724
rect 118697 518715 118755 518721
rect 122742 518712 122748 518724
rect 122800 518752 122806 518764
rect 122852 518752 122880 518792
rect 127710 518780 127716 518792
rect 127768 518780 127774 518832
rect 122800 518724 122880 518752
rect 122800 518712 122806 518724
rect 99377 518687 99435 518693
rect 99377 518653 99389 518687
rect 99423 518684 99435 518687
rect 115845 518687 115903 518693
rect 99423 518656 99512 518684
rect 99423 518653 99435 518656
rect 99377 518647 99435 518653
rect 99484 518616 99512 518656
rect 115845 518653 115857 518687
rect 115891 518684 115903 518687
rect 118513 518687 118571 518693
rect 118513 518684 118525 518687
rect 115891 518656 118525 518684
rect 115891 518653 115903 518656
rect 115845 518647 115903 518653
rect 118513 518653 118525 518656
rect 118559 518653 118571 518687
rect 118513 518647 118571 518653
rect 106277 518619 106335 518625
rect 106277 518616 106289 518619
rect 99484 518588 106289 518616
rect 106277 518585 106289 518588
rect 106323 518585 106335 518619
rect 106277 518579 106335 518585
rect 106277 518483 106335 518489
rect 106277 518449 106289 518483
rect 106323 518480 106335 518483
rect 115845 518483 115903 518489
rect 115845 518480 115857 518483
rect 106323 518452 115857 518480
rect 106323 518449 106335 518452
rect 106277 518443 106335 518449
rect 115845 518449 115857 518452
rect 115891 518449 115903 518483
rect 115845 518443 115903 518449
rect 97994 518372 98000 518424
rect 98052 518412 98058 518424
rect 126330 518412 126336 518424
rect 98052 518384 126336 518412
rect 98052 518372 98058 518384
rect 126330 518372 126336 518384
rect 126388 518372 126394 518424
rect 106642 518304 106648 518356
rect 106700 518344 106706 518356
rect 151078 518344 151084 518356
rect 106700 518316 151084 518344
rect 106700 518304 106706 518316
rect 151078 518304 151084 518316
rect 151136 518304 151142 518356
rect 100938 518236 100944 518288
rect 100996 518276 101002 518288
rect 157978 518276 157984 518288
rect 100996 518248 157984 518276
rect 100996 518236 101002 518248
rect 157978 518236 157984 518248
rect 158036 518236 158042 518288
rect 198090 518236 198096 518288
rect 198148 518276 198154 518288
rect 218974 518276 218980 518288
rect 198148 518248 218980 518276
rect 198148 518236 198154 518248
rect 218974 518236 218980 518248
rect 219032 518236 219038 518288
rect 391290 518236 391296 518288
rect 391348 518276 391354 518288
rect 479978 518276 479984 518288
rect 391348 518248 479984 518276
rect 391348 518236 391354 518248
rect 479978 518236 479984 518248
rect 480036 518236 480042 518288
rect 92290 518168 92296 518220
rect 92348 518208 92354 518220
rect 126974 518208 126980 518220
rect 92348 518180 126980 518208
rect 92348 518168 92354 518180
rect 126974 518168 126980 518180
rect 127032 518208 127038 518220
rect 297450 518208 297456 518220
rect 127032 518180 297456 518208
rect 127032 518168 127038 518180
rect 297450 518168 297456 518180
rect 297508 518168 297514 518220
rect 398098 518168 398104 518220
rect 398156 518208 398162 518220
rect 506842 518208 506848 518220
rect 398156 518180 506848 518208
rect 398156 518168 398162 518180
rect 506842 518168 506848 518180
rect 506900 518168 506906 518220
rect 205634 517488 205640 517540
rect 205692 517528 205698 517540
rect 206646 517528 206652 517540
rect 205692 517500 206652 517528
rect 205692 517488 205698 517500
rect 206646 517488 206652 517500
rect 206704 517488 206710 517540
rect 284938 516128 284944 516180
rect 284996 516168 285002 516180
rect 297818 516168 297824 516180
rect 284996 516140 297824 516168
rect 284996 516128 285002 516140
rect 297818 516128 297824 516140
rect 297876 516128 297882 516180
rect 153286 511980 153292 512032
rect 153344 512020 153350 512032
rect 153562 512020 153568 512032
rect 153344 511992 153568 512020
rect 153344 511980 153350 511992
rect 153562 511980 153568 511992
rect 153620 511980 153626 512032
rect 294690 509260 294696 509312
rect 294748 509300 294754 509312
rect 297726 509300 297732 509312
rect 294748 509272 297732 509300
rect 294748 509260 294754 509272
rect 297726 509260 297732 509272
rect 297784 509260 297790 509312
rect 192478 506472 192484 506524
rect 192536 506512 192542 506524
rect 297726 506512 297732 506524
rect 192536 506484 297732 506512
rect 192536 506472 192542 506484
rect 297726 506472 297732 506484
rect 297784 506472 297790 506524
rect 153562 505220 153568 505232
rect 153396 505192 153568 505220
rect 153396 505096 153424 505192
rect 153562 505180 153568 505192
rect 153620 505180 153626 505232
rect 128630 505044 128636 505096
rect 128688 505084 128694 505096
rect 128814 505084 128820 505096
rect 128688 505056 128820 505084
rect 128688 505044 128694 505056
rect 128814 505044 128820 505056
rect 128872 505044 128878 505096
rect 153378 505044 153384 505096
rect 153436 505044 153442 505096
rect 96522 500896 96528 500948
rect 96580 500936 96586 500948
rect 379514 500936 379520 500948
rect 96580 500908 379520 500936
rect 96580 500896 96586 500908
rect 379514 500896 379520 500908
rect 379572 500896 379578 500948
rect 103514 500828 103520 500880
rect 103572 500868 103578 500880
rect 104802 500868 104808 500880
rect 103572 500840 104808 500868
rect 103572 500828 103578 500840
rect 104802 500828 104808 500840
rect 104860 500868 104866 500880
rect 379422 500868 379428 500880
rect 104860 500840 379428 500868
rect 104860 500828 104866 500840
rect 379422 500828 379428 500840
rect 379480 500828 379486 500880
rect 69842 500216 69848 500268
rect 69900 500256 69906 500268
rect 95234 500256 95240 500268
rect 69900 500228 95240 500256
rect 69900 500216 69906 500228
rect 95234 500216 95240 500228
rect 95292 500256 95298 500268
rect 96522 500256 96528 500268
rect 95292 500228 96528 500256
rect 95292 500216 95298 500228
rect 96522 500216 96528 500228
rect 96580 500216 96586 500268
rect 118050 499468 118056 499520
rect 118108 499508 118114 499520
rect 302878 499508 302884 499520
rect 118108 499480 302884 499508
rect 118108 499468 118114 499480
rect 302878 499468 302884 499480
rect 302936 499468 302942 499520
rect 300486 499128 300492 499180
rect 300544 499168 300550 499180
rect 311894 499168 311900 499180
rect 300544 499140 311900 499168
rect 300544 499128 300550 499140
rect 311894 499128 311900 499140
rect 311952 499128 311958 499180
rect 298370 499060 298376 499112
rect 298428 499100 298434 499112
rect 310606 499100 310612 499112
rect 298428 499072 310612 499100
rect 298428 499060 298434 499072
rect 310606 499060 310612 499072
rect 310664 499060 310670 499112
rect 324222 499060 324228 499112
rect 324280 499100 324286 499112
rect 378410 499100 378416 499112
rect 324280 499072 378416 499100
rect 324280 499060 324286 499072
rect 378410 499060 378416 499072
rect 378468 499060 378474 499112
rect 298278 498992 298284 499044
rect 298336 499032 298342 499044
rect 314746 499032 314752 499044
rect 298336 499004 314752 499032
rect 298336 498992 298342 499004
rect 314746 498992 314752 499004
rect 314804 498992 314810 499044
rect 321462 498992 321468 499044
rect 321520 499032 321526 499044
rect 378318 499032 378324 499044
rect 321520 499004 378324 499032
rect 321520 498992 321526 499004
rect 378318 498992 378324 499004
rect 378376 498992 378382 499044
rect 298554 498924 298560 498976
rect 298612 498964 298618 498976
rect 316034 498964 316040 498976
rect 298612 498936 316040 498964
rect 298612 498924 298618 498936
rect 316034 498924 316040 498936
rect 316092 498924 316098 498976
rect 317322 498924 317328 498976
rect 317380 498964 317386 498976
rect 378226 498964 378232 498976
rect 317380 498936 378232 498964
rect 317380 498924 317386 498936
rect 378226 498924 378232 498936
rect 378284 498924 378290 498976
rect 298462 498856 298468 498908
rect 298520 498896 298526 498908
rect 309134 498896 309140 498908
rect 298520 498868 309140 498896
rect 298520 498856 298526 498868
rect 309134 498856 309140 498868
rect 309192 498856 309198 498908
rect 310422 498856 310428 498908
rect 310480 498896 310486 498908
rect 378594 498896 378600 498908
rect 310480 498868 378600 498896
rect 310480 498856 310486 498868
rect 378594 498856 378600 498868
rect 378652 498856 378658 498908
rect 298646 498788 298652 498840
rect 298704 498828 298710 498840
rect 306466 498828 306472 498840
rect 298704 498800 306472 498828
rect 298704 498788 298710 498800
rect 306466 498788 306472 498800
rect 306524 498788 306530 498840
rect 309042 498788 309048 498840
rect 309100 498828 309106 498840
rect 378502 498828 378508 498840
rect 309100 498800 378508 498828
rect 309100 498788 309106 498800
rect 378502 498788 378508 498800
rect 378560 498788 378566 498840
rect 300394 498584 300400 498636
rect 300452 498624 300458 498636
rect 302234 498624 302240 498636
rect 300452 498596 302240 498624
rect 300452 498584 300458 498596
rect 302234 498584 302240 498596
rect 302292 498584 302298 498636
rect 132126 498176 132132 498228
rect 132184 498216 132190 498228
rect 580166 498216 580172 498228
rect 132184 498188 580172 498216
rect 132184 498176 132190 498188
rect 580166 498176 580172 498188
rect 580224 498176 580230 498228
rect 129090 498108 129096 498160
rect 129148 498148 129154 498160
rect 364242 498148 364248 498160
rect 129148 498120 364248 498148
rect 129148 498108 129154 498120
rect 364242 498108 364248 498120
rect 364300 498108 364306 498160
rect 116026 498040 116032 498092
rect 116084 498080 116090 498092
rect 347314 498080 347320 498092
rect 116084 498052 347320 498080
rect 116084 498040 116090 498052
rect 347314 498040 347320 498052
rect 347372 498040 347378 498092
rect 120718 497972 120724 498024
rect 120776 498012 120782 498024
rect 121362 498012 121368 498024
rect 120776 497984 121368 498012
rect 120776 497972 120782 497984
rect 121362 497972 121368 497984
rect 121420 498012 121426 498024
rect 338850 498012 338856 498024
rect 121420 497984 338856 498012
rect 121420 497972 121426 497984
rect 338850 497972 338856 497984
rect 338908 497972 338914 498024
rect 126330 497904 126336 497956
rect 126388 497944 126394 497956
rect 334434 497944 334440 497956
rect 126388 497916 334440 497944
rect 126388 497904 126394 497916
rect 334434 497904 334440 497916
rect 334492 497904 334498 497956
rect 337470 497904 337476 497956
rect 337528 497944 337534 497956
rect 370682 497944 370688 497956
rect 337528 497916 370688 497944
rect 337528 497904 337534 497916
rect 370682 497904 370688 497916
rect 370740 497904 370746 497956
rect 152458 497836 152464 497888
rect 152516 497876 152522 497888
rect 153102 497876 153108 497888
rect 152516 497848 153108 497876
rect 152516 497836 152522 497848
rect 153102 497836 153108 497848
rect 153160 497876 153166 497888
rect 319714 497876 319720 497888
rect 153160 497848 319720 497876
rect 153160 497836 153166 497848
rect 319714 497836 319720 497848
rect 319772 497836 319778 497888
rect 320082 497836 320088 497888
rect 320140 497876 320146 497888
rect 357986 497876 357992 497888
rect 320140 497848 357992 497876
rect 320140 497836 320146 497848
rect 357986 497836 357992 497848
rect 358044 497836 358050 497888
rect 289722 497768 289728 497820
rect 289780 497808 289786 497820
rect 366450 497808 366456 497820
rect 289780 497780 366456 497808
rect 289780 497768 289786 497780
rect 366450 497768 366456 497780
rect 366508 497768 366514 497820
rect 284294 497700 284300 497752
rect 284352 497740 284358 497752
rect 368474 497740 368480 497752
rect 284352 497712 368480 497740
rect 284352 497700 284358 497712
rect 368474 497700 368480 497712
rect 368532 497700 368538 497752
rect 111702 497632 111708 497684
rect 111760 497672 111766 497684
rect 115290 497672 115296 497684
rect 111760 497644 115296 497672
rect 111760 497632 111766 497644
rect 115290 497632 115296 497644
rect 115348 497632 115354 497684
rect 291010 497632 291016 497684
rect 291068 497672 291074 497684
rect 377122 497672 377128 497684
rect 291068 497644 377128 497672
rect 291068 497632 291074 497644
rect 377122 497632 377128 497644
rect 377180 497632 377186 497684
rect 108942 497564 108948 497616
rect 109000 497604 109006 497616
rect 116026 497604 116032 497616
rect 109000 497576 116032 497604
rect 109000 497564 109006 497576
rect 116026 497564 116032 497576
rect 116084 497564 116090 497616
rect 284202 497564 284208 497616
rect 284260 497604 284266 497616
rect 374914 497604 374920 497616
rect 284260 497576 374920 497604
rect 284260 497564 284266 497576
rect 374914 497564 374920 497576
rect 374972 497564 374978 497616
rect 83918 497496 83924 497548
rect 83976 497536 83982 497548
rect 127066 497536 127072 497548
rect 83976 497508 127072 497536
rect 83976 497496 83982 497508
rect 127066 497496 127072 497508
rect 127124 497536 127130 497548
rect 360010 497536 360016 497548
rect 127124 497508 360016 497536
rect 127124 497496 127130 497508
rect 360010 497496 360016 497508
rect 360068 497496 360074 497548
rect 111794 497428 111800 497480
rect 111852 497468 111858 497480
rect 125962 497468 125968 497480
rect 111852 497440 125968 497468
rect 111852 497428 111858 497440
rect 125962 497428 125968 497440
rect 126020 497468 126026 497480
rect 372706 497468 372712 497480
rect 126020 497440 372712 497468
rect 126020 497428 126026 497440
rect 372706 497428 372712 497440
rect 372764 497428 372770 497480
rect 285582 497360 285588 497412
rect 285640 497400 285646 497412
rect 345106 497400 345112 497412
rect 285640 497372 345112 497400
rect 285640 497360 285646 497372
rect 345106 497360 345112 497372
rect 345164 497360 345170 497412
rect 292482 497292 292488 497344
rect 292540 497332 292546 497344
rect 351546 497332 351552 497344
rect 292540 497304 351552 497332
rect 292540 497292 292546 497304
rect 351546 497292 351552 497304
rect 351604 497292 351610 497344
rect 301498 497224 301504 497276
rect 301556 497264 301562 497276
rect 353570 497264 353576 497276
rect 301556 497236 353576 497264
rect 301556 497224 301562 497236
rect 353570 497224 353576 497236
rect 353628 497224 353634 497276
rect 295242 497156 295248 497208
rect 295300 497196 295306 497208
rect 340874 497196 340880 497208
rect 295300 497168 340880 497196
rect 295300 497156 295306 497168
rect 340874 497156 340880 497168
rect 340932 497156 340938 497208
rect 277302 497088 277308 497140
rect 277360 497128 277366 497140
rect 317506 497128 317512 497140
rect 277360 497100 317512 497128
rect 277360 497088 277366 497100
rect 317506 497088 317512 497100
rect 317564 497088 317570 497140
rect 319438 497088 319444 497140
rect 319496 497128 319502 497140
rect 349338 497128 349344 497140
rect 319496 497100 349344 497128
rect 319496 497088 319502 497100
rect 349338 497088 349344 497100
rect 349396 497088 349402 497140
rect 288342 497020 288348 497072
rect 288400 497060 288406 497072
rect 321738 497060 321744 497072
rect 288400 497032 321744 497060
rect 288400 497020 288406 497032
rect 321738 497020 321744 497032
rect 321796 497020 321802 497072
rect 334618 497020 334624 497072
rect 334676 497060 334682 497072
rect 362218 497060 362224 497072
rect 334676 497032 362224 497060
rect 334676 497020 334682 497032
rect 362218 497020 362224 497032
rect 362276 497020 362282 497072
rect 279510 496952 279516 497004
rect 279568 496992 279574 497004
rect 311066 496992 311072 497004
rect 279568 496964 311072 496992
rect 279568 496952 279574 496964
rect 311066 496952 311072 496964
rect 311124 496952 311130 497004
rect 333238 496952 333244 497004
rect 333296 496992 333302 497004
rect 355778 496992 355784 497004
rect 333296 496964 355784 496992
rect 333296 496952 333302 496964
rect 355778 496952 355784 496964
rect 355836 496952 355842 497004
rect 304258 496884 304264 496936
rect 304316 496924 304322 496936
rect 332410 496924 332416 496936
rect 304316 496896 332416 496924
rect 304316 496884 304322 496896
rect 332410 496884 332416 496896
rect 332468 496884 332474 496936
rect 126330 496816 126336 496868
rect 126388 496856 126394 496868
rect 126882 496856 126888 496868
rect 126388 496828 126888 496856
rect 126388 496816 126394 496828
rect 126882 496816 126888 496828
rect 126940 496816 126946 496868
rect 285030 496816 285036 496868
rect 285088 496856 285094 496868
rect 306834 496856 306840 496868
rect 285088 496828 306840 496856
rect 285088 496816 285094 496828
rect 306834 496816 306840 496828
rect 306892 496816 306898 496868
rect 308950 496816 308956 496868
rect 309008 496856 309014 496868
rect 316678 496856 316684 496868
rect 309008 496828 316684 496856
rect 309008 496816 309014 496828
rect 316678 496816 316684 496828
rect 316736 496816 316742 496868
rect 322198 496816 322204 496868
rect 322256 496856 322262 496868
rect 323946 496856 323952 496868
rect 322256 496828 323952 496856
rect 322256 496816 322262 496828
rect 323946 496816 323952 496828
rect 324004 496816 324010 496868
rect 330478 496816 330484 496868
rect 330536 496856 330542 496868
rect 336642 496856 336648 496868
rect 330536 496828 336648 496856
rect 330536 496816 330542 496828
rect 336642 496816 336648 496828
rect 336700 496816 336706 496868
rect 337378 496816 337384 496868
rect 337436 496856 337442 496868
rect 343082 496856 343088 496868
rect 337436 496828 343088 496856
rect 337436 496816 337442 496828
rect 343082 496816 343088 496828
rect 343140 496816 343146 496868
rect 3326 495456 3332 495508
rect 3384 495496 3390 495508
rect 31018 495496 31024 495508
rect 3384 495468 31024 495496
rect 3384 495456 3390 495468
rect 31018 495456 31024 495468
rect 31076 495456 31082 495508
rect 153378 495388 153384 495440
rect 153436 495428 153442 495440
rect 153562 495428 153568 495440
rect 153436 495400 153568 495428
rect 153436 495388 153442 495400
rect 153562 495388 153568 495400
rect 153620 495388 153626 495440
rect 153286 492600 153292 492652
rect 153344 492640 153350 492652
rect 153562 492640 153568 492652
rect 153344 492612 153568 492640
rect 153344 492600 153350 492612
rect 153562 492600 153568 492612
rect 153620 492600 153626 492652
rect 128630 491240 128636 491292
rect 128688 491280 128694 491292
rect 128722 491280 128728 491292
rect 128688 491252 128728 491280
rect 128688 491240 128694 491252
rect 128722 491240 128728 491252
rect 128780 491240 128786 491292
rect 284018 491280 284024 491292
rect 283979 491252 284024 491280
rect 284018 491240 284024 491252
rect 284076 491240 284082 491292
rect 299750 485800 299756 485852
rect 299808 485840 299814 485852
rect 300578 485840 300584 485852
rect 299808 485812 300584 485840
rect 299808 485800 299814 485812
rect 300578 485800 300584 485812
rect 300636 485800 300642 485852
rect 438210 485800 438216 485852
rect 438268 485840 438274 485852
rect 580166 485840 580172 485852
rect 438268 485812 580172 485840
rect 438268 485800 438274 485812
rect 580166 485800 580172 485812
rect 580224 485800 580230 485852
rect 284021 485775 284079 485781
rect 284021 485741 284033 485775
rect 284067 485772 284079 485775
rect 284110 485772 284116 485784
rect 284067 485744 284116 485772
rect 284067 485741 284079 485744
rect 284021 485735 284079 485741
rect 284110 485732 284116 485744
rect 284168 485732 284174 485784
rect 125962 481584 125968 481636
rect 126020 481624 126026 481636
rect 126054 481624 126060 481636
rect 126020 481596 126060 481624
rect 126020 481584 126026 481596
rect 126054 481584 126060 481596
rect 126112 481584 126118 481636
rect 284021 481627 284079 481633
rect 284021 481593 284033 481627
rect 284067 481624 284079 481627
rect 284110 481624 284116 481636
rect 284067 481596 284116 481624
rect 284067 481593 284079 481596
rect 284021 481587 284079 481593
rect 284110 481584 284116 481596
rect 284168 481584 284174 481636
rect 4062 480632 4068 480684
rect 4120 480672 4126 480684
rect 4982 480672 4988 480684
rect 4120 480644 4988 480672
rect 4120 480632 4126 480644
rect 4982 480632 4988 480644
rect 5040 480632 5046 480684
rect 153286 476076 153292 476128
rect 153344 476116 153350 476128
rect 153470 476116 153476 476128
rect 153344 476088 153476 476116
rect 153344 476076 153350 476088
rect 153470 476076 153476 476088
rect 153528 476076 153534 476128
rect 299566 476076 299572 476128
rect 299624 476116 299630 476128
rect 299750 476116 299756 476128
rect 299624 476088 299756 476116
rect 299624 476076 299630 476088
rect 299750 476076 299756 476088
rect 299808 476076 299814 476128
rect 153378 473328 153384 473340
rect 153339 473300 153384 473328
rect 153378 473288 153384 473300
rect 153436 473288 153442 473340
rect 299658 473328 299664 473340
rect 299619 473300 299664 473328
rect 299658 473288 299664 473300
rect 299716 473288 299722 473340
rect 153378 466392 153384 466404
rect 153339 466364 153384 466392
rect 153378 466352 153384 466364
rect 153436 466352 153442 466404
rect 299658 466392 299664 466404
rect 299619 466364 299664 466392
rect 299658 466352 299664 466364
rect 299716 466352 299722 466404
rect 284021 463811 284079 463817
rect 284021 463777 284033 463811
rect 284067 463808 284079 463811
rect 284110 463808 284116 463820
rect 284067 463780 284116 463808
rect 284067 463777 284079 463780
rect 284021 463771 284079 463777
rect 284110 463768 284116 463780
rect 284168 463768 284174 463820
rect 283834 463632 283840 463684
rect 283892 463672 283898 463684
rect 284110 463672 284116 463684
rect 283892 463644 284116 463672
rect 283892 463632 283898 463644
rect 284110 463632 284116 463644
rect 284168 463632 284174 463684
rect 133138 462340 133144 462392
rect 133196 462380 133202 462392
rect 579798 462380 579804 462392
rect 133196 462352 579804 462380
rect 133196 462340 133202 462352
rect 579798 462340 579804 462352
rect 579856 462340 579862 462392
rect 125962 456832 125968 456884
rect 126020 456832 126026 456884
rect 125980 456748 126008 456832
rect 299566 456764 299572 456816
rect 299624 456804 299630 456816
rect 299750 456804 299756 456816
rect 299624 456776 299756 456804
rect 299624 456764 299630 456776
rect 299750 456764 299756 456776
rect 299808 456764 299814 456816
rect 125962 456696 125968 456748
rect 126020 456696 126026 456748
rect 125962 453976 125968 454028
rect 126020 454016 126026 454028
rect 126054 454016 126060 454028
rect 126020 453988 126060 454016
rect 126020 453976 126026 453988
rect 126054 453976 126060 453988
rect 126112 453976 126118 454028
rect 284018 454016 284024 454028
rect 283979 453988 284024 454016
rect 284018 453976 284024 453988
rect 284076 453976 284082 454028
rect 299658 454016 299664 454028
rect 299619 453988 299664 454016
rect 299658 453976 299664 453988
rect 299716 453976 299722 454028
rect 126054 452588 126060 452600
rect 126015 452560 126060 452588
rect 126054 452548 126060 452560
rect 126112 452548 126118 452600
rect 3050 451324 3056 451376
rect 3108 451364 3114 451376
rect 267274 451364 267280 451376
rect 3108 451336 267280 451364
rect 3108 451324 3114 451336
rect 267274 451324 267280 451336
rect 267332 451324 267338 451376
rect 133230 451256 133236 451308
rect 133288 451296 133294 451308
rect 580166 451296 580172 451308
rect 133288 451268 580172 451296
rect 133288 451256 133294 451268
rect 580166 451256 580172 451268
rect 580224 451256 580230 451308
rect 299658 447080 299664 447092
rect 299619 447052 299664 447080
rect 299658 447040 299664 447052
rect 299716 447040 299722 447092
rect 284021 444499 284079 444505
rect 284021 444465 284033 444499
rect 284067 444496 284079 444499
rect 284110 444496 284116 444508
rect 284067 444468 284116 444496
rect 284067 444465 284079 444468
rect 284021 444459 284079 444465
rect 284110 444456 284116 444468
rect 284168 444456 284174 444508
rect 153378 444360 153384 444372
rect 153339 444332 153384 444360
rect 153378 444320 153384 444332
rect 153436 444320 153442 444372
rect 283834 444320 283840 444372
rect 283892 444360 283898 444372
rect 284110 444360 284116 444372
rect 283892 444332 284116 444360
rect 283892 444320 283898 444332
rect 284110 444320 284116 444332
rect 284168 444320 284174 444372
rect 126054 443816 126060 443828
rect 126015 443788 126060 443816
rect 126054 443776 126060 443788
rect 126112 443776 126118 443828
rect 436738 438880 436744 438932
rect 436796 438920 436802 438932
rect 580166 438920 580172 438932
rect 436796 438892 580172 438920
rect 436796 438880 436802 438892
rect 580166 438880 580172 438892
rect 580224 438880 580230 438932
rect 299566 437452 299572 437504
rect 299624 437492 299630 437504
rect 299750 437492 299756 437504
rect 299624 437464 299756 437492
rect 299624 437452 299630 437464
rect 299750 437452 299756 437464
rect 299808 437452 299814 437504
rect 153378 437424 153384 437436
rect 153339 437396 153384 437424
rect 153378 437384 153384 437396
rect 153436 437384 153442 437436
rect 125873 434707 125931 434713
rect 125873 434673 125885 434707
rect 125919 434704 125931 434707
rect 125962 434704 125968 434716
rect 125919 434676 125968 434704
rect 125919 434673 125931 434676
rect 125873 434667 125931 434673
rect 125962 434664 125968 434676
rect 126020 434664 126026 434716
rect 284018 434704 284024 434716
rect 283979 434676 284024 434704
rect 284018 434664 284024 434676
rect 284076 434664 284082 434716
rect 299658 434704 299664 434716
rect 299619 434676 299664 434704
rect 299658 434664 299664 434676
rect 299716 434664 299722 434716
rect 125870 427768 125876 427780
rect 125831 427740 125876 427768
rect 125870 427728 125876 427740
rect 125928 427728 125934 427780
rect 299658 427768 299664 427780
rect 299619 427740 299664 427768
rect 299658 427728 299664 427740
rect 299716 427728 299722 427780
rect 284021 425187 284079 425193
rect 284021 425153 284033 425187
rect 284067 425184 284079 425187
rect 284110 425184 284116 425196
rect 284067 425156 284116 425184
rect 284067 425153 284079 425156
rect 284021 425147 284079 425153
rect 284110 425144 284116 425156
rect 284168 425144 284174 425196
rect 125870 425008 125876 425060
rect 125928 425048 125934 425060
rect 125962 425048 125968 425060
rect 125928 425020 125968 425048
rect 125928 425008 125934 425020
rect 125962 425008 125968 425020
rect 126020 425008 126026 425060
rect 283834 425008 283840 425060
rect 283892 425048 283898 425060
rect 284110 425048 284116 425060
rect 283892 425020 284116 425048
rect 283892 425008 283898 425020
rect 284110 425008 284116 425020
rect 284168 425008 284174 425060
rect 4062 423648 4068 423700
rect 4120 423688 4126 423700
rect 5074 423688 5080 423700
rect 4120 423660 5080 423688
rect 4120 423648 4126 423660
rect 5074 423648 5080 423660
rect 5132 423648 5138 423700
rect 153286 418248 153292 418260
rect 153212 418220 153292 418248
rect 153212 418124 153240 418220
rect 153286 418208 153292 418220
rect 153344 418208 153350 418260
rect 299566 418140 299572 418192
rect 299624 418180 299630 418192
rect 299750 418180 299756 418192
rect 299624 418152 299756 418180
rect 299624 418140 299630 418152
rect 299750 418140 299756 418152
rect 299808 418140 299814 418192
rect 153194 418072 153200 418124
rect 153252 418072 153258 418124
rect 133046 415420 133052 415472
rect 133104 415460 133110 415472
rect 579798 415460 579804 415472
rect 133104 415432 579804 415460
rect 133104 415420 133110 415432
rect 579798 415420 579804 415432
rect 579856 415420 579862 415472
rect 126057 415395 126115 415401
rect 126057 415361 126069 415395
rect 126103 415392 126115 415395
rect 126146 415392 126152 415404
rect 126103 415364 126152 415392
rect 126103 415361 126115 415364
rect 126057 415355 126115 415361
rect 126146 415352 126152 415364
rect 126204 415352 126210 415404
rect 128541 415395 128599 415401
rect 128541 415361 128553 415395
rect 128587 415392 128599 415395
rect 128630 415392 128636 415404
rect 128587 415364 128636 415392
rect 128587 415361 128599 415364
rect 128541 415355 128599 415361
rect 128630 415352 128636 415364
rect 128688 415352 128694 415404
rect 153194 415352 153200 415404
rect 153252 415392 153258 415404
rect 153470 415392 153476 415404
rect 153252 415364 153476 415392
rect 153252 415352 153258 415364
rect 153470 415352 153476 415364
rect 153528 415352 153534 415404
rect 284018 415392 284024 415404
rect 283979 415364 284024 415392
rect 284018 415352 284024 415364
rect 284076 415352 284082 415404
rect 299658 415392 299664 415404
rect 299619 415364 299664 415392
rect 299658 415352 299664 415364
rect 299716 415352 299722 415404
rect 251726 410796 251732 410848
rect 251784 410836 251790 410848
rect 266354 410836 266360 410848
rect 251784 410808 266360 410836
rect 251784 410796 251790 410808
rect 266354 410796 266360 410808
rect 266412 410796 266418 410848
rect 246022 410728 246028 410780
rect 246080 410768 246086 410780
rect 267826 410768 267832 410780
rect 246080 410740 267832 410768
rect 246080 410728 246086 410740
rect 267826 410728 267832 410740
rect 267884 410728 267890 410780
rect 228910 410660 228916 410712
rect 228968 410700 228974 410712
rect 266998 410700 267004 410712
rect 228968 410672 267004 410700
rect 228968 410660 228974 410672
rect 266998 410660 267004 410672
rect 267056 410660 267062 410712
rect 223390 410592 223396 410644
rect 223448 410632 223454 410644
rect 266722 410632 266728 410644
rect 223448 410604 266728 410632
rect 223448 410592 223454 410604
rect 266722 410592 266728 410604
rect 266780 410592 266786 410644
rect 211982 410524 211988 410576
rect 212040 410564 212046 410576
rect 267090 410564 267096 410576
rect 212040 410536 267096 410564
rect 212040 410524 212046 410536
rect 267090 410524 267096 410536
rect 267148 410524 267154 410576
rect 206278 410456 206284 410508
rect 206336 410496 206342 410508
rect 266446 410496 266452 410508
rect 206336 410468 266452 410496
rect 206336 410456 206342 410468
rect 266446 410456 266452 410468
rect 266504 410456 266510 410508
rect 248966 410388 248972 410440
rect 249024 410428 249030 410440
rect 267734 410428 267740 410440
rect 249024 410400 267740 410428
rect 249024 410388 249030 410400
rect 267734 410388 267740 410400
rect 267792 410388 267798 410440
rect 243262 410320 243268 410372
rect 243320 410360 243326 410372
rect 266538 410360 266544 410372
rect 243320 410332 266544 410360
rect 243320 410320 243326 410332
rect 266538 410320 266544 410332
rect 266596 410320 266602 410372
rect 240318 410252 240324 410304
rect 240376 410292 240382 410304
rect 266630 410292 266636 410304
rect 240376 410264 266636 410292
rect 240376 410252 240382 410264
rect 266630 410252 266636 410264
rect 266688 410252 266694 410304
rect 237558 410184 237564 410236
rect 237616 410224 237622 410236
rect 267366 410224 267372 410236
rect 237616 410196 267372 410224
rect 237616 410184 237622 410196
rect 267366 410184 267372 410196
rect 267424 410184 267430 410236
rect 196894 410116 196900 410168
rect 196952 410156 196958 410168
rect 200574 410156 200580 410168
rect 196952 410128 200580 410156
rect 196952 410116 196958 410128
rect 200574 410116 200580 410128
rect 200632 410116 200638 410168
rect 234614 410116 234620 410168
rect 234672 410156 234678 410168
rect 266814 410156 266820 410168
rect 234672 410128 266820 410156
rect 234672 410116 234678 410128
rect 266814 410116 266820 410128
rect 266872 410116 266878 410168
rect 199746 410048 199752 410100
rect 199804 410088 199810 410100
rect 217686 410088 217692 410100
rect 199804 410060 217692 410088
rect 199804 410048 199810 410060
rect 217686 410048 217692 410060
rect 217744 410048 217750 410100
rect 257430 410048 257436 410100
rect 257488 410088 257494 410100
rect 267458 410088 267464 410100
rect 257488 410060 267464 410088
rect 257488 410048 257494 410060
rect 267458 410048 267464 410060
rect 267516 410048 267522 410100
rect 199838 409980 199844 410032
rect 199896 410020 199902 410032
rect 220446 410020 220452 410032
rect 199896 409992 220452 410020
rect 199896 409980 199902 409992
rect 220446 409980 220452 409992
rect 220504 409980 220510 410032
rect 254670 409980 254676 410032
rect 254728 410020 254734 410032
rect 268838 410020 268844 410032
rect 254728 409992 268844 410020
rect 254728 409980 254734 409992
rect 268838 409980 268844 409992
rect 268896 409980 268902 410032
rect 199930 409912 199936 409964
rect 199988 409952 199994 409964
rect 214742 409952 214748 409964
rect 199988 409924 214748 409952
rect 199988 409912 199994 409924
rect 214742 409912 214748 409924
rect 214800 409912 214806 409964
rect 260374 409912 260380 409964
rect 260432 409952 260438 409964
rect 267550 409952 267556 409964
rect 260432 409924 267556 409952
rect 260432 409912 260438 409924
rect 267550 409912 267556 409924
rect 267608 409912 267614 409964
rect 200022 409844 200028 409896
rect 200080 409884 200086 409896
rect 209038 409884 209044 409896
rect 200080 409856 209044 409884
rect 200080 409844 200086 409856
rect 209038 409844 209044 409856
rect 209096 409844 209102 409896
rect 265894 409844 265900 409896
rect 265952 409884 265958 409896
rect 268930 409884 268936 409896
rect 265952 409856 268936 409884
rect 265952 409844 265958 409856
rect 268930 409844 268936 409856
rect 268988 409844 268994 409896
rect 199562 409640 199568 409692
rect 199620 409680 199626 409692
rect 202874 409680 202880 409692
rect 199620 409652 202880 409680
rect 199620 409640 199626 409652
rect 202874 409640 202880 409652
rect 202932 409640 202938 409692
rect 199654 409572 199660 409624
rect 199712 409612 199718 409624
rect 205634 409612 205640 409624
rect 199712 409584 205640 409612
rect 199712 409572 199718 409584
rect 205634 409572 205640 409584
rect 205692 409572 205698 409624
rect 196802 409504 196808 409556
rect 196860 409544 196866 409556
rect 209774 409544 209780 409556
rect 196860 409516 209780 409544
rect 196860 409504 196866 409516
rect 209774 409504 209780 409516
rect 209832 409504 209838 409556
rect 195606 409436 195612 409488
rect 195664 409476 195670 409488
rect 212534 409476 212540 409488
rect 195664 409448 212540 409476
rect 195664 409436 195670 409448
rect 212534 409436 212540 409448
rect 212592 409436 212598 409488
rect 195790 409368 195796 409420
rect 195848 409408 195854 409420
rect 215294 409408 215300 409420
rect 195848 409380 215300 409408
rect 195848 409368 195854 409380
rect 215294 409368 215300 409380
rect 215352 409368 215358 409420
rect 196710 409300 196716 409352
rect 196768 409340 196774 409352
rect 222746 409340 222752 409352
rect 196768 409312 222752 409340
rect 196768 409300 196774 409312
rect 222746 409300 222752 409312
rect 222804 409300 222810 409352
rect 196618 409232 196624 409284
rect 196676 409272 196682 409284
rect 222838 409272 222844 409284
rect 196676 409244 222844 409272
rect 196676 409232 196682 409244
rect 222838 409232 222844 409244
rect 222896 409232 222902 409284
rect 195698 409164 195704 409216
rect 195756 409204 195762 409216
rect 222194 409204 222200 409216
rect 195756 409176 222200 409204
rect 195756 409164 195762 409176
rect 222194 409164 222200 409176
rect 222252 409164 222258 409216
rect 195514 409096 195520 409148
rect 195572 409136 195578 409148
rect 222286 409136 222292 409148
rect 195572 409108 222292 409136
rect 195572 409096 195578 409108
rect 222286 409096 222292 409108
rect 222344 409096 222350 409148
rect 188338 407804 188344 407856
rect 188396 407844 188402 407856
rect 377398 407844 377404 407856
rect 188396 407816 377404 407844
rect 188396 407804 188402 407816
rect 377398 407804 377404 407816
rect 377456 407804 377462 407856
rect 70210 407736 70216 407788
rect 70268 407776 70274 407788
rect 104802 407776 104808 407788
rect 70268 407748 104808 407776
rect 70268 407736 70274 407748
rect 104802 407736 104808 407748
rect 104860 407776 104866 407788
rect 393314 407776 393320 407788
rect 104860 407748 393320 407776
rect 104860 407736 104866 407748
rect 393314 407736 393320 407748
rect 393372 407736 393378 407788
rect 197998 407192 198004 407244
rect 198056 407232 198062 407244
rect 386414 407232 386420 407244
rect 198056 407204 386420 407232
rect 198056 407192 198062 407204
rect 386414 407192 386420 407204
rect 386472 407192 386478 407244
rect 130378 407124 130384 407176
rect 130436 407164 130442 407176
rect 358078 407164 358084 407176
rect 130436 407136 358084 407164
rect 130436 407124 130442 407136
rect 358078 407124 358084 407136
rect 358136 407124 358142 407176
rect 197722 406580 197728 406632
rect 197780 406620 197786 406632
rect 295334 406620 295340 406632
rect 197780 406592 295340 406620
rect 197780 406580 197786 406592
rect 295334 406580 295340 406592
rect 295392 406580 295398 406632
rect 70302 406512 70308 406564
rect 70360 406552 70366 406564
rect 295978 406552 295984 406564
rect 70360 406524 295984 406552
rect 70360 406512 70366 406524
rect 295978 406512 295984 406524
rect 296036 406512 296042 406564
rect 153102 406444 153108 406496
rect 153160 406484 153166 406496
rect 393406 406484 393412 406496
rect 153160 406456 393412 406484
rect 153160 406444 153166 406456
rect 393406 406444 393412 406456
rect 393464 406444 393470 406496
rect 295978 406376 295984 406428
rect 296036 406416 296042 406428
rect 344278 406416 344284 406428
rect 296036 406388 344284 406416
rect 296036 406376 296042 406388
rect 344278 406376 344284 406388
rect 344336 406376 344342 406428
rect 152458 405968 152464 406020
rect 152516 406008 152522 406020
rect 153102 406008 153108 406020
rect 152516 405980 153108 406008
rect 152516 405968 152522 405980
rect 153102 405968 153108 405980
rect 153160 405968 153166 406020
rect 126054 405736 126060 405748
rect 126015 405708 126060 405736
rect 126054 405696 126060 405708
rect 126112 405696 126118 405748
rect 128538 405736 128544 405748
rect 128499 405708 128544 405736
rect 128538 405696 128544 405708
rect 128596 405696 128602 405748
rect 284018 405736 284024 405748
rect 283979 405708 284024 405736
rect 284018 405696 284024 405708
rect 284076 405696 284082 405748
rect 295334 405696 295340 405748
rect 295392 405736 295398 405748
rect 296070 405736 296076 405748
rect 295392 405708 296076 405736
rect 295392 405696 295398 405708
rect 296070 405696 296076 405708
rect 296128 405696 296134 405748
rect 299661 405739 299719 405745
rect 299661 405705 299673 405739
rect 299707 405736 299719 405739
rect 299750 405736 299756 405748
rect 299707 405708 299756 405736
rect 299707 405705 299719 405708
rect 299661 405699 299719 405705
rect 299750 405696 299756 405708
rect 299808 405696 299814 405748
rect 128538 405600 128544 405612
rect 128499 405572 128544 405600
rect 128538 405560 128544 405572
rect 128596 405560 128602 405612
rect 386414 402908 386420 402960
rect 386472 402948 386478 402960
rect 387242 402948 387248 402960
rect 386472 402920 387248 402948
rect 386472 402908 386478 402920
rect 387242 402908 387248 402920
rect 387300 402908 387306 402960
rect 120902 399304 120908 399356
rect 120960 399344 120966 399356
rect 121362 399344 121368 399356
rect 120960 399316 121368 399344
rect 120960 399304 120966 399316
rect 121362 399304 121368 399316
rect 121420 399344 121426 399356
rect 125686 399344 125692 399356
rect 121420 399316 125692 399344
rect 121420 399304 121426 399316
rect 125686 399304 125692 399316
rect 125744 399304 125750 399356
rect 153378 398936 153384 398948
rect 153339 398908 153384 398936
rect 153378 398896 153384 398908
rect 153436 398896 153442 398948
rect 71682 398828 71688 398880
rect 71740 398868 71746 398880
rect 85482 398868 85488 398880
rect 71740 398840 85488 398868
rect 71740 398828 71746 398840
rect 85482 398828 85488 398840
rect 85540 398828 85546 398880
rect 85482 398692 85488 398744
rect 85540 398732 85546 398744
rect 90266 398732 90272 398744
rect 85540 398704 90272 398732
rect 85540 398692 85546 398704
rect 90266 398692 90272 398704
rect 90324 398692 90330 398744
rect 128541 398735 128599 398741
rect 128541 398701 128553 398735
rect 128587 398732 128599 398735
rect 128630 398732 128636 398744
rect 128587 398704 128636 398732
rect 128587 398701 128599 398704
rect 128541 398695 128599 398701
rect 128630 398692 128636 398704
rect 128688 398692 128694 398744
rect 379514 398624 379520 398676
rect 379572 398664 379578 398676
rect 380618 398664 380624 398676
rect 379572 398636 380624 398664
rect 379572 398624 379578 398636
rect 380618 398624 380624 398636
rect 380676 398624 380682 398676
rect 380434 398488 380440 398540
rect 380492 398528 380498 398540
rect 380618 398528 380624 398540
rect 380492 398500 380624 398528
rect 380492 398488 380498 398500
rect 380618 398488 380624 398500
rect 380676 398488 380682 398540
rect 380158 398352 380164 398404
rect 380216 398392 380222 398404
rect 380434 398392 380440 398404
rect 380216 398364 380440 398392
rect 380216 398352 380222 398364
rect 380434 398352 380440 398364
rect 380492 398352 380498 398404
rect 129458 398148 129464 398200
rect 129516 398188 129522 398200
rect 152458 398188 152464 398200
rect 129516 398160 152464 398188
rect 129516 398148 129522 398160
rect 152458 398148 152464 398160
rect 152516 398148 152522 398200
rect 75822 398080 75828 398132
rect 75880 398120 75886 398132
rect 115934 398120 115940 398132
rect 75880 398092 115940 398120
rect 75880 398080 75886 398092
rect 115934 398080 115940 398092
rect 115992 398120 115998 398132
rect 127250 398120 127256 398132
rect 115992 398092 127256 398120
rect 115992 398080 115998 398092
rect 127250 398080 127256 398092
rect 127308 398080 127314 398132
rect 134150 398080 134156 398132
rect 134208 398120 134214 398132
rect 191098 398120 191104 398132
rect 134208 398092 191104 398120
rect 134208 398080 134214 398092
rect 191098 398080 191104 398092
rect 191156 398080 191162 398132
rect 80790 397876 80796 397928
rect 80848 397916 80854 397928
rect 124858 397916 124864 397928
rect 80848 397888 124864 397916
rect 80848 397876 80854 397888
rect 124858 397876 124864 397888
rect 124916 397876 124922 397928
rect 100662 397808 100668 397860
rect 100720 397848 100726 397860
rect 113174 397848 113180 397860
rect 100720 397820 113180 397848
rect 100720 397808 100726 397820
rect 113174 397808 113180 397820
rect 113232 397848 113238 397860
rect 114462 397848 114468 397860
rect 113232 397820 114468 397848
rect 113232 397808 113238 397820
rect 114462 397808 114468 397820
rect 114520 397808 114526 397860
rect 110966 397740 110972 397792
rect 111024 397780 111030 397792
rect 111702 397780 111708 397792
rect 111024 397752 111708 397780
rect 111024 397740 111030 397752
rect 111702 397740 111708 397752
rect 111760 397780 111766 397792
rect 127158 397780 127164 397792
rect 111760 397752 127164 397780
rect 111760 397740 111766 397752
rect 127158 397740 127164 397752
rect 127216 397740 127222 397792
rect 105998 397672 106004 397724
rect 106056 397712 106062 397724
rect 127618 397712 127624 397724
rect 106056 397684 127624 397712
rect 106056 397672 106062 397684
rect 127618 397672 127624 397684
rect 127676 397672 127682 397724
rect 95878 397604 95884 397656
rect 95936 397644 95942 397656
rect 134150 397644 134156 397656
rect 95936 397616 134156 397644
rect 95936 397604 95942 397616
rect 134150 397604 134156 397616
rect 134208 397604 134214 397656
rect 85942 397536 85948 397588
rect 86000 397576 86006 397588
rect 129458 397576 129464 397588
rect 86000 397548 129464 397576
rect 86000 397536 86006 397548
rect 129458 397536 129464 397548
rect 129516 397536 129522 397588
rect 115842 397468 115848 397520
rect 115900 397508 115906 397520
rect 126330 397508 126336 397520
rect 115900 397480 126336 397508
rect 115900 397468 115906 397480
rect 126330 397468 126336 397480
rect 126388 397468 126394 397520
rect 124858 397400 124864 397452
rect 124916 397440 124922 397452
rect 126146 397440 126152 397452
rect 124916 397412 126152 397440
rect 124916 397400 124922 397412
rect 126146 397400 126152 397412
rect 126204 397400 126210 397452
rect 380066 397332 380072 397384
rect 380124 397372 380130 397384
rect 380250 397372 380256 397384
rect 380124 397344 380256 397372
rect 380124 397332 380130 397344
rect 380250 397332 380256 397344
rect 380308 397332 380314 397384
rect 69934 396788 69940 396840
rect 69992 396828 69998 396840
rect 117958 396828 117964 396840
rect 69992 396800 117964 396828
rect 69992 396788 69998 396800
rect 117958 396788 117964 396800
rect 118016 396828 118022 396840
rect 126514 396828 126520 396840
rect 118016 396800 126520 396828
rect 118016 396788 118022 396800
rect 126514 396788 126520 396800
rect 126572 396788 126578 396840
rect 114462 396720 114468 396772
rect 114520 396760 114526 396772
rect 128262 396760 128268 396772
rect 114520 396732 128268 396760
rect 114520 396720 114526 396732
rect 128262 396720 128268 396732
rect 128320 396760 128326 396772
rect 197998 396760 198004 396772
rect 128320 396732 198004 396760
rect 128320 396720 128326 396732
rect 197998 396720 198004 396732
rect 198056 396720 198062 396772
rect 153378 396080 153384 396092
rect 153339 396052 153384 396080
rect 153378 396040 153384 396052
rect 153436 396040 153442 396092
rect 133969 396015 134027 396021
rect 133969 395981 133981 396015
rect 134015 396012 134027 396015
rect 134150 396012 134156 396024
rect 134015 395984 134156 396012
rect 134015 395981 134027 395984
rect 133969 395975 134027 395981
rect 134150 395972 134156 395984
rect 134208 395972 134214 396024
rect 299566 396012 299572 396024
rect 299527 395984 299572 396012
rect 299566 395972 299572 395984
rect 299624 395972 299630 396024
rect 153289 395947 153347 395953
rect 153289 395913 153301 395947
rect 153335 395944 153347 395947
rect 153378 395944 153384 395956
rect 153335 395916 153384 395944
rect 153335 395913 153347 395916
rect 153289 395907 153347 395913
rect 153378 395904 153384 395916
rect 153436 395904 153442 395956
rect 84010 395836 84016 395888
rect 84068 395876 84074 395888
rect 84105 395879 84163 395885
rect 84105 395876 84117 395879
rect 84068 395848 84117 395876
rect 84068 395836 84074 395848
rect 84105 395845 84117 395848
rect 84151 395845 84163 395879
rect 84105 395839 84163 395845
rect 84013 395743 84071 395749
rect 84013 395709 84025 395743
rect 84059 395740 84071 395743
rect 84102 395740 84108 395752
rect 84059 395712 84108 395740
rect 84059 395709 84071 395712
rect 84013 395703 84071 395709
rect 84102 395700 84108 395712
rect 84160 395700 84166 395752
rect 70026 395632 70032 395684
rect 70084 395672 70090 395684
rect 108942 395672 108948 395684
rect 70084 395644 108948 395672
rect 70084 395632 70090 395644
rect 108942 395632 108948 395644
rect 109000 395672 109006 395684
rect 125870 395672 125876 395684
rect 109000 395644 125876 395672
rect 109000 395632 109006 395644
rect 125870 395632 125876 395644
rect 125928 395632 125934 395684
rect 84013 395607 84071 395613
rect 84013 395573 84025 395607
rect 84059 395573 84071 395607
rect 84013 395567 84071 395573
rect 84105 395607 84163 395613
rect 84105 395573 84117 395607
rect 84151 395604 84163 395607
rect 168650 395604 168656 395616
rect 84151 395576 168656 395604
rect 84151 395573 84163 395576
rect 84105 395567 84163 395573
rect 84028 395536 84056 395567
rect 168650 395564 168656 395576
rect 168708 395564 168714 395616
rect 179506 395536 179512 395548
rect 84028 395508 179512 395536
rect 179506 395496 179512 395508
rect 179564 395496 179570 395548
rect 349062 395428 349068 395480
rect 349120 395468 349126 395480
rect 361850 395468 361856 395480
rect 349120 395440 361856 395468
rect 349120 395428 349126 395440
rect 361850 395428 361856 395440
rect 361908 395428 361914 395480
rect 344278 395360 344284 395412
rect 344336 395400 344342 395412
rect 380250 395400 380256 395412
rect 344336 395372 380256 395400
rect 344336 395360 344342 395372
rect 380250 395360 380256 395372
rect 380308 395360 380314 395412
rect 296070 395292 296076 395344
rect 296128 395332 296134 395344
rect 364242 395332 364248 395344
rect 296128 395304 364248 395332
rect 296128 395292 296134 395304
rect 364242 395292 364248 395304
rect 364300 395292 364306 395344
rect 344922 395224 344928 395276
rect 344980 395264 344986 395276
rect 384850 395264 384856 395276
rect 344980 395236 384856 395264
rect 344980 395224 344986 395236
rect 384850 395224 384856 395236
rect 384908 395224 384914 395276
rect 355962 395156 355968 395208
rect 356020 395196 356026 395208
rect 389450 395196 389456 395208
rect 356020 395168 389456 395196
rect 356020 395156 356026 395168
rect 389450 395156 389456 395168
rect 389508 395156 389514 395208
rect 355870 395088 355876 395140
rect 355928 395128 355934 395140
rect 375650 395128 375656 395140
rect 355928 395100 375656 395128
rect 355928 395088 355934 395100
rect 375650 395088 375656 395100
rect 375708 395088 375714 395140
rect 353202 395020 353208 395072
rect 353260 395060 353266 395072
rect 378042 395060 378048 395072
rect 353260 395032 378048 395060
rect 353260 395020 353266 395032
rect 378042 395020 378048 395032
rect 378100 395020 378106 395072
rect 357345 394995 357403 395001
rect 357345 394961 357357 394995
rect 357391 394992 357403 394995
rect 382642 394992 382648 395004
rect 357391 394964 382648 394992
rect 357391 394961 357403 394964
rect 357345 394955 357403 394961
rect 382642 394952 382648 394964
rect 382700 394952 382706 395004
rect 347682 394884 347688 394936
rect 347740 394924 347746 394936
rect 373442 394924 373448 394936
rect 347740 394896 373448 394924
rect 347740 394884 347746 394896
rect 373442 394884 373448 394896
rect 373500 394884 373506 394936
rect 284018 394816 284024 394868
rect 284076 394816 284082 394868
rect 343542 394816 343548 394868
rect 343600 394856 343606 394868
rect 371050 394856 371056 394868
rect 343600 394828 371056 394856
rect 343600 394816 343606 394828
rect 371050 394816 371056 394828
rect 371108 394816 371114 394868
rect 284036 394732 284064 394816
rect 360010 394748 360016 394800
rect 360068 394788 360074 394800
rect 368842 394788 368848 394800
rect 360068 394760 368848 394788
rect 360068 394748 360074 394760
rect 368842 394748 368848 394760
rect 368900 394748 368906 394800
rect 284018 394680 284024 394732
rect 284076 394680 284082 394732
rect 360102 394680 360108 394732
rect 360160 394720 360166 394732
rect 366450 394720 366456 394732
rect 360160 394692 366456 394720
rect 360160 394680 360166 394692
rect 366450 394680 366456 394692
rect 366508 394680 366514 394732
rect 125778 394340 125784 394392
rect 125836 394380 125842 394392
rect 126146 394380 126152 394392
rect 125836 394352 126152 394380
rect 125836 394340 125842 394352
rect 126146 394340 126152 394352
rect 126204 394340 126210 394392
rect 315942 394068 315948 394120
rect 316000 394108 316006 394120
rect 380618 394108 380624 394120
rect 316000 394080 380624 394108
rect 316000 394068 316006 394080
rect 380618 394068 380624 394080
rect 380676 394068 380682 394120
rect 307662 394000 307668 394052
rect 307720 394040 307726 394052
rect 379422 394040 379428 394052
rect 307720 394012 379428 394040
rect 307720 394000 307726 394012
rect 379422 394000 379428 394012
rect 379480 394000 379486 394052
rect 271782 393932 271788 393984
rect 271840 393972 271846 393984
rect 380434 393972 380440 393984
rect 271840 393944 380440 393972
rect 271840 393932 271846 393944
rect 380434 393932 380440 393944
rect 380492 393932 380498 393984
rect 379422 393456 379428 393508
rect 379480 393496 379486 393508
rect 379698 393496 379704 393508
rect 379480 393468 379704 393496
rect 379480 393456 379486 393468
rect 379698 393456 379704 393468
rect 379756 393456 379762 393508
rect 380158 393388 380164 393440
rect 380216 393388 380222 393440
rect 379698 393320 379704 393372
rect 379756 393360 379762 393372
rect 380176 393360 380204 393388
rect 379756 393332 380204 393360
rect 379756 393320 379762 393332
rect 284018 393292 284024 393304
rect 283979 393264 284024 393292
rect 284018 393252 284024 393264
rect 284076 393252 284082 393304
rect 302142 393252 302148 393304
rect 302200 393292 302206 393304
rect 380342 393292 380348 393304
rect 302200 393264 380348 393292
rect 302200 393252 302206 393264
rect 380342 393252 380348 393264
rect 380400 393252 380406 393304
rect 300762 393184 300768 393236
rect 300820 393224 300826 393236
rect 379790 393224 379796 393236
rect 300820 393196 379796 393224
rect 300820 393184 300826 393196
rect 379790 393184 379796 393196
rect 379848 393184 379854 393236
rect 298646 393116 298652 393168
rect 298704 393156 298710 393168
rect 380526 393156 380532 393168
rect 298704 393128 380532 393156
rect 298704 393116 298710 393128
rect 380526 393116 380532 393128
rect 380584 393116 380590 393168
rect 297453 393091 297511 393097
rect 297453 393057 297465 393091
rect 297499 393088 297511 393091
rect 380066 393088 380072 393100
rect 297499 393060 380072 393088
rect 297499 393057 297511 393060
rect 297453 393051 297511 393057
rect 380066 393048 380072 393060
rect 380124 393048 380130 393100
rect 295150 392980 295156 393032
rect 295208 393020 295214 393032
rect 379514 393020 379520 393032
rect 295208 392992 379520 393020
rect 295208 392980 295214 392992
rect 379514 392980 379520 392992
rect 379572 392980 379578 393032
rect 292390 392912 292396 392964
rect 292448 392952 292454 392964
rect 377490 392952 377496 392964
rect 292448 392924 377496 392952
rect 292448 392912 292454 392924
rect 377490 392912 377496 392924
rect 377548 392912 377554 392964
rect 292298 392844 292304 392896
rect 292356 392884 292362 392896
rect 375929 392887 375987 392893
rect 375929 392884 375941 392887
rect 292356 392856 375941 392884
rect 292356 392844 292362 392856
rect 375929 392853 375941 392856
rect 375975 392853 375987 392887
rect 375929 392847 375987 392853
rect 376021 392887 376079 392893
rect 376021 392853 376033 392887
rect 376067 392884 376079 392887
rect 378134 392884 378140 392896
rect 376067 392856 378140 392884
rect 376067 392853 376079 392856
rect 376021 392847 376079 392853
rect 378134 392844 378140 392856
rect 378192 392844 378198 392896
rect 379422 392884 379428 392896
rect 379383 392856 379428 392884
rect 379422 392844 379428 392856
rect 379480 392844 379486 392896
rect 379606 392884 379612 392896
rect 379567 392856 379612 392884
rect 379606 392844 379612 392856
rect 379664 392844 379670 392896
rect 286870 392776 286876 392828
rect 286928 392816 286934 392828
rect 377030 392816 377036 392828
rect 286928 392788 377036 392816
rect 286928 392776 286934 392788
rect 377030 392776 377036 392788
rect 377088 392776 377094 392828
rect 377214 392816 377220 392828
rect 377175 392788 377220 392816
rect 377214 392776 377220 392788
rect 377272 392776 377278 392828
rect 379698 392816 379704 392828
rect 379659 392788 379704 392816
rect 379698 392776 379704 392788
rect 379756 392776 379762 392828
rect 379882 392776 379888 392828
rect 379940 392816 379946 392828
rect 379940 392788 380112 392816
rect 379940 392776 379946 392788
rect 288250 392708 288256 392760
rect 288308 392748 288314 392760
rect 375837 392751 375895 392757
rect 375837 392748 375849 392751
rect 288308 392720 375849 392748
rect 288308 392708 288314 392720
rect 375837 392717 375849 392720
rect 375883 392717 375895 392751
rect 375837 392711 375895 392717
rect 375929 392751 375987 392757
rect 375929 392717 375941 392751
rect 375975 392748 375987 392751
rect 379974 392748 379980 392760
rect 375975 392720 379980 392748
rect 375975 392717 375987 392720
rect 375929 392711 375987 392717
rect 379974 392708 379980 392720
rect 380032 392708 380038 392760
rect 281350 392640 281356 392692
rect 281408 392680 281414 392692
rect 379701 392683 379759 392689
rect 379701 392680 379713 392683
rect 281408 392652 379713 392680
rect 281408 392640 281414 392652
rect 379701 392649 379713 392652
rect 379747 392649 379759 392683
rect 379701 392643 379759 392649
rect 277210 392572 277216 392624
rect 277268 392612 277274 392624
rect 379609 392615 379667 392621
rect 379609 392612 379621 392615
rect 277268 392584 379621 392612
rect 277268 392572 277274 392584
rect 379609 392581 379621 392584
rect 379655 392581 379667 392615
rect 379609 392575 379667 392581
rect 302050 392504 302056 392556
rect 302108 392544 302114 392556
rect 375745 392547 375803 392553
rect 375745 392544 375757 392547
rect 302108 392516 375757 392544
rect 302108 392504 302114 392516
rect 375745 392513 375757 392516
rect 375791 392513 375803 392547
rect 375745 392507 375803 392513
rect 375837 392547 375895 392553
rect 375837 392513 375849 392547
rect 375883 392544 375895 392547
rect 380084 392544 380112 392788
rect 380710 392748 380716 392760
rect 380671 392720 380716 392748
rect 380710 392708 380716 392720
rect 380768 392708 380774 392760
rect 380802 392708 380808 392760
rect 380860 392708 380866 392760
rect 375883 392516 380112 392544
rect 375883 392513 375895 392516
rect 375837 392507 375895 392513
rect 300670 392436 300676 392488
rect 300728 392476 300734 392488
rect 376021 392479 376079 392485
rect 376021 392476 376033 392479
rect 300728 392448 376033 392476
rect 300728 392436 300734 392448
rect 376021 392445 376033 392448
rect 376067 392445 376079 392479
rect 376021 392439 376079 392445
rect 308950 392368 308956 392420
rect 309008 392408 309014 392420
rect 377217 392411 377275 392417
rect 377217 392408 377229 392411
rect 309008 392380 377229 392408
rect 309008 392368 309014 392380
rect 377217 392377 377229 392380
rect 377263 392377 377275 392411
rect 377217 392371 377275 392377
rect 314562 392300 314568 392352
rect 314620 392340 314626 392352
rect 375653 392343 375711 392349
rect 375653 392340 375665 392343
rect 314620 392312 375665 392340
rect 314620 392300 314626 392312
rect 375653 392309 375665 392312
rect 375699 392309 375711 392343
rect 375653 392303 375711 392309
rect 375745 392343 375803 392349
rect 375745 392309 375757 392343
rect 375791 392340 375803 392343
rect 380820 392340 380848 392708
rect 375791 392312 380848 392340
rect 375791 392309 375803 392312
rect 375745 392303 375803 392309
rect 322842 392232 322848 392284
rect 322900 392272 322906 392284
rect 379425 392275 379483 392281
rect 379425 392272 379437 392275
rect 322900 392244 379437 392272
rect 322900 392232 322906 392244
rect 379425 392241 379437 392244
rect 379471 392241 379483 392275
rect 379425 392235 379483 392241
rect 375653 392207 375711 392213
rect 375653 392173 375665 392207
rect 375699 392204 375711 392207
rect 380713 392207 380771 392213
rect 380713 392204 380725 392207
rect 375699 392176 380725 392204
rect 375699 392173 375711 392176
rect 375653 392167 375711 392173
rect 380713 392173 380725 392176
rect 380759 392173 380771 392207
rect 380713 392167 380771 392173
rect 302878 391212 302884 391264
rect 302936 391252 302942 391264
rect 357434 391252 357440 391264
rect 302936 391224 357440 391252
rect 302936 391212 302942 391224
rect 357434 391212 357440 391224
rect 357492 391212 357498 391264
rect 416590 389376 416596 389428
rect 416648 389416 416654 389428
rect 464246 389416 464252 389428
rect 416648 389388 464252 389416
rect 416648 389376 416654 389388
rect 464246 389376 464252 389388
rect 464304 389376 464310 389428
rect 418062 389308 418068 389360
rect 418120 389348 418126 389360
rect 487430 389348 487436 389360
rect 418120 389320 487436 389348
rect 418120 389308 418126 389320
rect 487430 389308 487436 389320
rect 487488 389308 487494 389360
rect 401502 389240 401508 389292
rect 401560 389280 401566 389292
rect 475838 389280 475844 389292
rect 401560 389252 475844 389280
rect 401560 389240 401566 389252
rect 475838 389240 475844 389252
rect 475896 389240 475902 389292
rect 416682 389172 416688 389224
rect 416740 389212 416746 389224
rect 499022 389212 499028 389224
rect 416740 389184 499028 389212
rect 416740 389172 416746 389184
rect 499022 389172 499028 389184
rect 499080 389172 499086 389224
rect 153286 389144 153292 389156
rect 153247 389116 153292 389144
rect 153286 389104 153292 389116
rect 153344 389104 153350 389156
rect 351822 387812 351828 387864
rect 351880 387852 351886 387864
rect 357434 387852 357440 387864
rect 351880 387824 357440 387852
rect 351880 387812 351886 387824
rect 357434 387812 357440 387824
rect 357492 387812 357498 387864
rect 357342 386560 357348 386572
rect 357303 386532 357348 386560
rect 357342 386520 357348 386532
rect 357400 386520 357406 386572
rect 128630 386384 128636 386436
rect 128688 386424 128694 386436
rect 128906 386424 128912 386436
rect 128688 386396 128912 386424
rect 128688 386384 128694 386396
rect 128906 386384 128912 386396
rect 128964 386384 128970 386436
rect 133966 386424 133972 386436
rect 133927 386396 133972 386424
rect 133966 386384 133972 386396
rect 134024 386384 134030 386436
rect 297450 386424 297456 386436
rect 297411 386396 297456 386424
rect 297450 386384 297456 386396
rect 297508 386384 297514 386436
rect 299569 386427 299627 386433
rect 299569 386393 299581 386427
rect 299615 386424 299627 386427
rect 299658 386424 299664 386436
rect 299615 386396 299664 386424
rect 299615 386393 299627 386396
rect 299569 386387 299627 386393
rect 299658 386384 299664 386396
rect 299716 386384 299722 386436
rect 357342 386356 357348 386368
rect 357303 386328 357348 386356
rect 357342 386316 357348 386328
rect 357400 386316 357406 386368
rect 133966 386288 133972 386300
rect 133927 386260 133972 386288
rect 133966 386248 133972 386260
rect 134024 386248 134030 386300
rect 284021 383707 284079 383713
rect 284021 383673 284033 383707
rect 284067 383704 284079 383707
rect 284110 383704 284116 383716
rect 284067 383676 284116 383704
rect 284067 383673 284079 383676
rect 284021 383667 284079 383673
rect 284110 383664 284116 383676
rect 284168 383664 284174 383716
rect 297450 383500 297456 383512
rect 297411 383472 297456 383500
rect 297450 383460 297456 383472
rect 297508 383460 297514 383512
rect 351178 380876 351184 380928
rect 351236 380916 351242 380928
rect 357434 380916 357440 380928
rect 351236 380888 357440 380916
rect 351236 380876 351242 380888
rect 357434 380876 357440 380888
rect 357492 380876 357498 380928
rect 153286 379448 153292 379500
rect 153344 379488 153350 379500
rect 153470 379488 153476 379500
rect 153344 379460 153476 379488
rect 153344 379448 153350 379460
rect 153470 379448 153476 379460
rect 153528 379448 153534 379500
rect 133969 376771 134027 376777
rect 133969 376737 133981 376771
rect 134015 376768 134027 376771
rect 134150 376768 134156 376780
rect 134015 376740 134156 376768
rect 134015 376737 134027 376740
rect 133969 376731 134027 376737
rect 134150 376728 134156 376740
rect 134208 376728 134214 376780
rect 357158 376728 357164 376780
rect 357216 376768 357222 376780
rect 357345 376771 357403 376777
rect 357345 376768 357357 376771
rect 357216 376740 357357 376768
rect 357216 376728 357222 376740
rect 357345 376737 357357 376740
rect 357391 376737 357403 376771
rect 357345 376731 357403 376737
rect 357250 376592 357256 376644
rect 357308 376632 357314 376644
rect 357345 376635 357403 376641
rect 357345 376632 357357 376635
rect 357308 376604 357357 376632
rect 357308 376592 357314 376604
rect 357345 376601 357357 376604
rect 357391 376601 357403 376635
rect 357345 376595 357403 376601
rect 297453 375411 297511 375417
rect 297453 375377 297465 375411
rect 297499 375408 297511 375411
rect 297634 375408 297640 375420
rect 297499 375380 297640 375408
rect 297499 375377 297511 375380
rect 297453 375371 297511 375377
rect 297634 375368 297640 375380
rect 297692 375368 297698 375420
rect 128814 375340 128820 375352
rect 128775 375312 128820 375340
rect 128814 375300 128820 375312
rect 128872 375300 128878 375352
rect 333882 374008 333888 374060
rect 333940 374048 333946 374060
rect 357434 374048 357440 374060
rect 333940 374020 357440 374048
rect 333940 374008 333946 374020
rect 357434 374008 357440 374020
rect 357492 374008 357498 374060
rect 413922 374008 413928 374060
rect 413980 374048 413986 374060
rect 456794 374048 456800 374060
rect 413980 374020 456800 374048
rect 413980 374008 413986 374020
rect 456794 374008 456800 374020
rect 456852 374008 456858 374060
rect 297542 370512 297548 370524
rect 297503 370484 297548 370512
rect 297542 370472 297548 370484
rect 297600 370472 297606 370524
rect 357342 367112 357348 367124
rect 357303 367084 357348 367112
rect 357342 367072 357348 367084
rect 357400 367072 357406 367124
rect 153562 367044 153568 367056
rect 153523 367016 153568 367044
rect 153562 367004 153568 367016
rect 153620 367004 153626 367056
rect 284021 367047 284079 367053
rect 284021 367013 284033 367047
rect 284067 367044 284079 367047
rect 284110 367044 284116 367056
rect 284067 367016 284116 367044
rect 284067 367013 284079 367016
rect 284021 367007 284079 367013
rect 284110 367004 284116 367016
rect 284168 367004 284174 367056
rect 390554 367004 390560 367056
rect 390612 367004 390618 367056
rect 390572 366976 390600 367004
rect 390738 366976 390744 366988
rect 390572 366948 390744 366976
rect 390738 366936 390744 366948
rect 390796 366936 390802 366988
rect 2774 365712 2780 365764
rect 2832 365752 2838 365764
rect 5166 365752 5172 365764
rect 2832 365724 5172 365752
rect 2832 365712 2838 365724
rect 5166 365712 5172 365724
rect 5224 365712 5230 365764
rect 128814 365752 128820 365764
rect 128775 365724 128820 365752
rect 128814 365712 128820 365724
rect 128872 365712 128878 365764
rect 129366 365644 129372 365696
rect 129424 365684 129430 365696
rect 197722 365684 197728 365696
rect 129424 365656 197728 365684
rect 129424 365644 129430 365656
rect 197722 365644 197728 365656
rect 197780 365644 197786 365696
rect 358538 364352 358544 364404
rect 358596 364392 358602 364404
rect 358722 364392 358728 364404
rect 358596 364364 358728 364392
rect 358596 364352 358602 364364
rect 358722 364352 358728 364364
rect 358780 364352 358786 364404
rect 299658 362284 299664 362296
rect 299619 362256 299664 362284
rect 299658 362244 299664 362256
rect 299716 362244 299722 362296
rect 360010 360136 360016 360188
rect 360068 360176 360074 360188
rect 364518 360176 364524 360188
rect 360068 360148 364524 360176
rect 360068 360136 360074 360148
rect 364518 360136 364524 360148
rect 364576 360136 364582 360188
rect 360102 360068 360108 360120
rect 360160 360108 360166 360120
rect 365714 360108 365720 360120
rect 360160 360080 365720 360108
rect 360160 360068 360166 360080
rect 365714 360068 365720 360080
rect 365772 360068 365778 360120
rect 126514 358708 126520 358760
rect 126572 358748 126578 358760
rect 128906 358748 128912 358760
rect 126572 358720 128912 358748
rect 126572 358708 126578 358720
rect 128906 358708 128912 358720
rect 128964 358708 128970 358760
rect 360102 358640 360108 358692
rect 360160 358680 360166 358692
rect 367370 358680 367376 358692
rect 360160 358652 367376 358680
rect 360160 358640 360166 358652
rect 367370 358640 367376 358652
rect 367428 358640 367434 358692
rect 359458 358572 359464 358624
rect 359516 358612 359522 358624
rect 369578 358612 369584 358624
rect 359516 358584 369584 358612
rect 359516 358572 359522 358584
rect 369578 358572 369584 358584
rect 369636 358572 369642 358624
rect 363690 358504 363696 358556
rect 363748 358544 363754 358556
rect 374178 358544 374184 358556
rect 363748 358516 374184 358544
rect 363748 358504 363754 358516
rect 374178 358504 374184 358516
rect 374236 358504 374242 358556
rect 362862 358436 362868 358488
rect 362920 358476 362926 358488
rect 378778 358476 378784 358488
rect 362920 358448 378784 358476
rect 362920 358436 362926 358448
rect 378778 358436 378784 358448
rect 378836 358436 378842 358488
rect 362218 358368 362224 358420
rect 362276 358408 362282 358420
rect 383378 358408 383384 358420
rect 362276 358380 383384 358408
rect 362276 358368 362282 358380
rect 383378 358368 383384 358380
rect 383436 358368 383442 358420
rect 354582 358300 354588 358352
rect 354640 358340 354646 358352
rect 376570 358340 376576 358352
rect 354640 358312 376576 358340
rect 354640 358300 354646 358312
rect 376570 358300 376576 358312
rect 376628 358300 376634 358352
rect 350442 358232 350448 358284
rect 350500 358272 350506 358284
rect 371970 358272 371976 358284
rect 350500 358244 371976 358272
rect 350500 358232 350506 358244
rect 371970 358232 371976 358244
rect 372028 358232 372034 358284
rect 342162 358164 342168 358216
rect 342220 358204 342226 358216
rect 364978 358204 364984 358216
rect 342220 358176 364984 358204
rect 342220 358164 342226 358176
rect 364978 358164 364984 358176
rect 365036 358164 365042 358216
rect 361482 358096 361488 358148
rect 361540 358136 361546 358148
rect 390370 358136 390376 358148
rect 361540 358108 390376 358136
rect 361540 358096 361546 358108
rect 390370 358096 390376 358108
rect 390428 358096 390434 358148
rect 333790 358028 333796 358080
rect 333848 358068 333854 358080
rect 387978 358068 387984 358080
rect 333848 358040 387984 358068
rect 333848 358028 333854 358040
rect 387978 358028 387984 358040
rect 388036 358028 388042 358080
rect 297726 357688 297732 357740
rect 297784 357688 297790 357740
rect 297744 357468 297772 357688
rect 153565 357459 153623 357465
rect 153565 357425 153577 357459
rect 153611 357456 153623 357459
rect 153654 357456 153660 357468
rect 153611 357428 153660 357456
rect 153611 357425 153623 357428
rect 153565 357419 153623 357425
rect 153654 357416 153660 357428
rect 153712 357416 153718 357468
rect 284018 357456 284024 357468
rect 283979 357428 284024 357456
rect 284018 357416 284024 357428
rect 284076 357416 284082 357468
rect 297545 357459 297603 357465
rect 297545 357425 297557 357459
rect 297591 357456 297603 357459
rect 297634 357456 297640 357468
rect 297591 357428 297640 357456
rect 297591 357425 297603 357428
rect 297545 357419 297603 357425
rect 297634 357416 297640 357428
rect 297692 357416 297698 357468
rect 297726 357416 297732 357468
rect 297784 357416 297790 357468
rect 299661 357459 299719 357465
rect 299661 357425 299673 357459
rect 299707 357456 299719 357459
rect 299750 357456 299756 357468
rect 299707 357428 299756 357456
rect 299707 357425 299719 357428
rect 299661 357419 299719 357425
rect 299750 357416 299756 357428
rect 299808 357416 299814 357468
rect 362770 357416 362776 357468
rect 362828 357456 362834 357468
rect 363598 357456 363604 357468
rect 362828 357428 363604 357456
rect 362828 357416 362834 357428
rect 363598 357416 363604 357428
rect 363656 357416 363662 357468
rect 412542 357416 412548 357468
rect 412600 357456 412606 357468
rect 456794 357456 456800 357468
rect 412600 357428 456800 357456
rect 412600 357416 412606 357428
rect 456794 357416 456800 357428
rect 456852 357416 456858 357468
rect 134242 357388 134248 357400
rect 134203 357360 134248 357388
rect 134242 357348 134248 357360
rect 134300 357348 134306 357400
rect 390738 357348 390744 357400
rect 390796 357388 390802 357400
rect 390922 357388 390928 357400
rect 390796 357360 390928 357388
rect 390796 357348 390802 357360
rect 390922 357348 390928 357360
rect 390980 357348 390986 357400
rect 185578 355988 185584 356040
rect 185636 356028 185642 356040
rect 188338 356028 188344 356040
rect 185636 356000 188344 356028
rect 185636 355988 185642 356000
rect 188338 355988 188344 356000
rect 188396 355988 188402 356040
rect 297545 356031 297603 356037
rect 297545 355997 297557 356031
rect 297591 356028 297603 356031
rect 297634 356028 297640 356040
rect 297591 356000 297640 356028
rect 297591 355997 297603 356000
rect 297545 355991 297603 355997
rect 297634 355988 297640 356000
rect 297692 355988 297698 356040
rect 390922 356028 390928 356040
rect 390883 356000 390928 356028
rect 390922 355988 390928 356000
rect 390980 355988 390986 356040
rect 267274 355308 267280 355360
rect 267332 355348 267338 355360
rect 436094 355348 436100 355360
rect 267332 355320 436100 355348
rect 267332 355308 267338 355320
rect 436094 355308 436100 355320
rect 436152 355308 436158 355360
rect 128998 350956 129004 351008
rect 129056 350996 129062 351008
rect 130378 350996 130384 351008
rect 129056 350968 130384 350996
rect 129056 350956 129062 350968
rect 130378 350956 130384 350968
rect 130436 350956 130442 351008
rect 134242 347800 134248 347812
rect 134203 347772 134248 347800
rect 134242 347760 134248 347772
rect 134300 347760 134306 347812
rect 153470 347760 153476 347812
rect 153528 347800 153534 347812
rect 153562 347800 153568 347812
rect 153528 347772 153568 347800
rect 153528 347760 153534 347772
rect 153562 347760 153568 347772
rect 153620 347760 153626 347812
rect 128814 347732 128820 347744
rect 128775 347704 128820 347732
rect 128814 347692 128820 347704
rect 128872 347692 128878 347744
rect 284021 347735 284079 347741
rect 284021 347701 284033 347735
rect 284067 347732 284079 347735
rect 284110 347732 284116 347744
rect 284067 347704 284116 347732
rect 284067 347701 284079 347704
rect 284021 347695 284079 347701
rect 284110 347692 284116 347704
rect 284168 347692 284174 347744
rect 297542 346440 297548 346452
rect 297503 346412 297548 346440
rect 297542 346400 297548 346412
rect 297600 346400 297606 346452
rect 390922 346440 390928 346452
rect 390883 346412 390928 346440
rect 390922 346400 390928 346412
rect 390980 346400 390986 346452
rect 358538 345040 358544 345092
rect 358596 345080 358602 345092
rect 358722 345080 358728 345092
rect 358596 345052 358728 345080
rect 358596 345040 358602 345052
rect 358722 345040 358728 345052
rect 358780 345040 358786 345092
rect 504818 345040 504824 345092
rect 504876 345080 504882 345092
rect 579982 345080 579988 345092
rect 504876 345052 579988 345080
rect 504876 345040 504882 345052
rect 579982 345040 579988 345052
rect 580040 345040 580046 345092
rect 132954 342864 132960 342916
rect 133012 342904 133018 342916
rect 192478 342904 192484 342916
rect 133012 342876 192484 342904
rect 133012 342864 133018 342876
rect 192478 342864 192484 342876
rect 192536 342864 192542 342916
rect 199286 342864 199292 342916
rect 199344 342904 199350 342916
rect 200206 342904 200212 342916
rect 199344 342876 200212 342904
rect 199344 342864 199350 342876
rect 200206 342864 200212 342876
rect 200264 342864 200270 342916
rect 128814 342456 128820 342508
rect 128872 342496 128878 342508
rect 132954 342496 132960 342508
rect 128872 342468 132960 342496
rect 128872 342456 128878 342468
rect 132954 342456 132960 342468
rect 133012 342456 133018 342508
rect 503806 341980 503812 342032
rect 503864 342020 503870 342032
rect 504174 342020 504180 342032
rect 503864 341992 504180 342020
rect 503864 341980 503870 341992
rect 504174 341980 504180 341992
rect 504232 341980 504238 342032
rect 131942 341640 131948 341692
rect 132000 341680 132006 341692
rect 580626 341680 580632 341692
rect 132000 341652 580632 341680
rect 132000 341640 132006 341652
rect 580626 341640 580632 341652
rect 580684 341640 580690 341692
rect 132034 341572 132040 341624
rect 132092 341612 132098 341624
rect 580810 341612 580816 341624
rect 132092 341584 580816 341612
rect 132092 341572 132098 341584
rect 580810 341572 580816 341584
rect 580868 341572 580874 341624
rect 131666 341504 131672 341556
rect 131724 341544 131730 341556
rect 580718 341544 580724 341556
rect 131724 341516 580724 341544
rect 131724 341504 131730 341516
rect 580718 341504 580724 341516
rect 580776 341504 580782 341556
rect 390922 340892 390928 340944
rect 390980 340892 390986 340944
rect 127158 340824 127164 340876
rect 127216 340864 127222 340876
rect 385034 340864 385040 340876
rect 127216 340836 385040 340864
rect 127216 340824 127222 340836
rect 385034 340824 385040 340836
rect 385092 340824 385098 340876
rect 390830 340824 390836 340876
rect 390888 340864 390894 340876
rect 390940 340864 390968 340892
rect 504726 340864 504732 340876
rect 390888 340836 390968 340864
rect 504100 340836 504732 340864
rect 390888 340824 390894 340836
rect 127250 340756 127256 340808
rect 127308 340796 127314 340808
rect 380894 340796 380900 340808
rect 127308 340768 380900 340796
rect 127308 340756 127314 340768
rect 380894 340756 380900 340768
rect 380952 340756 380958 340808
rect 503898 340756 503904 340808
rect 503956 340796 503962 340808
rect 504100 340796 504128 340836
rect 504726 340824 504732 340836
rect 504784 340824 504790 340876
rect 503956 340768 504128 340796
rect 503956 340756 503962 340768
rect 126882 340688 126888 340740
rect 126940 340728 126946 340740
rect 358170 340728 358176 340740
rect 126940 340700 358176 340728
rect 126940 340688 126946 340700
rect 358170 340688 358176 340700
rect 358228 340688 358234 340740
rect 128814 340620 128820 340672
rect 128872 340660 128878 340672
rect 360194 340660 360200 340672
rect 128872 340632 360200 340660
rect 128872 340620 128878 340632
rect 360194 340620 360200 340632
rect 360252 340620 360258 340672
rect 127710 340552 127716 340604
rect 127768 340592 127774 340604
rect 358078 340592 358084 340604
rect 127768 340564 358084 340592
rect 127768 340552 127774 340564
rect 358078 340552 358084 340564
rect 358136 340552 358142 340604
rect 128817 340527 128875 340533
rect 128817 340493 128829 340527
rect 128863 340524 128875 340527
rect 128906 340524 128912 340536
rect 128863 340496 128912 340524
rect 128863 340493 128875 340496
rect 128817 340487 128875 340493
rect 128906 340484 128912 340496
rect 128964 340484 128970 340536
rect 111702 340212 111708 340264
rect 111760 340252 111766 340264
rect 127158 340252 127164 340264
rect 111760 340224 127164 340252
rect 111760 340212 111766 340224
rect 127158 340212 127164 340224
rect 127216 340212 127222 340264
rect 110322 340144 110328 340196
rect 110380 340184 110386 340196
rect 127250 340184 127256 340196
rect 110380 340156 127256 340184
rect 110380 340144 110386 340156
rect 127250 340144 127256 340156
rect 127308 340144 127314 340196
rect 126054 340076 126060 340128
rect 126112 340116 126118 340128
rect 126882 340116 126888 340128
rect 126112 340088 126888 340116
rect 126112 340076 126118 340088
rect 126882 340076 126888 340088
rect 126940 340076 126946 340128
rect 198090 338988 198096 339040
rect 198148 339028 198154 339040
rect 209958 339028 209964 339040
rect 198148 339000 209964 339028
rect 198148 338988 198154 339000
rect 209958 338988 209964 339000
rect 210016 338988 210022 339040
rect 199470 338920 199476 338972
rect 199528 338960 199534 338972
rect 214098 338960 214104 338972
rect 199528 338932 214104 338960
rect 199528 338920 199534 338932
rect 214098 338920 214104 338932
rect 214156 338920 214162 338972
rect 257706 338920 257712 338972
rect 257764 338960 257770 338972
rect 267550 338960 267556 338972
rect 257764 338932 267556 338960
rect 257764 338920 257770 338932
rect 267550 338920 267556 338932
rect 267608 338920 267614 338972
rect 199378 338852 199384 338904
rect 199436 338892 199442 338904
rect 215294 338892 215300 338904
rect 199436 338864 215300 338892
rect 199436 338852 199442 338864
rect 215294 338852 215300 338864
rect 215352 338852 215358 338904
rect 253658 338852 253664 338904
rect 253716 338892 253722 338904
rect 268838 338892 268844 338904
rect 253716 338864 268844 338892
rect 253716 338852 253722 338864
rect 268838 338852 268844 338864
rect 268896 338852 268902 338904
rect 198182 338784 198188 338836
rect 198240 338824 198246 338836
rect 220814 338824 220820 338836
rect 198240 338796 220820 338824
rect 198240 338784 198246 338796
rect 220814 338784 220820 338796
rect 220872 338784 220878 338836
rect 244182 338784 244188 338836
rect 244240 338824 244246 338836
rect 267458 338824 267464 338836
rect 244240 338796 267464 338824
rect 244240 338784 244246 338796
rect 267458 338784 267464 338796
rect 267516 338784 267522 338836
rect 198274 338716 198280 338768
rect 198332 338756 198338 338768
rect 222194 338756 222200 338768
rect 198332 338728 222200 338756
rect 198332 338716 198338 338728
rect 222194 338716 222200 338728
rect 222252 338716 222258 338768
rect 237282 338716 237288 338768
rect 237340 338756 237346 338768
rect 267366 338756 267372 338768
rect 237340 338728 267372 338756
rect 237340 338716 237346 338728
rect 267366 338716 267372 338728
rect 267424 338716 267430 338768
rect 262122 338376 262128 338428
rect 262180 338416 262186 338428
rect 268930 338416 268936 338428
rect 262180 338388 268936 338416
rect 262180 338376 262186 338388
rect 268930 338376 268936 338388
rect 268988 338376 268994 338428
rect 284018 338212 284024 338224
rect 283979 338184 284024 338212
rect 284018 338172 284024 338184
rect 284076 338172 284082 338224
rect 153378 338104 153384 338156
rect 153436 338144 153442 338156
rect 153562 338144 153568 338156
rect 153436 338116 153568 338144
rect 153436 338104 153442 338116
rect 153562 338104 153568 338116
rect 153620 338104 153626 338156
rect 107562 338036 107568 338088
rect 107620 338076 107626 338088
rect 283929 338079 283987 338085
rect 283929 338076 283941 338079
rect 107620 338048 283941 338076
rect 107620 338036 107626 338048
rect 283929 338045 283941 338048
rect 283975 338045 283987 338079
rect 283929 338039 283987 338045
rect 284018 338036 284024 338088
rect 284076 338036 284082 338088
rect 284205 338079 284263 338085
rect 284205 338045 284217 338079
rect 284251 338076 284263 338079
rect 302878 338076 302884 338088
rect 284251 338048 302884 338076
rect 284251 338045 284263 338048
rect 284205 338039 284263 338045
rect 302878 338036 302884 338048
rect 302936 338036 302942 338088
rect 97902 337968 97908 338020
rect 97960 338008 97966 338020
rect 126974 338008 126980 338020
rect 97960 337980 126980 338008
rect 97960 337968 97966 337980
rect 126974 337968 126980 337980
rect 127032 337968 127038 338020
rect 128906 338008 128912 338020
rect 128867 337980 128912 338008
rect 128906 337968 128912 337980
rect 128964 337968 128970 338020
rect 231854 337968 231860 338020
rect 231912 338008 231918 338020
rect 248690 338008 248696 338020
rect 231912 337980 248696 338008
rect 231912 337968 231918 337980
rect 248690 337968 248696 337980
rect 248748 337968 248754 338020
rect 284036 338008 284064 338036
rect 284113 338011 284171 338017
rect 284113 338008 284125 338011
rect 284036 337980 284125 338008
rect 284113 337977 284125 337980
rect 284159 337977 284171 338011
rect 284113 337971 284171 337977
rect 87782 337900 87788 337952
rect 87840 337940 87846 337952
rect 96525 337943 96583 337949
rect 96525 337940 96537 337943
rect 87840 337912 96537 337940
rect 87840 337900 87846 337912
rect 96525 337909 96537 337912
rect 96571 337909 96583 337943
rect 96525 337903 96583 337909
rect 113082 337900 113088 337952
rect 113140 337940 113146 337952
rect 127066 337940 127072 337952
rect 113140 337912 127072 337940
rect 113140 337900 113146 337912
rect 127066 337900 127072 337912
rect 127124 337900 127130 337952
rect 220446 337900 220452 337952
rect 220504 337940 220510 337952
rect 238110 337940 238116 337952
rect 220504 337912 238116 337940
rect 220504 337900 220510 337912
rect 238110 337900 238116 337912
rect 238168 337900 238174 337952
rect 122742 337832 122748 337884
rect 122800 337872 122806 337884
rect 127710 337872 127716 337884
rect 122800 337844 127716 337872
rect 122800 337832 122806 337844
rect 127710 337832 127716 337844
rect 127768 337832 127774 337884
rect 209038 337832 209044 337884
rect 209096 337872 209102 337884
rect 220078 337872 220084 337884
rect 209096 337844 220084 337872
rect 209096 337832 209102 337844
rect 220078 337832 220084 337844
rect 220136 337832 220142 337884
rect 226150 337832 226156 337884
rect 226208 337872 226214 337884
rect 248506 337872 248512 337884
rect 226208 337844 248512 337872
rect 226208 337832 226214 337844
rect 248506 337832 248512 337844
rect 248564 337832 248570 337884
rect 250990 337832 250996 337884
rect 251048 337872 251054 337884
rect 260190 337872 260196 337884
rect 251048 337844 260196 337872
rect 251048 337832 251054 337844
rect 260190 337832 260196 337844
rect 260248 337832 260254 337884
rect 203334 337764 203340 337816
rect 203392 337804 203398 337816
rect 215938 337804 215944 337816
rect 203392 337776 215944 337804
rect 203392 337764 203398 337776
rect 215938 337764 215944 337776
rect 215996 337764 216002 337816
rect 217502 337764 217508 337816
rect 217560 337804 217566 337816
rect 241333 337807 241391 337813
rect 241333 337804 241345 337807
rect 217560 337776 241345 337804
rect 217560 337764 217566 337776
rect 241333 337773 241345 337776
rect 241379 337773 241391 337807
rect 241333 337767 241391 337773
rect 241422 337764 241428 337816
rect 241480 337804 241486 337816
rect 246022 337804 246028 337816
rect 241480 337776 246028 337804
rect 241480 337764 241486 337776
rect 246022 337764 246028 337776
rect 246080 337764 246086 337816
rect 253750 337764 253756 337816
rect 253808 337804 253814 337816
rect 263134 337804 263140 337816
rect 253808 337776 263140 337804
rect 253808 337764 253814 337776
rect 263134 337764 263140 337776
rect 263192 337764 263198 337816
rect 96525 337739 96583 337745
rect 96525 337705 96537 337739
rect 96571 337736 96583 337739
rect 96571 337708 99328 337736
rect 96571 337705 96583 337708
rect 96525 337699 96583 337705
rect 99300 337668 99328 337708
rect 200574 337696 200580 337748
rect 200632 337736 200638 337748
rect 238018 337736 238024 337748
rect 200632 337708 238024 337736
rect 200632 337696 200638 337708
rect 238018 337696 238024 337708
rect 238076 337696 238082 337748
rect 240042 337696 240048 337748
rect 240100 337736 240106 337748
rect 243078 337736 243084 337748
rect 240100 337708 243084 337736
rect 240100 337696 240106 337708
rect 243078 337696 243084 337708
rect 243136 337696 243142 337748
rect 247678 337696 247684 337748
rect 247736 337736 247742 337748
rect 257430 337736 257436 337748
rect 247736 337708 257436 337736
rect 247736 337696 247742 337708
rect 257430 337696 257436 337708
rect 257488 337696 257494 337748
rect 99377 337671 99435 337677
rect 99377 337668 99389 337671
rect 99300 337640 99389 337668
rect 99377 337637 99389 337640
rect 99423 337637 99435 337671
rect 99377 337631 99435 337637
rect 106277 337671 106335 337677
rect 106277 337637 106289 337671
rect 106323 337668 106335 337671
rect 117222 337668 117228 337680
rect 106323 337640 117228 337668
rect 106323 337637 106335 337640
rect 106277 337631 106335 337637
rect 117222 337628 117228 337640
rect 117280 337668 117286 337680
rect 126422 337668 126428 337680
rect 117280 337640 126428 337668
rect 117280 337628 117286 337640
rect 126422 337628 126428 337640
rect 126480 337628 126486 337680
rect 214742 337628 214748 337680
rect 214800 337668 214806 337680
rect 258718 337668 258724 337680
rect 214800 337640 258724 337668
rect 214800 337628 214806 337640
rect 258718 337628 258724 337640
rect 258776 337628 258782 337680
rect 206094 337560 206100 337612
rect 206152 337600 206158 337612
rect 255314 337600 255320 337612
rect 206152 337572 255320 337600
rect 206152 337560 206158 337572
rect 255314 337560 255320 337572
rect 255372 337560 255378 337612
rect 401410 337560 401416 337612
rect 401468 337600 401474 337612
rect 460566 337600 460572 337612
rect 401468 337572 460572 337600
rect 401468 337560 401474 337572
rect 460566 337560 460572 337572
rect 460624 337560 460630 337612
rect 99377 337535 99435 337541
rect 99377 337501 99389 337535
rect 99423 337532 99435 337535
rect 106277 337535 106335 337541
rect 106277 337532 106289 337535
rect 99423 337504 106289 337532
rect 99423 337501 99435 337504
rect 99377 337495 99435 337501
rect 106277 337501 106289 337504
rect 106323 337501 106335 337535
rect 106277 337495 106335 337501
rect 117958 337492 117964 337544
rect 118016 337532 118022 337544
rect 132678 337532 132684 337544
rect 118016 337504 132684 337532
rect 118016 337492 118022 337504
rect 132678 337492 132684 337504
rect 132736 337532 132742 337544
rect 297358 337532 297364 337544
rect 132736 337504 297364 337532
rect 132736 337492 132742 337504
rect 297358 337492 297364 337504
rect 297416 337492 297422 337544
rect 411162 337492 411168 337544
rect 411220 337532 411226 337544
rect 472158 337532 472164 337544
rect 411220 337504 472164 337532
rect 411220 337492 411226 337504
rect 472158 337492 472164 337504
rect 472216 337492 472222 337544
rect 72878 337424 72884 337476
rect 72936 337464 72942 337476
rect 103422 337464 103428 337476
rect 72936 337436 103428 337464
rect 72936 337424 72942 337436
rect 103422 337424 103428 337436
rect 103480 337464 103486 337476
rect 299750 337464 299756 337476
rect 103480 337436 299756 337464
rect 103480 337424 103486 337436
rect 299750 337424 299756 337436
rect 299808 337424 299814 337476
rect 408402 337424 408408 337476
rect 408460 337464 408466 337476
rect 483750 337464 483756 337476
rect 408460 337436 483756 337464
rect 408460 337424 408466 337436
rect 483750 337424 483756 337436
rect 483808 337424 483814 337476
rect 77846 337356 77852 337408
rect 77904 337396 77910 337408
rect 100662 337396 100668 337408
rect 77904 337368 100668 337396
rect 77904 337356 77910 337368
rect 100662 337356 100668 337368
rect 100720 337396 100726 337408
rect 329834 337396 329840 337408
rect 100720 337368 329840 337396
rect 100720 337356 100726 337368
rect 329834 337356 329840 337368
rect 329892 337356 329898 337408
rect 413830 337356 413836 337408
rect 413888 337396 413894 337408
rect 495342 337396 495348 337408
rect 413888 337368 495348 337396
rect 413888 337356 413894 337368
rect 495342 337356 495348 337368
rect 495400 337356 495406 337408
rect 228910 337288 228916 337340
rect 228968 337328 228974 337340
rect 232498 337328 232504 337340
rect 228968 337300 232504 337328
rect 228968 337288 228974 337300
rect 232498 337288 232504 337300
rect 232556 337288 232562 337340
rect 241333 337331 241391 337337
rect 241333 337297 241345 337331
rect 241379 337328 241391 337331
rect 244918 337328 244924 337340
rect 241379 337300 244924 337328
rect 241379 337297 241391 337300
rect 241333 337291 241391 337297
rect 244918 337288 244924 337300
rect 244976 337288 244982 337340
rect 237558 337220 237564 337272
rect 237616 337260 237622 337272
rect 243078 337260 243084 337272
rect 237616 337232 243084 337260
rect 237616 337220 237622 337232
rect 243078 337220 243084 337232
rect 243136 337220 243142 337272
rect 234614 337084 234620 337136
rect 234672 337124 234678 337136
rect 237742 337124 237748 337136
rect 234672 337096 237748 337124
rect 234672 337084 234678 337096
rect 237742 337084 237748 337096
rect 237800 337084 237806 337136
rect 251726 337084 251732 337136
rect 251784 337124 251790 337136
rect 252462 337124 252468 337136
rect 251784 337096 252468 337124
rect 251784 337084 251790 337096
rect 252462 337084 252468 337096
rect 252520 337084 252526 337136
rect 92750 336812 92756 336864
rect 92808 336852 92814 336864
rect 93762 336852 93768 336864
rect 92808 336824 93768 336852
rect 92808 336812 92814 336824
rect 93762 336812 93768 336824
rect 93820 336812 93826 336864
rect 102870 336812 102876 336864
rect 102928 336852 102934 336864
rect 103330 336852 103336 336864
rect 102928 336824 103336 336852
rect 102928 336812 102934 336824
rect 103330 336812 103336 336824
rect 103388 336812 103394 336864
rect 223206 336812 223212 336864
rect 223264 336852 223270 336864
rect 229738 336852 229744 336864
rect 223264 336824 229744 336852
rect 223264 336812 223270 336824
rect 229738 336812 229744 336824
rect 229796 336812 229802 336864
rect 244090 336812 244096 336864
rect 244148 336852 244154 336864
rect 248782 336852 248788 336864
rect 244148 336824 248788 336852
rect 244148 336812 244154 336824
rect 248782 336812 248788 336824
rect 248840 336812 248846 336864
rect 254486 336812 254492 336864
rect 254544 336852 254550 336864
rect 258258 336852 258264 336864
rect 254544 336824 258264 336852
rect 254544 336812 254550 336824
rect 258258 336812 258264 336824
rect 258316 336812 258322 336864
rect 2958 336744 2964 336796
rect 3016 336784 3022 336796
rect 434898 336784 434904 336796
rect 3016 336756 434904 336784
rect 3016 336744 3022 336756
rect 434898 336744 434904 336756
rect 434956 336744 434962 336796
rect 82722 336676 82728 336728
rect 82780 336716 82786 336728
rect 125962 336716 125968 336728
rect 82780 336688 125968 336716
rect 82780 336676 82786 336688
rect 125962 336676 125968 336688
rect 126020 336676 126026 336728
rect 257706 336676 257712 336728
rect 257764 336716 257770 336728
rect 257798 336716 257804 336728
rect 257764 336688 257804 336716
rect 257764 336676 257770 336688
rect 257798 336676 257804 336688
rect 257856 336676 257862 336728
rect 390922 336716 390928 336728
rect 390883 336688 390928 336716
rect 390922 336676 390928 336688
rect 390980 336676 390986 336728
rect 257709 335291 257767 335297
rect 257709 335257 257721 335291
rect 257755 335288 257767 335291
rect 257798 335288 257804 335300
rect 257755 335260 257804 335288
rect 257755 335257 257767 335260
rect 257709 335251 257767 335257
rect 257798 335248 257804 335260
rect 257856 335248 257862 335300
rect 503530 333276 503536 333328
rect 503588 333316 503594 333328
rect 503806 333316 503812 333328
rect 503588 333288 503812 333316
rect 503588 333276 503594 333288
rect 503806 333276 503812 333288
rect 503864 333276 503870 333328
rect 504358 333276 504364 333328
rect 504416 333316 504422 333328
rect 504818 333316 504824 333328
rect 504416 333288 504824 333316
rect 504416 333276 504422 333288
rect 504818 333276 504824 333288
rect 504876 333276 504882 333328
rect 128909 332367 128967 332373
rect 128909 332333 128921 332367
rect 128955 332364 128967 332367
rect 128998 332364 129004 332376
rect 128955 332336 129004 332364
rect 128955 332333 128967 332336
rect 128909 332327 128967 332333
rect 128998 332324 129004 332336
rect 129056 332324 129062 332376
rect 213917 331347 213975 331353
rect 213917 331313 213929 331347
rect 213963 331344 213975 331347
rect 214006 331344 214012 331356
rect 213963 331316 214012 331344
rect 213963 331313 213975 331316
rect 213917 331307 213975 331313
rect 214006 331304 214012 331316
rect 214064 331304 214070 331356
rect 128722 331276 128728 331288
rect 128683 331248 128728 331276
rect 128722 331236 128728 331248
rect 128780 331236 128786 331288
rect 503622 331168 503628 331220
rect 503680 331208 503686 331220
rect 503990 331208 503996 331220
rect 503680 331180 503996 331208
rect 503680 331168 503686 331180
rect 503990 331168 503996 331180
rect 504048 331168 504054 331220
rect 134242 331100 134248 331152
rect 134300 331100 134306 331152
rect 134260 331016 134288 331100
rect 134242 330964 134248 331016
rect 134300 330964 134306 331016
rect 284110 328556 284116 328568
rect 284071 328528 284116 328556
rect 284110 328516 284116 328528
rect 284168 328516 284174 328568
rect 128722 328488 128728 328500
rect 128683 328460 128728 328488
rect 128722 328448 128728 328460
rect 128780 328448 128786 328500
rect 209774 328448 209780 328500
rect 209832 328488 209838 328500
rect 209958 328488 209964 328500
rect 209832 328460 209964 328488
rect 209832 328448 209838 328460
rect 209958 328448 209964 328460
rect 210016 328448 210022 328500
rect 213914 328488 213920 328500
rect 213875 328460 213920 328488
rect 213914 328448 213920 328460
rect 213972 328448 213978 328500
rect 284021 328423 284079 328429
rect 284021 328389 284033 328423
rect 284067 328420 284079 328423
rect 284110 328420 284116 328432
rect 284067 328392 284116 328420
rect 284067 328389 284079 328392
rect 284021 328383 284079 328389
rect 284110 328380 284116 328392
rect 284168 328380 284174 328432
rect 390922 327128 390928 327140
rect 390883 327100 390928 327128
rect 390922 327088 390928 327100
rect 390980 327088 390986 327140
rect 358538 325660 358544 325712
rect 358596 325700 358602 325712
rect 358722 325700 358728 325712
rect 358596 325672 358728 325700
rect 358596 325660 358602 325672
rect 358722 325660 358728 325672
rect 358780 325660 358786 325712
rect 297634 323660 297640 323672
rect 297595 323632 297640 323660
rect 297634 323620 297640 323632
rect 297692 323620 297698 323672
rect 503898 321716 503904 321768
rect 503956 321756 503962 321768
rect 503956 321728 504001 321756
rect 503956 321716 503962 321728
rect 390833 321691 390891 321697
rect 390833 321657 390845 321691
rect 390879 321688 390891 321691
rect 390922 321688 390928 321700
rect 390879 321660 390928 321688
rect 390879 321657 390891 321660
rect 390833 321651 390891 321657
rect 390922 321648 390928 321660
rect 390980 321648 390986 321700
rect 503990 321688 503996 321700
rect 503951 321660 503996 321688
rect 503990 321648 503996 321660
rect 504048 321648 504054 321700
rect 132770 321580 132776 321632
rect 132828 321620 132834 321632
rect 579614 321620 579620 321632
rect 132828 321592 579620 321620
rect 132828 321580 132834 321592
rect 579614 321580 579620 321592
rect 579672 321580 579678 321632
rect 390830 321552 390836 321564
rect 390791 321524 390836 321552
rect 390830 321512 390836 321524
rect 390888 321512 390894 321564
rect 503898 321552 503904 321564
rect 503859 321524 503904 321552
rect 503898 321512 503904 321524
rect 503956 321512 503962 321564
rect 297634 318900 297640 318912
rect 297595 318872 297640 318900
rect 297634 318860 297640 318872
rect 297692 318860 297698 318912
rect 153378 318792 153384 318844
rect 153436 318832 153442 318844
rect 153470 318832 153476 318844
rect 153436 318804 153476 318832
rect 153436 318792 153442 318804
rect 153470 318792 153476 318804
rect 153528 318792 153534 318844
rect 284018 318832 284024 318844
rect 283979 318804 284024 318832
rect 284018 318792 284024 318804
rect 284076 318792 284082 318844
rect 503990 318832 503996 318844
rect 503951 318804 503996 318832
rect 503990 318792 503996 318804
rect 504048 318792 504054 318844
rect 128630 318724 128636 318776
rect 128688 318764 128694 318776
rect 128722 318764 128728 318776
rect 128688 318736 128728 318764
rect 128688 318724 128694 318736
rect 128722 318724 128728 318736
rect 128780 318724 128786 318776
rect 134153 318767 134211 318773
rect 134153 318733 134165 318767
rect 134199 318764 134211 318767
rect 134242 318764 134248 318776
rect 134199 318736 134248 318764
rect 134199 318733 134211 318736
rect 134153 318727 134211 318733
rect 134242 318724 134248 318736
rect 134300 318724 134306 318776
rect 209774 318764 209780 318776
rect 209735 318736 209780 318764
rect 209774 318724 209780 318736
rect 209832 318724 209838 318776
rect 503714 318764 503720 318776
rect 503675 318736 503720 318764
rect 503714 318724 503720 318736
rect 503772 318724 503778 318776
rect 257706 317472 257712 317484
rect 257667 317444 257712 317472
rect 257706 317432 257712 317444
rect 257764 317432 257770 317484
rect 128630 317404 128636 317416
rect 128591 317376 128636 317404
rect 128630 317364 128636 317376
rect 128688 317364 128694 317416
rect 153378 311924 153384 311976
rect 153436 311964 153442 311976
rect 153470 311964 153476 311976
rect 153436 311936 153476 311964
rect 153436 311924 153442 311936
rect 153470 311924 153476 311936
rect 153528 311924 153534 311976
rect 297542 311924 297548 311976
rect 297600 311924 297606 311976
rect 297560 311828 297588 311924
rect 503622 311856 503628 311908
rect 503680 311896 503686 311908
rect 503990 311896 503996 311908
rect 503680 311868 503996 311896
rect 503680 311856 503686 311868
rect 503990 311856 503996 311868
rect 504048 311856 504054 311908
rect 297634 311828 297640 311840
rect 297560 311800 297640 311828
rect 297634 311788 297640 311800
rect 297692 311788 297698 311840
rect 503622 311720 503628 311772
rect 503680 311760 503686 311772
rect 503990 311760 503996 311772
rect 503680 311732 503996 311760
rect 503680 311720 503686 311732
rect 503990 311720 503996 311732
rect 504048 311720 504054 311772
rect 131850 310496 131856 310548
rect 131908 310536 131914 310548
rect 579706 310536 579712 310548
rect 131908 310508 579712 310536
rect 131908 310496 131914 310508
rect 579706 310496 579712 310508
rect 579764 310496 579770 310548
rect 283926 309204 283932 309256
rect 283984 309244 283990 309256
rect 284110 309244 284116 309256
rect 283984 309216 284116 309244
rect 283984 309204 283990 309216
rect 284110 309204 284116 309216
rect 284168 309204 284174 309256
rect 128633 309179 128691 309185
rect 128633 309145 128645 309179
rect 128679 309176 128691 309179
rect 128722 309176 128728 309188
rect 128679 309148 128728 309176
rect 128679 309145 128691 309148
rect 128633 309139 128691 309145
rect 128722 309136 128728 309148
rect 128780 309136 128786 309188
rect 134150 309176 134156 309188
rect 134111 309148 134156 309176
rect 134150 309136 134156 309148
rect 134208 309136 134214 309188
rect 209774 309176 209780 309188
rect 209735 309148 209780 309176
rect 209774 309136 209780 309148
rect 209832 309136 209838 309188
rect 503717 309179 503775 309185
rect 503717 309145 503729 309179
rect 503763 309176 503775 309179
rect 503806 309176 503812 309188
rect 503763 309148 503812 309176
rect 503763 309145 503775 309148
rect 503717 309139 503775 309145
rect 503806 309136 503812 309148
rect 503864 309136 503870 309188
rect 284021 309111 284079 309117
rect 284021 309077 284033 309111
rect 284067 309108 284079 309111
rect 284110 309108 284116 309120
rect 284067 309080 284116 309108
rect 284067 309077 284079 309080
rect 284021 309071 284079 309077
rect 284110 309068 284116 309080
rect 284168 309068 284174 309120
rect 390833 309111 390891 309117
rect 390833 309077 390845 309111
rect 390879 309108 390891 309111
rect 390922 309108 390928 309120
rect 390879 309080 390928 309108
rect 390879 309077 390891 309080
rect 390833 309071 390891 309077
rect 390922 309068 390928 309080
rect 390980 309068 390986 309120
rect 504358 309108 504364 309120
rect 504319 309080 504364 309108
rect 504358 309068 504364 309080
rect 504416 309068 504422 309120
rect 132678 308252 132684 308304
rect 132736 308292 132742 308304
rect 132862 308292 132868 308304
rect 132736 308264 132868 308292
rect 132736 308252 132742 308264
rect 132862 308252 132868 308264
rect 132920 308252 132926 308304
rect 297818 308048 297824 308100
rect 297876 308048 297882 308100
rect 297836 307828 297864 308048
rect 4062 307776 4068 307828
rect 4120 307816 4126 307828
rect 5258 307816 5264 307828
rect 4120 307788 5264 307816
rect 4120 307776 4126 307788
rect 5258 307776 5264 307788
rect 5316 307776 5322 307828
rect 297818 307776 297824 307828
rect 297876 307776 297882 307828
rect 128722 307748 128728 307760
rect 128683 307720 128728 307748
rect 128722 307708 128728 307720
rect 128780 307708 128786 307760
rect 257798 307748 257804 307760
rect 257759 307720 257804 307748
rect 257798 307708 257804 307720
rect 257856 307708 257862 307760
rect 297545 307751 297603 307757
rect 297545 307717 297557 307751
rect 297591 307748 297603 307751
rect 297634 307748 297640 307760
rect 297591 307720 297640 307748
rect 297591 307717 297603 307720
rect 297545 307711 297603 307717
rect 297634 307708 297640 307720
rect 297692 307708 297698 307760
rect 358538 306348 358544 306400
rect 358596 306388 358602 306400
rect 358722 306388 358728 306400
rect 358596 306360 358728 306388
rect 358596 306348 358602 306360
rect 358722 306348 358728 306360
rect 358780 306348 358786 306400
rect 153286 302200 153292 302252
rect 153344 302240 153350 302252
rect 153470 302240 153476 302252
rect 153344 302212 153476 302240
rect 153344 302200 153350 302212
rect 153470 302200 153476 302212
rect 153528 302200 153534 302252
rect 128722 302172 128728 302184
rect 128683 302144 128728 302172
rect 128722 302132 128728 302144
rect 128780 302132 128786 302184
rect 134150 302132 134156 302184
rect 134208 302172 134214 302184
rect 134334 302172 134340 302184
rect 134208 302144 134340 302172
rect 134208 302132 134214 302144
rect 134334 302132 134340 302144
rect 134392 302132 134398 302184
rect 284018 299588 284024 299600
rect 283979 299560 284024 299588
rect 284018 299548 284024 299560
rect 284076 299548 284082 299600
rect 390830 299520 390836 299532
rect 390791 299492 390836 299520
rect 390830 299480 390836 299492
rect 390888 299480 390894 299532
rect 504361 299523 504419 299529
rect 504361 299489 504373 299523
rect 504407 299520 504419 299523
rect 504450 299520 504456 299532
rect 504407 299492 504456 299520
rect 504407 299489 504419 299492
rect 504361 299483 504419 299489
rect 504450 299480 504456 299492
rect 504508 299480 504514 299532
rect 209774 299452 209780 299464
rect 209735 299424 209780 299452
rect 209774 299412 209780 299424
rect 209832 299412 209838 299464
rect 284018 299452 284024 299464
rect 283979 299424 284024 299452
rect 284018 299412 284024 299424
rect 284076 299412 284082 299464
rect 257801 298163 257859 298169
rect 257801 298129 257813 298163
rect 257847 298160 257859 298163
rect 257890 298160 257896 298172
rect 257847 298132 257896 298160
rect 257847 298129 257859 298132
rect 257801 298123 257859 298129
rect 257890 298120 257896 298132
rect 257948 298120 257954 298172
rect 297542 298160 297548 298172
rect 297503 298132 297548 298160
rect 297542 298120 297548 298132
rect 297600 298120 297606 298172
rect 128722 298092 128728 298104
rect 128683 298064 128728 298092
rect 128722 298052 128728 298064
rect 128780 298052 128786 298104
rect 134245 298095 134303 298101
rect 134245 298061 134257 298095
rect 134291 298092 134303 298095
rect 134334 298092 134340 298104
rect 134291 298064 134340 298092
rect 134291 298061 134303 298064
rect 134245 298055 134303 298061
rect 134334 298052 134340 298064
rect 134392 298052 134398 298104
rect 3326 293972 3332 294024
rect 3384 294012 3390 294024
rect 434530 294012 434536 294024
rect 3384 293984 434536 294012
rect 3384 293972 3390 293984
rect 434530 293972 434536 293984
rect 434588 293972 434594 294024
rect 504266 292544 504272 292596
rect 504324 292584 504330 292596
rect 504450 292584 504456 292596
rect 504324 292556 504456 292584
rect 504324 292544 504330 292556
rect 504450 292544 504456 292556
rect 504508 292544 504514 292596
rect 128722 292448 128728 292460
rect 128683 292420 128728 292448
rect 128722 292408 128728 292420
rect 128780 292408 128786 292460
rect 284021 289935 284079 289941
rect 284021 289901 284033 289935
rect 284067 289932 284079 289935
rect 284110 289932 284116 289944
rect 284067 289904 284116 289932
rect 284067 289901 284079 289904
rect 284021 289895 284079 289901
rect 284110 289892 284116 289904
rect 284168 289892 284174 289944
rect 209774 289864 209780 289876
rect 209735 289836 209780 289864
rect 209774 289824 209780 289836
rect 209832 289824 209838 289876
rect 284021 289799 284079 289805
rect 284021 289765 284033 289799
rect 284067 289796 284079 289799
rect 284110 289796 284116 289808
rect 284067 289768 284116 289796
rect 284067 289765 284079 289768
rect 284021 289759 284079 289765
rect 284110 289756 284116 289768
rect 284168 289756 284174 289808
rect 390833 289799 390891 289805
rect 390833 289765 390845 289799
rect 390879 289796 390891 289799
rect 390922 289796 390928 289808
rect 390879 289768 390928 289796
rect 390879 289765 390891 289768
rect 390833 289759 390891 289765
rect 390922 289756 390928 289768
rect 390980 289756 390986 289808
rect 134242 288436 134248 288448
rect 134203 288408 134248 288436
rect 134242 288396 134248 288408
rect 134300 288396 134306 288448
rect 257798 288396 257804 288448
rect 257856 288436 257862 288448
rect 257890 288436 257896 288448
rect 257856 288408 257896 288436
rect 257856 288396 257862 288408
rect 257890 288396 257896 288408
rect 257948 288396 257954 288448
rect 504266 288436 504272 288448
rect 504227 288408 504272 288436
rect 504266 288396 504272 288408
rect 504324 288396 504330 288448
rect 297545 288371 297603 288377
rect 297545 288337 297557 288371
rect 297591 288368 297603 288371
rect 297634 288368 297640 288380
rect 297591 288340 297640 288368
rect 297591 288337 297603 288340
rect 297545 288331 297603 288337
rect 297634 288328 297640 288340
rect 297692 288328 297698 288380
rect 257798 288300 257804 288312
rect 257759 288272 257804 288300
rect 257798 288260 257804 288272
rect 257856 288260 257862 288312
rect 358538 287036 358544 287088
rect 358596 287076 358602 287088
rect 358722 287076 358728 287088
rect 358596 287048 358728 287076
rect 358596 287036 358602 287048
rect 358722 287036 358728 287048
rect 358780 287036 358786 287088
rect 503714 283024 503720 283076
rect 503772 283064 503778 283076
rect 503772 283036 503852 283064
rect 503772 283024 503778 283036
rect 503824 283008 503852 283036
rect 503806 282956 503812 283008
rect 503864 282956 503870 283008
rect 128630 282928 128636 282940
rect 128591 282900 128636 282928
rect 128630 282888 128636 282900
rect 128688 282888 128694 282940
rect 153286 282888 153292 282940
rect 153344 282928 153350 282940
rect 153470 282928 153476 282940
rect 153344 282900 153476 282928
rect 153344 282888 153350 282900
rect 153470 282888 153476 282900
rect 153528 282888 153534 282940
rect 284018 280276 284024 280288
rect 283979 280248 284024 280276
rect 284018 280236 284024 280248
rect 284076 280236 284082 280288
rect 357250 280236 357256 280288
rect 357308 280276 357314 280288
rect 357342 280276 357348 280288
rect 357308 280248 357348 280276
rect 357308 280236 357314 280248
rect 357342 280236 357348 280248
rect 357400 280236 357406 280288
rect 504269 280279 504327 280285
rect 504269 280245 504281 280279
rect 504315 280276 504327 280279
rect 504450 280276 504456 280288
rect 504315 280248 504456 280276
rect 504315 280245 504327 280248
rect 504269 280239 504327 280245
rect 504450 280236 504456 280248
rect 504508 280236 504514 280288
rect 390830 280208 390836 280220
rect 390791 280180 390836 280208
rect 390830 280168 390836 280180
rect 390888 280168 390894 280220
rect 153378 280140 153384 280152
rect 153339 280112 153384 280140
rect 153378 280100 153384 280112
rect 153436 280100 153442 280152
rect 209774 280140 209780 280152
rect 209735 280112 209780 280140
rect 209774 280100 209780 280112
rect 209832 280100 209838 280152
rect 284018 280140 284024 280152
rect 283979 280112 284024 280140
rect 284018 280100 284024 280112
rect 284076 280100 284082 280152
rect 357250 280140 357256 280152
rect 357211 280112 357256 280140
rect 357250 280100 357256 280112
rect 357308 280100 357314 280152
rect 134150 278808 134156 278860
rect 134208 278848 134214 278860
rect 134242 278848 134248 278860
rect 134208 278820 134248 278848
rect 134208 278808 134214 278820
rect 134242 278808 134248 278820
rect 134300 278808 134306 278860
rect 128630 278780 128636 278792
rect 128591 278752 128636 278780
rect 128630 278740 128636 278752
rect 128688 278740 128694 278792
rect 257801 278783 257859 278789
rect 257801 278749 257813 278783
rect 257847 278780 257859 278783
rect 257890 278780 257896 278792
rect 257847 278752 257896 278780
rect 257847 278749 257859 278752
rect 257801 278743 257859 278749
rect 257890 278740 257896 278752
rect 257948 278740 257954 278792
rect 134242 278712 134248 278724
rect 134203 278684 134248 278712
rect 134242 278672 134248 278684
rect 134300 278672 134306 278724
rect 504450 278712 504456 278724
rect 504411 278684 504456 278712
rect 504450 278672 504456 278684
rect 504508 278672 504514 278724
rect 132678 274660 132684 274712
rect 132736 274700 132742 274712
rect 579614 274700 579620 274712
rect 132736 274672 579620 274700
rect 132736 274660 132742 274672
rect 579614 274660 579620 274672
rect 579672 274660 579678 274712
rect 128630 273340 128636 273352
rect 128591 273312 128636 273340
rect 128630 273300 128636 273312
rect 128688 273300 128694 273352
rect 503622 273300 503628 273352
rect 503680 273340 503686 273352
rect 503990 273340 503996 273352
rect 503680 273312 503996 273340
rect 503680 273300 503686 273312
rect 503990 273300 503996 273312
rect 504048 273300 504054 273352
rect 153381 273275 153439 273281
rect 153381 273241 153393 273275
rect 153427 273272 153439 273275
rect 153562 273272 153568 273284
rect 153427 273244 153568 273272
rect 153427 273241 153439 273244
rect 153381 273235 153439 273241
rect 153562 273232 153568 273244
rect 153620 273232 153626 273284
rect 503622 273164 503628 273216
rect 503680 273204 503686 273216
rect 503990 273204 503996 273216
rect 503680 273176 503996 273204
rect 503680 273164 503686 273176
rect 503990 273164 503996 273176
rect 504048 273164 504054 273216
rect 209774 270552 209780 270564
rect 209735 270524 209780 270552
rect 209774 270512 209780 270524
rect 209832 270512 209838 270564
rect 284018 270552 284024 270564
rect 283979 270524 284024 270552
rect 284018 270512 284024 270524
rect 284076 270512 284082 270564
rect 297545 270555 297603 270561
rect 297545 270521 297557 270555
rect 297591 270552 297603 270555
rect 297634 270552 297640 270564
rect 297591 270524 297640 270552
rect 297591 270521 297603 270524
rect 297545 270515 297603 270521
rect 297634 270512 297640 270524
rect 297692 270512 297698 270564
rect 357253 270555 357311 270561
rect 357253 270521 357265 270555
rect 357299 270552 357311 270555
rect 357342 270552 357348 270564
rect 357299 270524 357348 270552
rect 357299 270521 357311 270524
rect 357253 270515 357311 270521
rect 357342 270512 357348 270524
rect 357400 270512 357406 270564
rect 128630 270484 128636 270496
rect 128591 270456 128636 270484
rect 128630 270444 128636 270456
rect 128688 270444 128694 270496
rect 153562 270484 153568 270496
rect 153523 270456 153568 270484
rect 153562 270444 153568 270456
rect 153620 270444 153626 270496
rect 257798 270484 257804 270496
rect 257759 270456 257804 270484
rect 257798 270444 257804 270456
rect 257856 270444 257862 270496
rect 390922 270484 390928 270496
rect 390883 270456 390928 270484
rect 390922 270444 390928 270456
rect 390980 270444 390986 270496
rect 134242 269124 134248 269136
rect 134203 269096 134248 269124
rect 134242 269084 134248 269096
rect 134300 269084 134306 269136
rect 504453 269127 504511 269133
rect 504453 269093 504465 269127
rect 504499 269124 504511 269127
rect 504634 269124 504640 269136
rect 504499 269096 504640 269124
rect 504499 269093 504511 269096
rect 504453 269087 504511 269093
rect 504634 269084 504640 269096
rect 504692 269084 504698 269136
rect 358538 267724 358544 267776
rect 358596 267764 358602 267776
rect 358722 267764 358728 267776
rect 358596 267736 358728 267764
rect 358596 267724 358602 267736
rect 358722 267724 358728 267736
rect 358780 267724 358786 267776
rect 2774 264936 2780 264988
rect 2832 264976 2838 264988
rect 5442 264976 5448 264988
rect 2832 264948 5448 264976
rect 2832 264936 2838 264948
rect 5442 264936 5448 264948
rect 5500 264936 5506 264988
rect 284018 263684 284024 263696
rect 283979 263656 284024 263684
rect 284018 263644 284024 263656
rect 284076 263644 284082 263696
rect 297542 263684 297548 263696
rect 297503 263656 297548 263684
rect 297542 263644 297548 263656
rect 297600 263644 297606 263696
rect 503714 263644 503720 263696
rect 503772 263684 503778 263696
rect 503990 263684 503996 263696
rect 503772 263656 503996 263684
rect 503772 263644 503778 263656
rect 503990 263644 503996 263656
rect 504048 263644 504054 263696
rect 131574 263576 131580 263628
rect 131632 263616 131638 263628
rect 580166 263616 580172 263628
rect 131632 263588 580172 263616
rect 131632 263576 131638 263588
rect 580166 263576 580172 263588
rect 580224 263576 580230 263628
rect 257798 263548 257804 263560
rect 257759 263520 257804 263548
rect 257798 263508 257804 263520
rect 257856 263508 257862 263560
rect 503714 263508 503720 263560
rect 503772 263548 503778 263560
rect 503990 263548 503996 263560
rect 503772 263520 503996 263548
rect 503772 263508 503778 263520
rect 503990 263508 503996 263520
rect 504048 263508 504054 263560
rect 390922 263480 390928 263492
rect 390883 263452 390928 263480
rect 390922 263440 390928 263452
rect 390980 263440 390986 263492
rect 284018 260964 284024 260976
rect 283979 260936 284024 260964
rect 284018 260924 284024 260936
rect 284076 260924 284082 260976
rect 153565 260899 153623 260905
rect 153565 260865 153577 260899
rect 153611 260896 153623 260899
rect 153654 260896 153660 260908
rect 153611 260868 153660 260896
rect 153611 260865 153623 260868
rect 153565 260859 153623 260865
rect 153654 260856 153660 260868
rect 153712 260856 153718 260908
rect 297542 260896 297548 260908
rect 297503 260868 297548 260896
rect 297542 260856 297548 260868
rect 297600 260856 297606 260908
rect 134245 260831 134303 260837
rect 134245 260797 134257 260831
rect 134291 260828 134303 260831
rect 134334 260828 134340 260840
rect 134291 260800 134340 260828
rect 134291 260797 134303 260800
rect 134245 260791 134303 260797
rect 134334 260788 134340 260800
rect 134392 260788 134398 260840
rect 209774 260828 209780 260840
rect 209735 260800 209780 260828
rect 209774 260788 209780 260800
rect 209832 260788 209838 260840
rect 257798 260828 257804 260840
rect 257759 260800 257804 260828
rect 257798 260788 257804 260800
rect 257856 260788 257862 260840
rect 284018 260788 284024 260840
rect 284076 260828 284082 260840
rect 284294 260828 284300 260840
rect 284076 260800 284300 260828
rect 284076 260788 284082 260800
rect 284294 260788 284300 260800
rect 284352 260788 284358 260840
rect 390922 260828 390928 260840
rect 390883 260800 390928 260828
rect 390922 260788 390928 260800
rect 390980 260788 390986 260840
rect 504266 260828 504272 260840
rect 504227 260800 504272 260828
rect 504266 260788 504272 260800
rect 504324 260788 504330 260840
rect 128633 259403 128691 259409
rect 128633 259369 128645 259403
rect 128679 259400 128691 259403
rect 128722 259400 128728 259412
rect 128679 259372 128728 259400
rect 128679 259369 128691 259372
rect 128633 259363 128691 259369
rect 128722 259360 128728 259372
rect 128780 259360 128786 259412
rect 284110 254600 284116 254652
rect 284168 254640 284174 254652
rect 284294 254640 284300 254652
rect 284168 254612 284300 254640
rect 284168 254600 284174 254612
rect 284294 254600 284300 254612
rect 284352 254600 284358 254652
rect 153654 254028 153660 254040
rect 153580 254000 153660 254028
rect 153580 253904 153608 254000
rect 153654 253988 153660 254000
rect 153712 253988 153718 254040
rect 503622 253988 503628 254040
rect 503680 254028 503686 254040
rect 503990 254028 503996 254040
rect 503680 254000 503996 254028
rect 503680 253988 503686 254000
rect 503990 253988 503996 254000
rect 504048 253988 504054 254040
rect 153562 253852 153568 253904
rect 153620 253852 153626 253904
rect 503622 253852 503628 253904
rect 503680 253892 503686 253904
rect 503990 253892 503996 253904
rect 503680 253864 503996 253892
rect 503680 253852 503686 253864
rect 503990 253852 503996 253864
rect 504048 253852 504054 253904
rect 257798 253824 257804 253836
rect 257759 253796 257804 253824
rect 257798 253784 257804 253796
rect 257856 253784 257862 253836
rect 390922 253824 390928 253836
rect 390883 253796 390928 253824
rect 390922 253784 390928 253796
rect 390980 253784 390986 253836
rect 504266 253824 504272 253836
rect 504227 253796 504272 253824
rect 504266 253784 504272 253796
rect 504324 253784 504330 253836
rect 284202 251404 284208 251456
rect 284260 251404 284266 251456
rect 209774 251308 209780 251320
rect 209735 251280 209780 251308
rect 209774 251268 209780 251280
rect 209832 251268 209838 251320
rect 284220 251252 284248 251404
rect 297358 251268 297364 251320
rect 297416 251308 297422 251320
rect 297634 251308 297640 251320
rect 297416 251280 297640 251308
rect 297416 251268 297422 251280
rect 297634 251268 297640 251280
rect 297692 251268 297698 251320
rect 347792 251280 357296 251308
rect 3326 251200 3332 251252
rect 3384 251240 3390 251252
rect 284113 251243 284171 251249
rect 284113 251240 284125 251243
rect 3384 251212 284125 251240
rect 3384 251200 3390 251212
rect 284113 251209 284125 251212
rect 284159 251209 284171 251243
rect 284113 251203 284171 251209
rect 284202 251200 284208 251252
rect 284260 251200 284266 251252
rect 284389 251243 284447 251249
rect 284389 251209 284401 251243
rect 284435 251240 284447 251243
rect 347792 251240 347820 251280
rect 284435 251212 347820 251240
rect 357268 251240 357296 251280
rect 358372 251280 358676 251308
rect 358372 251240 358400 251280
rect 357268 251212 358400 251240
rect 358648 251240 358676 251280
rect 435082 251240 435088 251252
rect 358648 251212 435088 251240
rect 284435 251209 284447 251212
rect 284389 251203 284447 251209
rect 435082 251200 435088 251212
rect 435140 251200 435146 251252
rect 257709 251175 257767 251181
rect 257709 251141 257721 251175
rect 257755 251172 257767 251175
rect 257798 251172 257804 251184
rect 257755 251144 257804 251172
rect 257755 251141 257767 251144
rect 257709 251135 257767 251141
rect 257798 251132 257804 251144
rect 257856 251132 257862 251184
rect 357158 251132 357164 251184
rect 357216 251172 357222 251184
rect 357342 251172 357348 251184
rect 357216 251144 357348 251172
rect 357216 251132 357222 251144
rect 357342 251132 357348 251144
rect 357400 251132 357406 251184
rect 358446 251132 358452 251184
rect 358504 251172 358510 251184
rect 358630 251172 358636 251184
rect 358504 251144 358636 251172
rect 358504 251132 358510 251144
rect 358630 251132 358636 251144
rect 358688 251132 358694 251184
rect 390922 251172 390928 251184
rect 390883 251144 390928 251172
rect 390922 251132 390928 251144
rect 390980 251132 390986 251184
rect 504266 251172 504272 251184
rect 504227 251144 504272 251172
rect 504266 251132 504272 251144
rect 504324 251132 504330 251184
rect 134242 250628 134248 250640
rect 134203 250600 134248 250628
rect 134242 250588 134248 250600
rect 134300 250588 134306 250640
rect 503714 244400 503720 244452
rect 503772 244440 503778 244452
rect 503772 244412 503852 244440
rect 503772 244400 503778 244412
rect 503824 244384 503852 244412
rect 297634 244332 297640 244384
rect 297692 244332 297698 244384
rect 503806 244332 503812 244384
rect 503864 244332 503870 244384
rect 297652 244248 297680 244332
rect 297634 244196 297640 244248
rect 297692 244196 297698 244248
rect 128630 241584 128636 241596
rect 128591 241556 128636 241584
rect 128630 241544 128636 241556
rect 128688 241544 128694 241596
rect 257706 241516 257712 241528
rect 257667 241488 257712 241516
rect 257706 241476 257712 241488
rect 257764 241476 257770 241528
rect 390925 241519 390983 241525
rect 390925 241485 390937 241519
rect 390971 241516 390983 241519
rect 391014 241516 391020 241528
rect 390971 241488 391020 241516
rect 390971 241485 390983 241488
rect 390925 241479 390983 241485
rect 391014 241476 391020 241488
rect 391072 241476 391078 241528
rect 504269 241519 504327 241525
rect 504269 241485 504281 241519
rect 504315 241516 504327 241519
rect 504450 241516 504456 241528
rect 504315 241488 504456 241516
rect 504315 241485 504327 241488
rect 504269 241479 504327 241485
rect 504450 241476 504456 241488
rect 504508 241476 504514 241528
rect 134058 240116 134064 240168
rect 134116 240156 134122 240168
rect 134334 240156 134340 240168
rect 134116 240128 134340 240156
rect 134116 240116 134122 240128
rect 134334 240116 134340 240128
rect 134392 240116 134398 240168
rect 134245 235331 134303 235337
rect 134245 235297 134257 235331
rect 134291 235328 134303 235331
rect 134334 235328 134340 235340
rect 134291 235300 134340 235328
rect 134291 235297 134303 235300
rect 134245 235291 134303 235297
rect 134334 235288 134340 235300
rect 134392 235288 134398 235340
rect 153286 234676 153292 234728
rect 153344 234676 153350 234728
rect 503622 234676 503628 234728
rect 503680 234716 503686 234728
rect 503990 234716 503996 234728
rect 503680 234688 503996 234716
rect 503680 234676 503686 234688
rect 503990 234676 503996 234688
rect 504048 234676 504054 234728
rect 504450 234716 504456 234728
rect 504376 234688 504456 234716
rect 128722 234648 128728 234660
rect 128648 234620 128728 234648
rect 128648 234592 128676 234620
rect 128722 234608 128728 234620
rect 128780 234608 128786 234660
rect 153304 234592 153332 234676
rect 257706 234608 257712 234660
rect 257764 234608 257770 234660
rect 128630 234540 128636 234592
rect 128688 234540 128694 234592
rect 153286 234540 153292 234592
rect 153344 234540 153350 234592
rect 257724 234512 257752 234608
rect 504376 234592 504404 234688
rect 504450 234676 504456 234688
rect 504508 234676 504514 234728
rect 503622 234540 503628 234592
rect 503680 234580 503686 234592
rect 503990 234580 503996 234592
rect 503680 234552 503996 234580
rect 503680 234540 503686 234552
rect 503990 234540 503996 234552
rect 504048 234540 504054 234592
rect 504358 234540 504364 234592
rect 504416 234540 504422 234592
rect 257798 234512 257804 234524
rect 257724 234484 257804 234512
rect 257798 234472 257804 234484
rect 257856 234472 257862 234524
rect 357158 234472 357164 234524
rect 357216 234512 357222 234524
rect 357342 234512 357348 234524
rect 357216 234484 357348 234512
rect 357216 234472 357222 234484
rect 357342 234472 357348 234484
rect 357400 234472 357406 234524
rect 358446 234472 358452 234524
rect 358504 234512 358510 234524
rect 358630 234512 358636 234524
rect 358504 234484 358636 234512
rect 358504 234472 358510 234484
rect 358630 234472 358636 234484
rect 358688 234472 358694 234524
rect 209774 231820 209780 231872
rect 209832 231860 209838 231872
rect 209958 231860 209964 231872
rect 209832 231832 209964 231860
rect 209832 231820 209838 231832
rect 209958 231820 209964 231832
rect 210016 231820 210022 231872
rect 284110 231820 284116 231872
rect 284168 231860 284174 231872
rect 284294 231860 284300 231872
rect 284168 231832 284300 231860
rect 284168 231820 284174 231832
rect 284294 231820 284300 231832
rect 284352 231820 284358 231872
rect 390830 231820 390836 231872
rect 390888 231860 390894 231872
rect 391014 231860 391020 231872
rect 390888 231832 391020 231860
rect 390888 231820 390894 231832
rect 391014 231820 391020 231832
rect 391072 231820 391078 231872
rect 504358 231792 504364 231804
rect 504319 231764 504364 231792
rect 504358 231752 504364 231764
rect 504416 231752 504422 231804
rect 297358 230460 297364 230512
rect 297416 230500 297422 230512
rect 297450 230500 297456 230512
rect 297416 230472 297456 230500
rect 297416 230460 297422 230472
rect 297450 230460 297456 230472
rect 297508 230460 297514 230512
rect 131298 227740 131304 227792
rect 131356 227780 131362 227792
rect 580166 227780 580172 227792
rect 131356 227752 580172 227780
rect 131356 227740 131362 227752
rect 580166 227740 580172 227752
rect 580224 227740 580230 227792
rect 390554 226992 390560 227044
rect 390612 227032 390618 227044
rect 390830 227032 390836 227044
rect 390612 227004 390836 227032
rect 390612 226992 390618 227004
rect 390830 226992 390836 227004
rect 390888 226992 390894 227044
rect 503714 225088 503720 225140
rect 503772 225128 503778 225140
rect 503772 225100 503852 225128
rect 503772 225088 503778 225100
rect 503824 225072 503852 225100
rect 503806 225020 503812 225072
rect 503864 225020 503870 225072
rect 153194 224992 153200 225004
rect 153155 224964 153200 224992
rect 153194 224952 153200 224964
rect 153252 224952 153258 225004
rect 257706 224992 257712 225004
rect 257667 224964 257712 224992
rect 257706 224952 257712 224964
rect 257764 224952 257770 225004
rect 2958 222164 2964 222216
rect 3016 222204 3022 222216
rect 14458 222204 14464 222216
rect 3016 222176 14464 222204
rect 3016 222164 3022 222176
rect 14458 222164 14464 222176
rect 14516 222164 14522 222216
rect 134242 222204 134248 222216
rect 134203 222176 134248 222204
rect 134242 222164 134248 222176
rect 134300 222164 134306 222216
rect 153194 222204 153200 222216
rect 153155 222176 153200 222204
rect 153194 222164 153200 222176
rect 153252 222164 153258 222216
rect 257706 222204 257712 222216
rect 257667 222176 257712 222204
rect 257706 222164 257712 222176
rect 257764 222164 257770 222216
rect 297358 222164 297364 222216
rect 297416 222204 297422 222216
rect 297450 222204 297456 222216
rect 297416 222176 297456 222204
rect 297416 222164 297422 222176
rect 297450 222164 297456 222176
rect 297508 222164 297514 222216
rect 504361 222207 504419 222213
rect 504361 222173 504373 222207
rect 504407 222204 504419 222207
rect 504450 222204 504456 222216
rect 504407 222176 504456 222204
rect 504407 222173 504419 222176
rect 504361 222167 504419 222173
rect 504450 222164 504456 222176
rect 504508 222164 504514 222216
rect 364518 222136 364524 222148
rect 364479 222108 364524 222136
rect 364518 222096 364524 222108
rect 364576 222096 364582 222148
rect 390554 219376 390560 219428
rect 390612 219416 390618 219428
rect 390738 219416 390744 219428
rect 390612 219388 390744 219416
rect 390612 219376 390618 219388
rect 390738 219376 390744 219388
rect 390796 219376 390802 219428
rect 131482 216656 131488 216708
rect 131540 216696 131546 216708
rect 579614 216696 579620 216708
rect 131540 216668 579620 216696
rect 131540 216656 131546 216668
rect 579614 216656 579620 216668
rect 579672 216656 579678 216708
rect 283926 215364 283932 215416
rect 283984 215364 283990 215416
rect 503622 215364 503628 215416
rect 503680 215404 503686 215416
rect 503990 215404 503996 215416
rect 503680 215376 503996 215404
rect 503680 215364 503686 215376
rect 503990 215364 503996 215376
rect 504048 215364 504054 215416
rect 504450 215404 504456 215416
rect 504284 215376 504456 215404
rect 153194 215296 153200 215348
rect 153252 215296 153258 215348
rect 257706 215296 257712 215348
rect 257764 215296 257770 215348
rect 153212 215200 153240 215296
rect 153286 215200 153292 215212
rect 153212 215172 153292 215200
rect 153286 215160 153292 215172
rect 153344 215160 153350 215212
rect 257724 215200 257752 215296
rect 283944 215280 283972 215364
rect 504284 215280 504312 215376
rect 504450 215364 504456 215376
rect 504508 215364 504514 215416
rect 283926 215228 283932 215280
rect 283984 215228 283990 215280
rect 308858 215228 308864 215280
rect 308916 215268 308922 215280
rect 309042 215268 309048 215280
rect 308916 215240 309048 215268
rect 308916 215228 308922 215240
rect 309042 215228 309048 215240
rect 309100 215228 309106 215280
rect 503622 215228 503628 215280
rect 503680 215268 503686 215280
rect 503990 215268 503996 215280
rect 503680 215240 503996 215268
rect 503680 215228 503686 215240
rect 503990 215228 503996 215240
rect 504048 215228 504054 215280
rect 504266 215228 504272 215280
rect 504324 215228 504330 215280
rect 257798 215200 257804 215212
rect 257724 215172 257804 215200
rect 257798 215160 257804 215172
rect 257856 215160 257862 215212
rect 209774 212508 209780 212560
rect 209832 212548 209838 212560
rect 209958 212548 209964 212560
rect 209832 212520 209964 212548
rect 209832 212508 209838 212520
rect 209958 212508 209964 212520
rect 210016 212508 210022 212560
rect 297358 212508 297364 212560
rect 297416 212548 297422 212560
rect 297634 212548 297640 212560
rect 297416 212520 297640 212548
rect 297416 212508 297422 212520
rect 297634 212508 297640 212520
rect 297692 212508 297698 212560
rect 357158 212508 357164 212560
rect 357216 212548 357222 212560
rect 357250 212548 357256 212560
rect 357216 212520 357256 212548
rect 357216 212508 357222 212520
rect 357250 212508 357256 212520
rect 357308 212508 357314 212560
rect 364521 212551 364579 212557
rect 364521 212517 364533 212551
rect 364567 212548 364579 212551
rect 364702 212548 364708 212560
rect 364567 212520 364708 212548
rect 364567 212517 364579 212520
rect 364521 212511 364579 212517
rect 364702 212508 364708 212520
rect 364760 212508 364766 212560
rect 153286 212480 153292 212492
rect 153247 212452 153292 212480
rect 153286 212440 153292 212452
rect 153344 212440 153350 212492
rect 298554 210400 298560 210452
rect 298612 210440 298618 210452
rect 299014 210440 299020 210452
rect 298612 210412 299020 210440
rect 298612 210400 298618 210412
rect 299014 210400 299020 210412
rect 299072 210400 299078 210452
rect 297542 210264 297548 210316
rect 297600 210304 297606 210316
rect 298002 210304 298008 210316
rect 297600 210276 298008 210304
rect 297600 210264 297606 210276
rect 298002 210264 298008 210276
rect 298060 210264 298066 210316
rect 390554 209788 390560 209840
rect 390612 209828 390618 209840
rect 390738 209828 390744 209840
rect 390612 209800 390744 209828
rect 390612 209788 390618 209800
rect 390738 209788 390744 209800
rect 390796 209788 390802 209840
rect 243998 209720 244004 209772
rect 244056 209760 244062 209772
rect 244182 209760 244188 209772
rect 244056 209732 244188 209760
rect 244056 209720 244062 209732
rect 244182 209720 244188 209732
rect 244240 209720 244246 209772
rect 301866 208496 301872 208548
rect 301924 208536 301930 208548
rect 302142 208536 302148 208548
rect 301924 208508 302148 208536
rect 301924 208496 301930 208508
rect 302142 208496 302148 208508
rect 302200 208496 302206 208548
rect 2958 207000 2964 207052
rect 3016 207040 3022 207052
rect 435174 207040 435180 207052
rect 3016 207012 435180 207040
rect 3016 207000 3022 207012
rect 435174 207000 435180 207012
rect 435232 207000 435238 207052
rect 503714 205776 503720 205828
rect 503772 205816 503778 205828
rect 503772 205788 503852 205816
rect 503772 205776 503778 205788
rect 503824 205760 503852 205788
rect 503806 205708 503812 205760
rect 503864 205708 503870 205760
rect 257706 205680 257712 205692
rect 257667 205652 257712 205680
rect 257706 205640 257712 205652
rect 257764 205640 257770 205692
rect 503714 205640 503720 205692
rect 503772 205680 503778 205692
rect 503990 205680 503996 205692
rect 503772 205652 503996 205680
rect 503772 205640 503778 205652
rect 503990 205640 503996 205652
rect 504048 205640 504054 205692
rect 504174 205680 504180 205692
rect 504135 205652 504180 205680
rect 504174 205640 504180 205652
rect 504232 205640 504238 205692
rect 196710 205300 196716 205352
rect 196768 205340 196774 205352
rect 226886 205340 226892 205352
rect 196768 205312 226892 205340
rect 196768 205300 196774 205312
rect 226886 205300 226892 205312
rect 226944 205300 226950 205352
rect 196618 205232 196624 205284
rect 196676 205272 196682 205284
rect 227898 205272 227904 205284
rect 196676 205244 227904 205272
rect 196676 205232 196682 205244
rect 227898 205232 227904 205244
rect 227956 205232 227962 205284
rect 195882 205164 195888 205216
rect 195940 205204 195946 205216
rect 228634 205204 228640 205216
rect 195940 205176 228640 205204
rect 195940 205164 195946 205176
rect 228634 205164 228640 205176
rect 228692 205164 228698 205216
rect 195606 205096 195612 205148
rect 195664 205136 195670 205148
rect 229554 205136 229560 205148
rect 195664 205108 229560 205136
rect 195664 205096 195670 205108
rect 229554 205096 229560 205108
rect 229612 205096 229618 205148
rect 195790 205028 195796 205080
rect 195848 205068 195854 205080
rect 230474 205068 230480 205080
rect 195848 205040 230480 205068
rect 195848 205028 195854 205040
rect 230474 205028 230480 205040
rect 230532 205028 230538 205080
rect 195514 204960 195520 205012
rect 195572 205000 195578 205012
rect 231210 205000 231216 205012
rect 195572 204972 231216 205000
rect 195572 204960 195578 204972
rect 231210 204960 231216 204972
rect 231268 204960 231274 205012
rect 195698 204892 195704 204944
rect 195756 204932 195762 204944
rect 233234 204932 233240 204944
rect 195756 204904 233240 204932
rect 195756 204892 195762 204904
rect 233234 204892 233240 204904
rect 233292 204892 233298 204944
rect 266354 204892 266360 204944
rect 266412 204932 266418 204944
rect 267458 204932 267464 204944
rect 266412 204904 267464 204932
rect 266412 204892 266418 204904
rect 267458 204892 267464 204904
rect 267516 204892 267522 204944
rect 255774 204144 255780 204196
rect 255832 204184 255838 204196
rect 268286 204184 268292 204196
rect 255832 204156 268292 204184
rect 255832 204144 255838 204156
rect 268286 204144 268292 204156
rect 268344 204144 268350 204196
rect 253566 204076 253572 204128
rect 253624 204116 253630 204128
rect 269022 204116 269028 204128
rect 253624 204088 269028 204116
rect 253624 204076 253630 204088
rect 269022 204076 269028 204088
rect 269080 204076 269086 204128
rect 250530 204008 250536 204060
rect 250588 204048 250594 204060
rect 268010 204048 268016 204060
rect 250588 204020 268016 204048
rect 250588 204008 250594 204020
rect 268010 204008 268016 204020
rect 268068 204008 268074 204060
rect 199010 203940 199016 203992
rect 199068 203980 199074 203992
rect 238754 203980 238760 203992
rect 199068 203952 238760 203980
rect 199068 203940 199074 203952
rect 238754 203940 238760 203952
rect 238812 203940 238818 203992
rect 247586 203940 247592 203992
rect 247644 203980 247650 203992
rect 268194 203980 268200 203992
rect 247644 203952 268200 203980
rect 247644 203940 247650 203952
rect 268194 203940 268200 203952
rect 268252 203940 268258 203992
rect 197722 203872 197728 203924
rect 197780 203912 197786 203924
rect 257154 203912 257160 203924
rect 197780 203884 257160 203912
rect 197780 203872 197786 203884
rect 257154 203872 257160 203884
rect 257212 203872 257218 203924
rect 197998 203804 198004 203856
rect 198056 203844 198062 203856
rect 260374 203844 260380 203856
rect 198056 203816 260380 203844
rect 198056 203804 198062 203816
rect 260374 203804 260380 203816
rect 260432 203804 260438 203856
rect 198458 203736 198464 203788
rect 198516 203776 198522 203788
rect 262766 203776 262772 203788
rect 198516 203748 262772 203776
rect 198516 203736 198522 203748
rect 262766 203736 262772 203748
rect 262824 203736 262830 203788
rect 197446 203668 197452 203720
rect 197504 203708 197510 203720
rect 262950 203708 262956 203720
rect 197504 203680 262956 203708
rect 197504 203668 197510 203680
rect 262950 203668 262956 203680
rect 263008 203668 263014 203720
rect 197814 203600 197820 203652
rect 197872 203640 197878 203652
rect 265250 203640 265256 203652
rect 197872 203612 265256 203640
rect 197872 203600 197878 203612
rect 265250 203600 265256 203612
rect 265308 203600 265314 203652
rect 198366 203532 198372 203584
rect 198424 203572 198430 203584
rect 267366 203572 267372 203584
rect 198424 203544 267372 203572
rect 198424 203532 198430 203544
rect 267366 203532 267372 203544
rect 267424 203532 267430 203584
rect 153289 202895 153347 202901
rect 153289 202861 153301 202895
rect 153335 202892 153347 202895
rect 153378 202892 153384 202904
rect 153335 202864 153384 202892
rect 153335 202861 153347 202864
rect 153289 202855 153347 202861
rect 153378 202852 153384 202864
rect 153436 202852 153442 202904
rect 257706 202892 257712 202904
rect 239600 202864 240272 202892
rect 257667 202864 257712 202892
rect 199930 202784 199936 202836
rect 199988 202824 199994 202836
rect 239600 202824 239628 202864
rect 199988 202796 239628 202824
rect 199988 202784 199994 202796
rect 239674 202784 239680 202836
rect 239732 202824 239738 202836
rect 240134 202824 240140 202836
rect 239732 202796 240140 202824
rect 239732 202784 239738 202796
rect 240134 202784 240140 202796
rect 240192 202784 240198 202836
rect 196894 202716 196900 202768
rect 196952 202756 196958 202768
rect 196952 202728 239076 202756
rect 196952 202716 196958 202728
rect 200022 202648 200028 202700
rect 200080 202688 200086 202700
rect 238941 202691 238999 202697
rect 238941 202688 238953 202691
rect 200080 202660 238953 202688
rect 200080 202648 200086 202660
rect 238941 202657 238953 202660
rect 238987 202657 238999 202691
rect 239048 202688 239076 202728
rect 239214 202716 239220 202768
rect 239272 202756 239278 202768
rect 240042 202756 240048 202768
rect 239272 202728 240048 202756
rect 239272 202716 239278 202728
rect 240042 202716 240048 202728
rect 240100 202716 240106 202768
rect 240244 202756 240272 202864
rect 257706 202852 257712 202864
rect 257764 202852 257770 202904
rect 283650 202852 283656 202904
rect 283708 202892 283714 202904
rect 283742 202892 283748 202904
rect 283708 202864 283748 202892
rect 283708 202852 283714 202864
rect 283742 202852 283748 202864
rect 283800 202852 283806 202904
rect 297450 202852 297456 202904
rect 297508 202892 297514 202904
rect 297634 202892 297640 202904
rect 297508 202864 297640 202892
rect 297508 202852 297514 202864
rect 297634 202852 297640 202864
rect 297692 202852 297698 202904
rect 504174 202892 504180 202904
rect 504135 202864 504180 202892
rect 504174 202852 504180 202864
rect 504232 202852 504238 202904
rect 240502 202784 240508 202836
rect 240560 202824 240566 202836
rect 241422 202824 241428 202836
rect 240560 202796 241428 202824
rect 240560 202784 240566 202796
rect 241422 202784 241428 202796
rect 241480 202784 241486 202836
rect 267918 202824 267924 202836
rect 258644 202796 267924 202824
rect 240244 202728 241652 202756
rect 241514 202688 241520 202700
rect 239048 202660 241520 202688
rect 238941 202651 238999 202657
rect 241514 202648 241520 202660
rect 241572 202648 241578 202700
rect 241624 202688 241652 202728
rect 242066 202716 242072 202768
rect 242124 202756 242130 202768
rect 247678 202756 247684 202768
rect 242124 202728 247684 202756
rect 242124 202716 242130 202728
rect 247678 202716 247684 202728
rect 247736 202716 247742 202768
rect 251818 202716 251824 202768
rect 251876 202756 251882 202768
rect 258644 202756 258672 202796
rect 267918 202784 267924 202796
rect 267976 202784 267982 202836
rect 270954 202784 270960 202836
rect 271012 202824 271018 202836
rect 271782 202824 271788 202836
rect 271012 202796 271788 202824
rect 271012 202784 271018 202796
rect 271782 202784 271788 202796
rect 271840 202784 271846 202836
rect 272242 202784 272248 202836
rect 272300 202824 272306 202836
rect 273162 202824 273168 202836
rect 272300 202796 273168 202824
rect 272300 202784 272306 202796
rect 273162 202784 273168 202796
rect 273220 202784 273226 202836
rect 273990 202784 273996 202836
rect 274048 202824 274054 202836
rect 274542 202824 274548 202836
rect 274048 202796 274548 202824
rect 274048 202784 274054 202796
rect 274542 202784 274548 202796
rect 274600 202784 274606 202836
rect 277026 202784 277032 202836
rect 277084 202824 277090 202836
rect 277302 202824 277308 202836
rect 277084 202796 277308 202824
rect 277084 202784 277090 202796
rect 277302 202784 277308 202796
rect 277360 202784 277366 202836
rect 278682 202784 278688 202836
rect 278740 202824 278746 202836
rect 279418 202824 279424 202836
rect 278740 202796 279424 202824
rect 278740 202784 278746 202796
rect 279418 202784 279424 202796
rect 279476 202784 279482 202836
rect 280522 202784 280528 202836
rect 280580 202824 280586 202836
rect 281350 202824 281356 202836
rect 280580 202796 281356 202824
rect 280580 202784 280586 202796
rect 281350 202784 281356 202796
rect 281408 202784 281414 202836
rect 298646 202784 298652 202836
rect 298704 202824 298710 202836
rect 299106 202824 299112 202836
rect 298704 202796 299112 202824
rect 298704 202784 298710 202796
rect 299106 202784 299112 202796
rect 299164 202784 299170 202836
rect 300118 202784 300124 202836
rect 300176 202824 300182 202836
rect 300762 202824 300768 202836
rect 300176 202796 300768 202824
rect 300176 202784 300182 202796
rect 300762 202784 300768 202796
rect 300820 202784 300826 202836
rect 301406 202784 301412 202836
rect 301464 202824 301470 202836
rect 302050 202824 302056 202836
rect 301464 202796 302056 202824
rect 301464 202784 301470 202796
rect 302050 202784 302056 202796
rect 302108 202784 302114 202836
rect 309134 202784 309140 202836
rect 309192 202824 309198 202836
rect 309594 202824 309600 202836
rect 309192 202796 309600 202824
rect 309192 202784 309198 202796
rect 309594 202784 309600 202796
rect 309652 202784 309658 202836
rect 311894 202784 311900 202836
rect 311952 202824 311958 202836
rect 312538 202824 312544 202836
rect 311952 202796 312544 202824
rect 311952 202784 311958 202796
rect 312538 202784 312544 202796
rect 312596 202784 312602 202836
rect 313550 202784 313556 202836
rect 313608 202824 313614 202836
rect 314562 202824 314568 202836
rect 313608 202796 314568 202824
rect 313608 202784 313614 202796
rect 314562 202784 314568 202796
rect 314620 202784 314626 202836
rect 314746 202784 314752 202836
rect 314804 202824 314810 202836
rect 315574 202824 315580 202836
rect 314804 202796 315580 202824
rect 314804 202784 314810 202796
rect 315574 202784 315580 202796
rect 315632 202784 315638 202836
rect 316678 202784 316684 202836
rect 316736 202824 316742 202836
rect 321646 202824 321652 202836
rect 316736 202796 321652 202824
rect 316736 202784 316742 202796
rect 321646 202784 321652 202796
rect 321704 202784 321710 202836
rect 341334 202784 341340 202836
rect 341392 202824 341398 202836
rect 342162 202824 342168 202836
rect 341392 202796 342168 202824
rect 341392 202784 341398 202796
rect 342162 202784 342168 202796
rect 342220 202784 342226 202836
rect 363414 202824 363420 202836
rect 361316 202796 363420 202824
rect 251876 202728 258672 202756
rect 251876 202716 251882 202728
rect 258718 202716 258724 202768
rect 258776 202756 258782 202768
rect 263870 202756 263876 202768
rect 258776 202728 263876 202756
rect 258776 202716 258782 202728
rect 263870 202716 263876 202728
rect 263928 202716 263934 202768
rect 266354 202716 266360 202768
rect 266412 202756 266418 202768
rect 267182 202756 267188 202768
rect 266412 202728 267188 202756
rect 266412 202716 266418 202728
rect 267182 202716 267188 202728
rect 267240 202716 267246 202768
rect 271414 202716 271420 202768
rect 271472 202756 271478 202768
rect 272518 202756 272524 202768
rect 271472 202728 272524 202756
rect 271472 202716 271478 202728
rect 272518 202716 272524 202728
rect 272576 202716 272582 202768
rect 279234 202716 279240 202768
rect 279292 202756 279298 202768
rect 280062 202756 280068 202768
rect 279292 202728 280068 202756
rect 279292 202716 279298 202728
rect 280062 202716 280068 202728
rect 280120 202716 280126 202768
rect 282270 202716 282276 202768
rect 282328 202756 282334 202768
rect 284938 202756 284944 202768
rect 282328 202728 284944 202756
rect 282328 202716 282334 202728
rect 284938 202716 284944 202728
rect 284996 202716 285002 202768
rect 297910 202716 297916 202768
rect 297968 202756 297974 202768
rect 298830 202756 298836 202768
rect 297968 202728 298836 202756
rect 297968 202716 297974 202728
rect 298830 202716 298836 202728
rect 298888 202716 298894 202768
rect 299474 202716 299480 202768
rect 299532 202756 299538 202768
rect 313642 202756 313648 202768
rect 299532 202728 313648 202756
rect 299532 202716 299538 202728
rect 313642 202716 313648 202728
rect 313700 202716 313706 202768
rect 318610 202716 318616 202768
rect 318668 202756 318674 202768
rect 333238 202756 333244 202768
rect 318668 202728 333244 202756
rect 318668 202716 318674 202728
rect 333238 202716 333244 202728
rect 333296 202716 333302 202768
rect 245194 202688 245200 202700
rect 241624 202660 245200 202688
rect 245194 202648 245200 202660
rect 245252 202648 245258 202700
rect 250898 202648 250904 202700
rect 250956 202688 250962 202700
rect 258629 202691 258687 202697
rect 258629 202688 258641 202691
rect 250956 202660 258641 202688
rect 250956 202648 250962 202660
rect 258629 202657 258641 202660
rect 258675 202657 258687 202691
rect 258629 202651 258687 202657
rect 258813 202691 258871 202697
rect 258813 202657 258825 202691
rect 258859 202688 258871 202691
rect 268378 202688 268384 202700
rect 258859 202660 268384 202688
rect 258859 202657 258871 202660
rect 258813 202651 258871 202657
rect 268378 202648 268384 202660
rect 268436 202648 268442 202700
rect 299198 202648 299204 202700
rect 299256 202688 299262 202700
rect 304350 202688 304356 202700
rect 299256 202660 304356 202688
rect 299256 202648 299262 202660
rect 304350 202648 304356 202660
rect 304408 202648 304414 202700
rect 304902 202648 304908 202700
rect 304960 202688 304966 202700
rect 309134 202688 309140 202700
rect 304960 202660 309140 202688
rect 304960 202648 304966 202660
rect 309134 202648 309140 202660
rect 309192 202648 309198 202700
rect 311158 202648 311164 202700
rect 311216 202688 311222 202700
rect 330478 202688 330484 202700
rect 311216 202660 330484 202688
rect 311216 202648 311222 202660
rect 330478 202648 330484 202660
rect 330536 202648 330542 202700
rect 358722 202648 358728 202700
rect 358780 202688 358786 202700
rect 361316 202688 361344 202796
rect 363414 202784 363420 202796
rect 363472 202784 363478 202836
rect 375742 202784 375748 202836
rect 375800 202824 375806 202836
rect 391198 202824 391204 202836
rect 375800 202796 391204 202824
rect 375800 202784 375806 202796
rect 391198 202784 391204 202796
rect 391256 202784 391262 202836
rect 400582 202784 400588 202836
rect 400640 202824 400646 202836
rect 401410 202824 401416 202836
rect 400640 202796 401416 202824
rect 400640 202784 400646 202796
rect 401410 202784 401416 202796
rect 401468 202784 401474 202836
rect 413186 202784 413192 202836
rect 413244 202824 413250 202836
rect 413922 202824 413928 202836
rect 413244 202796 413928 202824
rect 413244 202784 413250 202796
rect 413922 202784 413928 202796
rect 413980 202784 413986 202836
rect 415762 202784 415768 202836
rect 415820 202824 415826 202836
rect 416590 202824 416596 202836
rect 415820 202796 416596 202824
rect 415820 202784 415826 202796
rect 416590 202784 416596 202796
rect 416648 202784 416654 202836
rect 417510 202784 417516 202836
rect 417568 202824 417574 202836
rect 418062 202824 418068 202836
rect 417568 202796 418068 202824
rect 417568 202784 417574 202796
rect 418062 202784 418068 202796
rect 418120 202784 418126 202836
rect 374454 202716 374460 202768
rect 374512 202756 374518 202768
rect 391290 202756 391296 202768
rect 374512 202728 391296 202756
rect 374512 202716 374518 202728
rect 391290 202716 391296 202728
rect 391348 202716 391354 202768
rect 504174 202716 504180 202768
rect 504232 202756 504238 202768
rect 504450 202756 504456 202768
rect 504232 202728 504456 202756
rect 504232 202716 504238 202728
rect 504450 202716 504456 202728
rect 504508 202716 504514 202768
rect 358780 202660 361344 202688
rect 358780 202648 358786 202660
rect 361390 202648 361396 202700
rect 361448 202688 361454 202700
rect 362218 202688 362224 202700
rect 361448 202660 362224 202688
rect 361448 202648 361454 202660
rect 362218 202648 362224 202660
rect 362276 202648 362282 202700
rect 376478 202648 376484 202700
rect 376536 202688 376542 202700
rect 398098 202688 398104 202700
rect 376536 202660 398104 202688
rect 376536 202648 376542 202660
rect 398098 202648 398104 202660
rect 398156 202648 398162 202700
rect 160738 202580 160744 202632
rect 160796 202620 160802 202632
rect 169110 202620 169116 202632
rect 160796 202592 169116 202620
rect 160796 202580 160802 202592
rect 169110 202580 169116 202592
rect 169168 202580 169174 202632
rect 197630 202580 197636 202632
rect 197688 202620 197694 202632
rect 197688 202592 240180 202620
rect 197688 202580 197694 202592
rect 157978 202512 157984 202564
rect 158036 202552 158042 202564
rect 176930 202552 176936 202564
rect 158036 202524 176936 202552
rect 158036 202512 158042 202524
rect 176930 202512 176936 202524
rect 176988 202512 176994 202564
rect 197538 202512 197544 202564
rect 197596 202552 197602 202564
rect 240045 202555 240103 202561
rect 240045 202552 240057 202555
rect 197596 202524 240057 202552
rect 197596 202512 197602 202524
rect 240045 202521 240057 202524
rect 240091 202521 240103 202555
rect 240152 202552 240180 202592
rect 244642 202580 244648 202632
rect 244700 202620 244706 202632
rect 268102 202620 268108 202632
rect 244700 202592 268108 202620
rect 244700 202580 244706 202592
rect 268102 202580 268108 202592
rect 268160 202580 268166 202632
rect 299382 202580 299388 202632
rect 299440 202620 299446 202632
rect 320634 202620 320640 202632
rect 299440 202592 320640 202620
rect 299440 202580 299446 202592
rect 320634 202580 320640 202592
rect 320692 202580 320698 202632
rect 359642 202580 359648 202632
rect 359700 202620 359706 202632
rect 360102 202620 360108 202632
rect 359700 202592 360108 202620
rect 359700 202580 359706 202592
rect 360102 202580 360108 202592
rect 360160 202580 360166 202632
rect 360562 202580 360568 202632
rect 360620 202620 360626 202632
rect 361482 202620 361488 202632
rect 360620 202592 361488 202620
rect 360620 202580 360626 202592
rect 361482 202580 361488 202592
rect 361540 202580 361546 202632
rect 362310 202580 362316 202632
rect 362368 202620 362374 202632
rect 362862 202620 362868 202632
rect 362368 202592 362868 202620
rect 362368 202580 362374 202592
rect 362862 202580 362868 202592
rect 362920 202580 362926 202632
rect 363598 202580 363604 202632
rect 363656 202620 363662 202632
rect 364334 202620 364340 202632
rect 363656 202592 364340 202620
rect 363656 202580 363662 202592
rect 364334 202580 364340 202592
rect 364392 202580 364398 202632
rect 367002 202580 367008 202632
rect 367060 202620 367066 202632
rect 395338 202620 395344 202632
rect 367060 202592 395344 202620
rect 367060 202580 367066 202592
rect 395338 202580 395344 202592
rect 395396 202580 395402 202632
rect 244734 202552 244740 202564
rect 240152 202524 244740 202552
rect 240045 202515 240103 202521
rect 244734 202512 244740 202524
rect 244792 202512 244798 202564
rect 247494 202512 247500 202564
rect 247552 202552 247558 202564
rect 267826 202552 267832 202564
rect 247552 202524 267832 202552
rect 247552 202512 247558 202524
rect 267826 202512 267832 202524
rect 267884 202512 267890 202564
rect 298922 202512 298928 202564
rect 298980 202552 298986 202564
rect 303062 202552 303068 202564
rect 298980 202524 303068 202552
rect 298980 202512 298986 202524
rect 303062 202512 303068 202524
rect 303120 202512 303126 202564
rect 303154 202512 303160 202564
rect 303212 202552 303218 202564
rect 304258 202552 304264 202564
rect 303212 202524 304264 202552
rect 303212 202512 303218 202524
rect 304258 202512 304264 202524
rect 304316 202512 304322 202564
rect 306650 202512 306656 202564
rect 306708 202552 306714 202564
rect 307662 202552 307668 202564
rect 306708 202524 307668 202552
rect 306708 202512 306714 202524
rect 307662 202512 307668 202524
rect 307720 202512 307726 202564
rect 307757 202555 307815 202561
rect 307757 202521 307769 202555
rect 307803 202552 307815 202555
rect 325694 202552 325700 202564
rect 307803 202524 325700 202552
rect 307803 202521 307815 202524
rect 307757 202515 307815 202521
rect 325694 202512 325700 202524
rect 325752 202512 325758 202564
rect 346670 202512 346676 202564
rect 346728 202552 346734 202564
rect 351178 202552 351184 202564
rect 346728 202524 351184 202552
rect 346728 202512 346734 202524
rect 351178 202512 351184 202524
rect 351236 202512 351242 202564
rect 357894 202512 357900 202564
rect 357952 202552 357958 202564
rect 393314 202552 393320 202564
rect 357952 202524 393320 202552
rect 357952 202512 357958 202524
rect 393314 202512 393320 202524
rect 393372 202512 393378 202564
rect 159358 202444 159364 202496
rect 159416 202484 159422 202496
rect 178034 202484 178040 202496
rect 159416 202456 178040 202484
rect 159416 202444 159422 202456
rect 178034 202444 178040 202456
rect 178092 202444 178098 202496
rect 197354 202444 197360 202496
rect 197412 202484 197418 202496
rect 251910 202484 251916 202496
rect 197412 202456 251916 202484
rect 197412 202444 197418 202456
rect 251910 202444 251916 202456
rect 251968 202444 251974 202496
rect 252462 202444 252468 202496
rect 252520 202484 252526 202496
rect 268470 202484 268476 202496
rect 252520 202456 268476 202484
rect 252520 202444 252526 202456
rect 268470 202444 268476 202456
rect 268528 202444 268534 202496
rect 286226 202444 286232 202496
rect 286284 202484 286290 202496
rect 286870 202484 286876 202496
rect 286284 202456 286876 202484
rect 286284 202444 286290 202456
rect 286870 202444 286876 202456
rect 286928 202444 286934 202496
rect 287514 202444 287520 202496
rect 287572 202484 287578 202496
rect 288250 202484 288256 202496
rect 287572 202456 288256 202484
rect 287572 202444 287578 202456
rect 288250 202444 288256 202456
rect 288308 202444 288314 202496
rect 289446 202444 289452 202496
rect 289504 202484 289510 202496
rect 289722 202484 289728 202496
rect 289504 202456 289728 202484
rect 289504 202444 289510 202456
rect 289722 202444 289728 202456
rect 289780 202444 289786 202496
rect 290550 202444 290556 202496
rect 290608 202484 290614 202496
rect 291010 202484 291016 202496
rect 290608 202456 291016 202484
rect 290608 202444 290614 202456
rect 291010 202444 291016 202456
rect 291068 202444 291074 202496
rect 292206 202444 292212 202496
rect 292264 202484 292270 202496
rect 292390 202484 292396 202496
rect 292264 202456 292396 202484
rect 292264 202444 292270 202456
rect 292390 202444 292396 202456
rect 292448 202444 292454 202496
rect 298738 202484 298744 202496
rect 292500 202456 298744 202484
rect 153838 202376 153844 202428
rect 153896 202416 153902 202428
rect 182174 202416 182180 202428
rect 153896 202388 182180 202416
rect 153896 202376 153902 202388
rect 182174 202376 182180 202388
rect 182232 202376 182238 202428
rect 199194 202376 199200 202428
rect 199252 202416 199258 202428
rect 254026 202416 254032 202428
rect 199252 202388 254032 202416
rect 199252 202376 199258 202388
rect 254026 202376 254032 202388
rect 254084 202376 254090 202428
rect 255958 202376 255964 202428
rect 256016 202416 256022 202428
rect 258905 202419 258963 202425
rect 258905 202416 258917 202419
rect 256016 202388 258917 202416
rect 256016 202376 256022 202388
rect 258905 202385 258917 202388
rect 258951 202385 258963 202419
rect 258905 202379 258963 202385
rect 258997 202419 259055 202425
rect 258997 202385 259009 202419
rect 259043 202416 259055 202419
rect 268562 202416 268568 202428
rect 259043 202388 268568 202416
rect 259043 202385 259055 202388
rect 258997 202379 259055 202385
rect 268562 202376 268568 202388
rect 268620 202376 268626 202428
rect 275278 202376 275284 202428
rect 275336 202416 275342 202428
rect 285030 202416 285036 202428
rect 275336 202388 285036 202416
rect 275336 202376 275342 202388
rect 285030 202376 285036 202388
rect 285088 202376 285094 202428
rect 289262 202376 289268 202428
rect 289320 202416 289326 202428
rect 292500 202416 292528 202456
rect 298738 202444 298744 202456
rect 298796 202444 298802 202496
rect 299290 202444 299296 202496
rect 299348 202484 299354 202496
rect 325142 202484 325148 202496
rect 299348 202456 325148 202484
rect 299348 202444 299354 202456
rect 325142 202444 325148 202456
rect 325200 202444 325206 202496
rect 352742 202444 352748 202496
rect 352800 202484 352806 202496
rect 353202 202484 353208 202496
rect 352800 202456 353208 202484
rect 352800 202444 352806 202456
rect 353202 202444 353208 202456
rect 353260 202444 353266 202496
rect 358722 202444 358728 202496
rect 358780 202484 358786 202496
rect 359458 202484 359464 202496
rect 358780 202456 359464 202484
rect 358780 202444 358786 202456
rect 359458 202444 359464 202456
rect 359516 202444 359522 202496
rect 359553 202487 359611 202493
rect 359553 202453 359565 202487
rect 359599 202484 359611 202487
rect 393498 202484 393504 202496
rect 359599 202456 393504 202484
rect 359599 202453 359611 202456
rect 359553 202447 359611 202453
rect 393498 202444 393504 202456
rect 393556 202444 393562 202496
rect 289320 202388 292528 202416
rect 289320 202376 289326 202388
rect 298002 202376 298008 202428
rect 298060 202416 298066 202428
rect 306929 202419 306987 202425
rect 306929 202416 306941 202419
rect 298060 202388 306941 202416
rect 298060 202376 298066 202388
rect 306929 202385 306941 202388
rect 306975 202385 306987 202419
rect 306929 202379 306987 202385
rect 310606 202376 310612 202428
rect 310664 202416 310670 202428
rect 311250 202416 311256 202428
rect 310664 202388 311256 202416
rect 310664 202376 310670 202388
rect 311250 202376 311256 202388
rect 311308 202376 311314 202428
rect 311345 202419 311403 202425
rect 311345 202385 311357 202419
rect 311391 202416 311403 202419
rect 325694 202416 325700 202428
rect 311391 202388 325700 202416
rect 311391 202385 311403 202388
rect 311345 202379 311403 202385
rect 325694 202376 325700 202388
rect 325752 202376 325758 202428
rect 333146 202376 333152 202428
rect 333204 202416 333210 202428
rect 333882 202416 333888 202428
rect 333204 202388 333888 202416
rect 333204 202376 333210 202388
rect 333882 202376 333888 202388
rect 333940 202376 333946 202428
rect 348326 202376 348332 202428
rect 348384 202416 348390 202428
rect 390646 202416 390652 202428
rect 348384 202388 390652 202416
rect 348384 202376 348390 202388
rect 390646 202376 390652 202388
rect 390704 202376 390710 202428
rect 400950 202376 400956 202428
rect 401008 202416 401014 202428
rect 401502 202416 401508 202428
rect 401008 202388 401508 202416
rect 401008 202376 401014 202388
rect 401502 202376 401508 202388
rect 401560 202376 401566 202428
rect 140038 202308 140044 202360
rect 140096 202348 140102 202360
rect 168374 202348 168380 202360
rect 140096 202320 168380 202348
rect 140096 202308 140102 202320
rect 168374 202308 168380 202320
rect 168432 202308 168438 202360
rect 199102 202308 199108 202360
rect 199160 202348 199166 202360
rect 258442 202348 258448 202360
rect 199160 202320 258448 202348
rect 199160 202308 199166 202320
rect 258442 202308 258448 202320
rect 258500 202308 258506 202360
rect 261938 202348 261944 202360
rect 258552 202320 261944 202348
rect 151078 202240 151084 202292
rect 151136 202280 151142 202292
rect 181254 202280 181260 202292
rect 151136 202252 181260 202280
rect 151136 202240 151142 202252
rect 181254 202240 181260 202252
rect 181312 202240 181318 202292
rect 198918 202240 198924 202292
rect 198976 202280 198982 202292
rect 257065 202283 257123 202289
rect 257065 202280 257077 202283
rect 198976 202252 257077 202280
rect 198976 202240 198982 202252
rect 257065 202249 257077 202252
rect 257111 202249 257123 202283
rect 258552 202280 258580 202320
rect 261938 202308 261944 202320
rect 261996 202308 262002 202360
rect 265158 202308 265164 202360
rect 265216 202348 265222 202360
rect 266906 202348 266912 202360
rect 265216 202320 266912 202348
rect 265216 202308 265222 202320
rect 266906 202308 266912 202320
rect 266964 202308 266970 202360
rect 280982 202308 280988 202360
rect 281040 202348 281046 202360
rect 281442 202348 281448 202360
rect 281040 202320 281448 202348
rect 281040 202308 281046 202320
rect 281442 202308 281448 202320
rect 281500 202308 281506 202360
rect 282730 202308 282736 202360
rect 282788 202348 282794 202360
rect 294598 202348 294604 202360
rect 282788 202320 294604 202348
rect 282788 202308 282794 202320
rect 294598 202308 294604 202320
rect 294656 202308 294662 202360
rect 298554 202308 298560 202360
rect 298612 202348 298618 202360
rect 304994 202348 305000 202360
rect 298612 202320 305000 202348
rect 298612 202308 298618 202320
rect 304994 202308 305000 202320
rect 305052 202308 305058 202360
rect 307021 202351 307079 202357
rect 307021 202317 307033 202351
rect 307067 202348 307079 202351
rect 334618 202348 334624 202360
rect 307067 202320 334624 202348
rect 307067 202317 307079 202320
rect 307021 202311 307079 202317
rect 334618 202308 334624 202320
rect 334676 202308 334682 202360
rect 345750 202308 345756 202360
rect 345808 202348 345814 202360
rect 392026 202348 392032 202360
rect 345808 202320 392032 202348
rect 345808 202308 345814 202320
rect 392026 202308 392032 202320
rect 392084 202308 392090 202360
rect 257065 202243 257123 202249
rect 257172 202252 258580 202280
rect 258629 202283 258687 202289
rect 103330 202172 103336 202224
rect 103388 202212 103394 202224
rect 142522 202212 142528 202224
rect 103388 202184 142528 202212
rect 103388 202172 103394 202184
rect 142522 202172 142528 202184
rect 142580 202172 142586 202224
rect 146938 202172 146944 202224
rect 146996 202212 147002 202224
rect 180334 202212 180340 202224
rect 146996 202184 180340 202212
rect 146996 202172 147002 202184
rect 180334 202172 180340 202184
rect 180392 202172 180398 202224
rect 198826 202172 198832 202224
rect 198884 202212 198890 202224
rect 257172 202212 257200 202252
rect 258629 202249 258641 202283
rect 258675 202280 258687 202283
rect 266814 202280 266820 202292
rect 258675 202252 266820 202280
rect 258675 202249 258687 202252
rect 258629 202243 258687 202249
rect 266814 202240 266820 202252
rect 266872 202240 266878 202292
rect 283558 202240 283564 202292
rect 283616 202280 283622 202292
rect 337378 202280 337384 202292
rect 283616 202252 337384 202280
rect 283616 202240 283622 202252
rect 337378 202240 337384 202252
rect 337436 202240 337442 202292
rect 344002 202240 344008 202292
rect 344060 202280 344066 202292
rect 390554 202280 390560 202292
rect 344060 202252 390560 202280
rect 344060 202240 344066 202252
rect 390554 202240 390560 202252
rect 390612 202240 390618 202292
rect 414934 202240 414940 202292
rect 414992 202280 414998 202292
rect 503898 202280 503904 202292
rect 414992 202252 503904 202280
rect 414992 202240 414998 202252
rect 503898 202240 503904 202252
rect 503956 202240 503962 202292
rect 198884 202184 257200 202212
rect 257249 202215 257307 202221
rect 198884 202172 198890 202184
rect 257249 202181 257261 202215
rect 257295 202212 257307 202215
rect 260190 202212 260196 202224
rect 257295 202184 260196 202212
rect 257295 202181 257307 202184
rect 257249 202175 257307 202181
rect 260190 202172 260196 202184
rect 260248 202172 260254 202224
rect 275738 202172 275744 202224
rect 275796 202212 275802 202224
rect 287698 202212 287704 202224
rect 275796 202184 287704 202212
rect 275796 202172 275802 202184
rect 287698 202172 287704 202184
rect 287756 202172 287762 202224
rect 288802 202172 288808 202224
rect 288860 202212 288866 202224
rect 322198 202212 322204 202224
rect 288860 202184 322204 202212
rect 288860 202172 288866 202184
rect 322198 202172 322204 202184
rect 322256 202172 322262 202224
rect 332502 202172 332508 202224
rect 332560 202212 332566 202224
rect 391934 202212 391940 202224
rect 332560 202184 391940 202212
rect 332560 202172 332566 202184
rect 391934 202172 391940 202184
rect 391992 202172 391998 202224
rect 411070 202172 411076 202224
rect 411128 202212 411134 202224
rect 503806 202212 503812 202224
rect 411128 202184 503812 202212
rect 411128 202172 411134 202184
rect 503806 202172 503812 202184
rect 503864 202172 503870 202224
rect 93762 202104 93768 202156
rect 93820 202144 93826 202156
rect 134702 202144 134708 202156
rect 93820 202116 134708 202144
rect 93820 202104 93826 202116
rect 134702 202104 134708 202116
rect 134760 202104 134766 202156
rect 144178 202104 144184 202156
rect 144236 202144 144242 202156
rect 178678 202144 178684 202156
rect 144236 202116 178684 202144
rect 144236 202104 144242 202116
rect 178678 202104 178684 202116
rect 178736 202104 178742 202156
rect 197906 202104 197912 202156
rect 197964 202144 197970 202156
rect 269482 202144 269488 202156
rect 197964 202116 269488 202144
rect 197964 202104 197970 202116
rect 269482 202104 269488 202116
rect 269540 202104 269546 202156
rect 271690 202104 271696 202156
rect 271748 202144 271754 202156
rect 337470 202144 337476 202156
rect 271748 202116 337476 202144
rect 271748 202104 271754 202116
rect 337470 202104 337476 202116
rect 337528 202104 337534 202156
rect 342070 202104 342076 202156
rect 342128 202144 342134 202156
rect 393406 202144 393412 202156
rect 342128 202116 393412 202144
rect 342128 202104 342134 202116
rect 393406 202104 393412 202116
rect 393464 202104 393470 202156
rect 409230 202104 409236 202156
rect 409288 202144 409294 202156
rect 503714 202144 503720 202156
rect 409288 202116 503720 202144
rect 409288 202104 409294 202116
rect 503714 202104 503720 202116
rect 503772 202104 503778 202156
rect 200022 202036 200028 202088
rect 200080 202076 200086 202088
rect 215205 202079 215263 202085
rect 215205 202076 215217 202079
rect 200080 202048 215217 202076
rect 200080 202036 200086 202048
rect 215205 202045 215217 202048
rect 215251 202045 215263 202079
rect 215205 202039 215263 202045
rect 219253 202079 219311 202085
rect 219253 202045 219265 202079
rect 219299 202076 219311 202079
rect 233881 202079 233939 202085
rect 233881 202076 233893 202079
rect 219299 202048 233893 202076
rect 219299 202045 219311 202048
rect 219253 202039 219311 202045
rect 233881 202045 233893 202048
rect 233927 202045 233939 202079
rect 233881 202039 233939 202045
rect 236638 202036 236644 202088
rect 236696 202076 236702 202088
rect 237282 202076 237288 202088
rect 236696 202048 237288 202076
rect 236696 202036 236702 202048
rect 237282 202036 237288 202048
rect 237340 202036 237346 202088
rect 240962 202036 240968 202088
rect 241020 202076 241026 202088
rect 267274 202076 267280 202088
rect 241020 202048 267280 202076
rect 241020 202036 241026 202048
rect 267274 202036 267280 202048
rect 267332 202036 267338 202088
rect 299014 202036 299020 202088
rect 299072 202076 299078 202088
rect 311986 202076 311992 202088
rect 299072 202048 311992 202076
rect 299072 202036 299078 202048
rect 311986 202036 311992 202048
rect 312044 202036 312050 202088
rect 315298 202036 315304 202088
rect 315356 202076 315362 202088
rect 319438 202076 319444 202088
rect 315356 202048 319444 202076
rect 315356 202036 315362 202048
rect 319438 202036 319444 202048
rect 319496 202036 319502 202088
rect 351730 202036 351736 202088
rect 351788 202076 351794 202088
rect 359553 202079 359611 202085
rect 359553 202076 359565 202079
rect 351788 202048 359565 202076
rect 351788 202036 351794 202048
rect 359553 202045 359565 202048
rect 359599 202045 359611 202079
rect 359553 202039 359611 202045
rect 362862 202036 362868 202088
rect 362920 202076 362926 202088
rect 363690 202076 363696 202088
rect 362920 202048 363696 202076
rect 362920 202036 362926 202048
rect 363690 202036 363696 202048
rect 363748 202036 363754 202088
rect 199930 201968 199936 202020
rect 199988 202008 199994 202020
rect 219345 202011 219403 202017
rect 199988 201980 214512 202008
rect 199988 201968 199994 201980
rect 198642 201900 198648 201952
rect 198700 201940 198706 201952
rect 214285 201943 214343 201949
rect 214285 201940 214297 201943
rect 198700 201912 214297 201940
rect 198700 201900 198706 201912
rect 214285 201909 214297 201912
rect 214331 201909 214343 201943
rect 214285 201903 214343 201909
rect 198734 201832 198740 201884
rect 198792 201872 198798 201884
rect 211706 201872 211712 201884
rect 198792 201844 211712 201872
rect 198792 201832 198798 201844
rect 211706 201832 211712 201844
rect 211764 201832 211770 201884
rect 214484 201872 214512 201980
rect 219345 201977 219357 202011
rect 219391 202008 219403 202011
rect 232409 202011 232467 202017
rect 232409 202008 232421 202011
rect 219391 201980 232421 202008
rect 219391 201977 219403 201980
rect 219345 201971 219403 201977
rect 232409 201977 232421 201980
rect 232455 201977 232467 202011
rect 232409 201971 232467 201977
rect 232498 201968 232504 202020
rect 232556 202008 232562 202020
rect 236730 202008 236736 202020
rect 232556 201980 236736 202008
rect 232556 201968 232562 201980
rect 236730 201968 236736 201980
rect 236788 201968 236794 202020
rect 238110 201968 238116 202020
rect 238168 202008 238174 202020
rect 257525 202011 257583 202017
rect 257525 202008 257537 202011
rect 238168 201980 257537 202008
rect 238168 201968 238174 201980
rect 257525 201977 257537 201980
rect 257571 201977 257583 202011
rect 257525 201971 257583 201977
rect 258350 201968 258356 202020
rect 258408 202008 258414 202020
rect 258905 202011 258963 202017
rect 258408 201980 258856 202008
rect 258408 201968 258414 201980
rect 214561 201943 214619 201949
rect 214561 201909 214573 201943
rect 214607 201940 214619 201943
rect 216030 201940 216036 201952
rect 214607 201912 216036 201940
rect 214607 201909 214619 201912
rect 214561 201903 214619 201909
rect 216030 201900 216036 201912
rect 216088 201900 216094 201952
rect 247770 201940 247776 201952
rect 216140 201912 247776 201940
rect 215849 201875 215907 201881
rect 215849 201872 215861 201875
rect 214484 201844 215861 201872
rect 215849 201841 215861 201844
rect 215895 201841 215907 201875
rect 215849 201835 215907 201841
rect 215938 201832 215944 201884
rect 215996 201872 216002 201884
rect 216140 201872 216168 201912
rect 247770 201900 247776 201912
rect 247828 201900 247834 201952
rect 251450 201900 251456 201952
rect 251508 201940 251514 201952
rect 258828 201940 258856 201980
rect 258905 201977 258917 202011
rect 258951 202008 258963 202011
rect 268654 202008 268660 202020
rect 258951 201980 268660 202008
rect 258951 201977 258963 201980
rect 258905 201971 258963 201977
rect 268654 201968 268660 201980
rect 268712 201968 268718 202020
rect 291378 201968 291384 202020
rect 291436 202008 291442 202020
rect 292482 202008 292488 202020
rect 291436 201980 292488 202008
rect 291436 201968 291442 201980
rect 292482 201968 292488 201980
rect 292540 201968 292546 202020
rect 296162 201968 296168 202020
rect 296220 202008 296226 202020
rect 301498 202008 301504 202020
rect 296220 201980 301504 202008
rect 296220 201968 296226 201980
rect 301498 201968 301504 201980
rect 301556 201968 301562 202020
rect 306929 202011 306987 202017
rect 306929 201977 306941 202011
rect 306975 202008 306987 202011
rect 315390 202008 315396 202020
rect 306975 201980 315396 202008
rect 306975 201977 306987 201980
rect 306929 201971 306987 201977
rect 315390 201968 315396 201980
rect 315448 201968 315454 202020
rect 266538 201940 266544 201952
rect 251508 201912 258764 201940
rect 258828 201912 266544 201940
rect 251508 201900 251514 201912
rect 215996 201844 216168 201872
rect 216217 201875 216275 201881
rect 215996 201832 216002 201844
rect 216217 201841 216229 201875
rect 216263 201872 216275 201875
rect 242158 201872 242164 201884
rect 216263 201844 242164 201872
rect 216263 201841 216275 201844
rect 216217 201835 216275 201841
rect 242158 201832 242164 201844
rect 242216 201832 242222 201884
rect 248966 201832 248972 201884
rect 249024 201872 249030 201884
rect 258736 201872 258764 201912
rect 266538 201900 266544 201912
rect 266596 201900 266602 201952
rect 298370 201900 298376 201952
rect 298428 201940 298434 201952
rect 307021 201943 307079 201949
rect 307021 201940 307033 201943
rect 298428 201912 307033 201940
rect 298428 201900 298434 201912
rect 307021 201909 307033 201912
rect 307067 201909 307079 201943
rect 307021 201903 307079 201909
rect 249024 201844 258672 201872
rect 258736 201844 261064 201872
rect 249024 201832 249030 201844
rect 196802 201764 196808 201816
rect 196860 201804 196866 201816
rect 196860 201776 220768 201804
rect 196860 201764 196866 201776
rect 199286 201696 199292 201748
rect 199344 201736 199350 201748
rect 219526 201736 219532 201748
rect 199344 201708 219532 201736
rect 199344 201696 199350 201708
rect 219526 201696 219532 201708
rect 219584 201696 219590 201748
rect 220740 201736 220768 201776
rect 220814 201764 220820 201816
rect 220872 201804 220878 201816
rect 221274 201804 221280 201816
rect 220872 201776 221280 201804
rect 220872 201764 220878 201776
rect 221274 201764 221280 201776
rect 221332 201764 221338 201816
rect 229738 201764 229744 201816
rect 229796 201804 229802 201816
rect 237374 201804 237380 201816
rect 229796 201776 237380 201804
rect 229796 201764 229802 201776
rect 237374 201764 237380 201776
rect 237432 201764 237438 201816
rect 238018 201764 238024 201816
rect 238076 201804 238082 201816
rect 238076 201776 255176 201804
rect 238076 201764 238082 201776
rect 223022 201736 223028 201748
rect 220740 201708 223028 201736
rect 223022 201696 223028 201708
rect 223080 201696 223086 201748
rect 223117 201739 223175 201745
rect 223117 201705 223129 201739
rect 223163 201736 223175 201739
rect 223163 201708 241192 201736
rect 223163 201705 223175 201708
rect 223117 201699 223175 201705
rect 199562 201628 199568 201680
rect 199620 201668 199626 201680
rect 218606 201668 218612 201680
rect 199620 201640 218612 201668
rect 199620 201628 199626 201640
rect 218606 201628 218612 201640
rect 218664 201628 218670 201680
rect 233881 201671 233939 201677
rect 233881 201637 233893 201671
rect 233927 201668 233939 201671
rect 241054 201668 241060 201680
rect 233927 201640 241060 201668
rect 233927 201637 233939 201640
rect 233881 201631 233939 201637
rect 241054 201628 241060 201640
rect 241112 201628 241118 201680
rect 241164 201668 241192 201708
rect 242986 201696 242992 201748
rect 243044 201736 243050 201748
rect 244090 201736 244096 201748
rect 243044 201708 244096 201736
rect 243044 201696 243050 201708
rect 244090 201696 244096 201708
rect 244148 201696 244154 201748
rect 244918 201696 244924 201748
rect 244976 201736 244982 201748
rect 246022 201736 246028 201748
rect 244976 201708 246028 201736
rect 244976 201696 244982 201708
rect 246022 201696 246028 201708
rect 246080 201696 246086 201748
rect 250070 201696 250076 201748
rect 250128 201736 250134 201748
rect 250990 201736 250996 201748
rect 250128 201708 250996 201736
rect 250128 201696 250134 201708
rect 250990 201696 250996 201708
rect 251048 201696 251054 201748
rect 253106 201696 253112 201748
rect 253164 201736 253170 201748
rect 253750 201736 253756 201748
rect 253164 201708 253756 201736
rect 253164 201696 253170 201708
rect 253750 201696 253756 201708
rect 253808 201696 253814 201748
rect 255148 201736 255176 201776
rect 255222 201764 255228 201816
rect 255280 201804 255286 201816
rect 258537 201807 258595 201813
rect 258537 201804 258549 201807
rect 255280 201776 258549 201804
rect 255280 201764 255286 201776
rect 258537 201773 258549 201776
rect 258583 201773 258595 201807
rect 258644 201804 258672 201844
rect 258813 201807 258871 201813
rect 258813 201804 258825 201807
rect 258644 201776 258825 201804
rect 258537 201767 258595 201773
rect 258813 201773 258825 201776
rect 258859 201773 258871 201807
rect 258813 201767 258871 201773
rect 259454 201736 259460 201748
rect 255148 201708 259460 201736
rect 259454 201696 259460 201708
rect 259512 201696 259518 201748
rect 259549 201739 259607 201745
rect 259549 201705 259561 201739
rect 259595 201736 259607 201739
rect 260929 201739 260987 201745
rect 260929 201736 260941 201739
rect 259595 201708 260941 201736
rect 259595 201705 259607 201708
rect 259549 201699 259607 201705
rect 260929 201705 260941 201708
rect 260975 201705 260987 201739
rect 261036 201736 261064 201844
rect 266262 201832 266268 201884
rect 266320 201872 266326 201884
rect 269114 201872 269120 201884
rect 266320 201844 269120 201872
rect 266320 201832 266326 201844
rect 269114 201832 269120 201844
rect 269172 201832 269178 201884
rect 297726 201832 297732 201884
rect 297784 201872 297790 201884
rect 311345 201875 311403 201881
rect 311345 201872 311357 201875
rect 297784 201844 311357 201872
rect 297784 201832 297790 201844
rect 311345 201841 311357 201844
rect 311391 201841 311403 201875
rect 311345 201835 311403 201841
rect 264882 201764 264888 201816
rect 264940 201804 264946 201816
rect 267734 201804 267740 201816
rect 264940 201776 267740 201804
rect 264940 201764 264946 201776
rect 267734 201764 267740 201776
rect 267792 201764 267798 201816
rect 298646 201764 298652 201816
rect 298704 201804 298710 201816
rect 307757 201807 307815 201813
rect 307757 201804 307769 201807
rect 298704 201776 307769 201804
rect 298704 201764 298710 201776
rect 307757 201773 307769 201776
rect 307803 201773 307815 201807
rect 307757 201767 307815 201773
rect 314930 201764 314936 201816
rect 314988 201804 314994 201816
rect 315942 201804 315948 201816
rect 314988 201776 315948 201804
rect 314988 201764 314994 201776
rect 315942 201764 315948 201776
rect 316000 201764 316006 201816
rect 266630 201736 266636 201748
rect 261036 201708 266636 201736
rect 260929 201699 260987 201705
rect 266630 201696 266636 201708
rect 266688 201696 266694 201748
rect 267090 201696 267096 201748
rect 267148 201736 267154 201748
rect 268194 201736 268200 201748
rect 267148 201708 268200 201736
rect 267148 201696 267154 201708
rect 268194 201696 268200 201708
rect 268252 201696 268258 201748
rect 297818 201696 297824 201748
rect 297876 201736 297882 201748
rect 303890 201736 303896 201748
rect 297876 201708 303896 201736
rect 297876 201696 297882 201708
rect 303890 201696 303896 201708
rect 303948 201696 303954 201748
rect 306466 201696 306472 201748
rect 306524 201736 306530 201748
rect 307294 201736 307300 201748
rect 306524 201708 307300 201736
rect 306524 201696 306530 201708
rect 307294 201696 307300 201708
rect 307352 201696 307358 201748
rect 350994 201696 351000 201748
rect 351052 201736 351058 201748
rect 351822 201736 351828 201748
rect 351052 201708 351828 201736
rect 351052 201696 351058 201708
rect 351822 201696 351828 201708
rect 351880 201696 351886 201748
rect 355318 201696 355324 201748
rect 355376 201736 355382 201748
rect 355962 201736 355968 201748
rect 355376 201708 355968 201736
rect 355376 201696 355382 201708
rect 355962 201696 355968 201708
rect 356020 201696 356026 201748
rect 243170 201668 243176 201680
rect 241164 201640 243176 201668
rect 243170 201628 243176 201640
rect 243228 201628 243234 201680
rect 252370 201628 252376 201680
rect 252428 201668 252434 201680
rect 263594 201668 263600 201680
rect 252428 201640 263600 201668
rect 252428 201628 252434 201640
rect 263594 201628 263600 201640
rect 263652 201628 263658 201680
rect 273622 201628 273628 201680
rect 273680 201668 273686 201680
rect 279510 201668 279516 201680
rect 273680 201640 279516 201668
rect 273680 201628 273686 201640
rect 279510 201628 279516 201640
rect 279568 201628 279574 201680
rect 297542 201628 297548 201680
rect 297600 201668 297606 201680
rect 305638 201668 305644 201680
rect 297600 201640 305644 201668
rect 297600 201628 297606 201640
rect 305638 201628 305644 201640
rect 305696 201628 305702 201680
rect 353570 201628 353576 201680
rect 353628 201668 353634 201680
rect 356698 201668 356704 201680
rect 353628 201640 356704 201668
rect 353628 201628 353634 201640
rect 356698 201628 356704 201640
rect 356756 201628 356762 201680
rect 126330 201560 126336 201612
rect 126388 201600 126394 201612
rect 134150 201600 134156 201612
rect 126388 201572 134156 201600
rect 126388 201560 126394 201572
rect 134150 201560 134156 201572
rect 134208 201560 134214 201612
rect 199654 201560 199660 201612
rect 199712 201600 199718 201612
rect 216858 201600 216864 201612
rect 199712 201572 216864 201600
rect 199712 201560 199718 201572
rect 216858 201560 216864 201572
rect 216916 201560 216922 201612
rect 216953 201603 217011 201609
rect 216953 201569 216965 201603
rect 216999 201600 217011 201603
rect 219253 201603 219311 201609
rect 219253 201600 219265 201603
rect 216999 201572 219265 201600
rect 216999 201569 217011 201572
rect 216953 201563 217011 201569
rect 219253 201569 219265 201572
rect 219299 201569 219311 201603
rect 219253 201563 219311 201569
rect 232409 201603 232467 201609
rect 232409 201569 232421 201603
rect 232455 201600 232467 201603
rect 238202 201600 238208 201612
rect 232455 201572 238208 201600
rect 232455 201569 232467 201572
rect 232409 201563 232467 201569
rect 238202 201560 238208 201572
rect 238260 201560 238266 201612
rect 240045 201603 240103 201609
rect 240045 201569 240057 201603
rect 240091 201600 240103 201603
rect 245654 201600 245660 201612
rect 240091 201572 245660 201600
rect 240091 201569 240103 201572
rect 240045 201563 240103 201569
rect 245654 201560 245660 201572
rect 245712 201560 245718 201612
rect 257525 201603 257583 201609
rect 257525 201569 257537 201603
rect 257571 201600 257583 201603
rect 260834 201600 260840 201612
rect 257571 201572 260840 201600
rect 257571 201569 257583 201572
rect 257525 201563 257583 201569
rect 260834 201560 260840 201572
rect 260892 201560 260898 201612
rect 260929 201603 260987 201609
rect 260929 201569 260941 201603
rect 260975 201600 260987 201603
rect 266722 201600 266728 201612
rect 260975 201572 266728 201600
rect 260975 201569 260987 201572
rect 260929 201563 260987 201569
rect 266722 201560 266728 201572
rect 266780 201560 266786 201612
rect 266998 201560 267004 201612
rect 267056 201600 267062 201612
rect 267734 201600 267740 201612
rect 267056 201572 267740 201600
rect 267056 201560 267062 201572
rect 267734 201560 267740 201572
rect 267792 201560 267798 201612
rect 293770 201560 293776 201612
rect 293828 201600 293834 201612
rect 294690 201600 294696 201612
rect 293828 201572 294696 201600
rect 293828 201560 293834 201572
rect 294690 201560 294696 201572
rect 294748 201560 294754 201612
rect 308398 201560 308404 201612
rect 308456 201600 308462 201612
rect 308950 201600 308956 201612
rect 308456 201572 308956 201600
rect 308456 201560 308462 201572
rect 308950 201560 308956 201572
rect 309008 201560 309014 201612
rect 314654 201600 314660 201612
rect 309060 201572 314660 201600
rect 127618 201492 127624 201544
rect 127676 201532 127682 201544
rect 134334 201532 134340 201544
rect 127676 201504 134340 201532
rect 127676 201492 127682 201504
rect 134334 201492 134340 201504
rect 134392 201492 134398 201544
rect 198550 201492 198556 201544
rect 198608 201532 198614 201544
rect 202874 201532 202880 201544
rect 198608 201504 202880 201532
rect 198608 201492 198614 201504
rect 202874 201492 202880 201504
rect 202932 201492 202938 201544
rect 212442 201492 212448 201544
rect 212500 201532 212506 201544
rect 216217 201535 216275 201541
rect 216217 201532 216229 201535
rect 212500 201504 216229 201532
rect 212500 201492 212506 201504
rect 216217 201501 216229 201504
rect 216263 201501 216275 201535
rect 219345 201535 219403 201541
rect 219345 201532 219357 201535
rect 216217 201495 216275 201501
rect 216324 201504 219357 201532
rect 215849 201467 215907 201473
rect 215849 201433 215861 201467
rect 215895 201464 215907 201467
rect 216324 201464 216352 201504
rect 219345 201501 219357 201504
rect 219391 201501 219403 201535
rect 219345 201495 219403 201501
rect 220078 201492 220084 201544
rect 220136 201532 220142 201544
rect 223117 201535 223175 201541
rect 223117 201532 223129 201535
rect 220136 201504 223129 201532
rect 220136 201492 220142 201504
rect 223117 201501 223129 201504
rect 223163 201501 223175 201535
rect 223117 201495 223175 201501
rect 238941 201535 238999 201541
rect 238941 201501 238953 201535
rect 238987 201532 238999 201535
rect 246482 201532 246488 201544
rect 238987 201504 246488 201532
rect 238987 201501 238999 201504
rect 238941 201495 238999 201501
rect 246482 201492 246488 201504
rect 246540 201492 246546 201544
rect 254854 201492 254860 201544
rect 254912 201532 254918 201544
rect 259549 201535 259607 201541
rect 259549 201532 259561 201535
rect 254912 201504 259561 201532
rect 254912 201492 254918 201504
rect 259549 201501 259561 201504
rect 259595 201501 259607 201535
rect 259549 201495 259607 201501
rect 260098 201492 260104 201544
rect 260156 201532 260162 201544
rect 267642 201532 267648 201544
rect 260156 201504 267648 201532
rect 260156 201492 260162 201504
rect 267642 201492 267648 201504
rect 267700 201492 267706 201544
rect 293034 201492 293040 201544
rect 293092 201532 293098 201544
rect 293862 201532 293868 201544
rect 293092 201504 293868 201532
rect 293092 201492 293098 201504
rect 293862 201492 293868 201504
rect 293920 201492 293926 201544
rect 294414 201492 294420 201544
rect 294472 201532 294478 201544
rect 295242 201532 295248 201544
rect 294472 201504 295248 201532
rect 294472 201492 294478 201504
rect 295242 201492 295248 201504
rect 295300 201492 295306 201544
rect 295794 201492 295800 201544
rect 295852 201532 295858 201544
rect 296622 201532 296628 201544
rect 295852 201504 296628 201532
rect 295852 201492 295858 201504
rect 296622 201492 296628 201504
rect 296680 201492 296686 201544
rect 307018 201492 307024 201544
rect 307076 201532 307082 201544
rect 309060 201532 309088 201572
rect 314654 201560 314660 201572
rect 314712 201560 314718 201612
rect 307076 201504 309088 201532
rect 307076 201492 307082 201504
rect 316034 201492 316040 201544
rect 316092 201532 316098 201544
rect 317138 201532 317144 201544
rect 316092 201504 317144 201532
rect 316092 201492 316098 201504
rect 317138 201492 317144 201504
rect 317196 201492 317202 201544
rect 319070 201492 319076 201544
rect 319128 201532 319134 201544
rect 320082 201532 320088 201544
rect 319128 201504 320088 201532
rect 319128 201492 319134 201504
rect 320082 201492 320088 201504
rect 320140 201492 320146 201544
rect 320542 201492 320548 201544
rect 320600 201532 320606 201544
rect 321462 201532 321468 201544
rect 320600 201504 321468 201532
rect 320600 201492 320606 201504
rect 321462 201492 321468 201504
rect 321520 201492 321526 201544
rect 324038 201492 324044 201544
rect 324096 201532 324102 201544
rect 327074 201532 327080 201544
rect 324096 201504 327080 201532
rect 324096 201492 324102 201504
rect 327074 201492 327080 201504
rect 327132 201492 327138 201544
rect 410150 201492 410156 201544
rect 410208 201532 410214 201544
rect 411162 201532 411168 201544
rect 410208 201504 411168 201532
rect 410208 201492 410214 201504
rect 411162 201492 411168 201504
rect 411220 201492 411226 201544
rect 215895 201436 216352 201464
rect 215895 201433 215907 201436
rect 215849 201427 215907 201433
rect 215205 201399 215263 201405
rect 215205 201365 215217 201399
rect 215251 201396 215263 201399
rect 216953 201399 217011 201405
rect 216953 201396 216965 201399
rect 215251 201368 216965 201396
rect 215251 201365 215263 201368
rect 215205 201359 215263 201365
rect 216953 201365 216965 201368
rect 216999 201365 217011 201399
rect 216953 201359 217011 201365
rect 133506 201152 133512 201204
rect 133564 201192 133570 201204
rect 153378 201192 153384 201204
rect 133564 201164 153384 201192
rect 133564 201152 133570 201164
rect 153378 201152 153384 201164
rect 153436 201152 153442 201204
rect 3878 201084 3884 201136
rect 3936 201124 3942 201136
rect 436554 201124 436560 201136
rect 3936 201096 436560 201124
rect 3936 201084 3942 201096
rect 436554 201084 436560 201096
rect 436612 201084 436618 201136
rect 3602 201016 3608 201068
rect 3660 201056 3666 201068
rect 436462 201056 436468 201068
rect 3660 201028 436468 201056
rect 3660 201016 3666 201028
rect 436462 201016 436468 201028
rect 436520 201016 436526 201068
rect 3418 200948 3424 201000
rect 3476 200988 3482 201000
rect 436370 200988 436376 201000
rect 3476 200960 436376 200988
rect 3476 200948 3482 200960
rect 436370 200948 436376 200960
rect 436428 200948 436434 201000
rect 132402 200880 132408 200932
rect 132460 200920 132466 200932
rect 580258 200920 580264 200932
rect 132460 200892 580264 200920
rect 132460 200880 132466 200892
rect 580258 200880 580264 200892
rect 580316 200880 580322 200932
rect 132218 200812 132224 200864
rect 132276 200852 132282 200864
rect 580442 200852 580448 200864
rect 132276 200824 580448 200852
rect 132276 200812 132282 200824
rect 580442 200812 580448 200824
rect 580500 200812 580506 200864
rect 131390 200744 131396 200796
rect 131448 200784 131454 200796
rect 580350 200784 580356 200796
rect 131448 200756 580356 200784
rect 131448 200744 131454 200756
rect 580350 200744 580356 200756
rect 580408 200744 580414 200796
rect 209866 200200 209872 200252
rect 209924 200240 209930 200252
rect 210280 200240 210286 200252
rect 209924 200212 210286 200240
rect 209924 200200 209930 200212
rect 210280 200200 210286 200212
rect 210338 200200 210344 200252
rect 213914 200200 213920 200252
rect 213972 200240 213978 200252
rect 214604 200240 214610 200252
rect 213972 200212 214610 200240
rect 213972 200200 213978 200212
rect 214604 200200 214610 200212
rect 214662 200200 214668 200252
rect 3234 200132 3240 200184
rect 3292 200172 3298 200184
rect 436646 200172 436652 200184
rect 3292 200144 436652 200172
rect 3292 200132 3298 200144
rect 436646 200132 436652 200144
rect 436704 200132 436710 200184
rect 134061 200107 134119 200113
rect 134061 200073 134073 200107
rect 134107 200104 134119 200107
rect 134242 200104 134248 200116
rect 134107 200076 134248 200104
rect 134107 200073 134119 200076
rect 134061 200067 134119 200073
rect 134242 200064 134248 200076
rect 134300 200064 134306 200116
rect 238754 199860 238760 199912
rect 238812 199900 238818 199912
rect 239490 199900 239496 199912
rect 238812 199872 239496 199900
rect 238812 199860 238818 199872
rect 239490 199860 239496 199872
rect 239548 199860 239554 199912
rect 243078 199860 243084 199912
rect 243136 199900 243142 199912
rect 243814 199900 243820 199912
rect 243136 199872 243820 199900
rect 243136 199860 243142 199872
rect 243814 199860 243820 199872
rect 243872 199860 243878 199912
rect 133598 199792 133604 199844
rect 133656 199832 133662 199844
rect 580258 199832 580264 199844
rect 133656 199804 580264 199832
rect 133656 199792 133662 199804
rect 580258 199792 580264 199804
rect 580316 199792 580322 199844
rect 131390 198296 131396 198348
rect 131448 198336 131454 198348
rect 131485 198339 131543 198345
rect 131485 198336 131497 198339
rect 131448 198308 131497 198336
rect 131448 198296 131454 198308
rect 131485 198305 131497 198308
rect 131531 198305 131543 198339
rect 131485 198299 131543 198305
rect 3418 197344 3424 197396
rect 3476 197384 3482 197396
rect 131390 197384 131396 197396
rect 3476 197356 131396 197384
rect 3476 197344 3482 197356
rect 131390 197344 131396 197356
rect 131448 197344 131454 197396
rect 5350 196256 5356 196308
rect 5408 196296 5414 196308
rect 131390 196296 131396 196308
rect 5408 196268 131396 196296
rect 5408 196256 5414 196268
rect 131390 196256 131396 196268
rect 131448 196256 131454 196308
rect 17218 196052 17224 196104
rect 17276 196092 17282 196104
rect 130838 196092 130844 196104
rect 17276 196064 130844 196092
rect 17276 196052 17282 196064
rect 130838 196052 130844 196064
rect 130896 196052 130902 196104
rect 131758 196092 131764 196104
rect 131719 196064 131764 196092
rect 131758 196052 131764 196064
rect 131816 196052 131822 196104
rect 132862 196092 132868 196104
rect 132823 196064 132868 196092
rect 132862 196052 132868 196064
rect 132920 196052 132926 196104
rect 128538 195984 128544 196036
rect 128596 195984 128602 196036
rect 131390 195984 131396 196036
rect 131448 196024 131454 196036
rect 131485 196027 131543 196033
rect 131485 196024 131497 196027
rect 131448 195996 131497 196024
rect 131448 195984 131454 195996
rect 131485 195993 131497 195996
rect 131531 195993 131543 196027
rect 131485 195987 131543 195993
rect 128556 195888 128584 195984
rect 131758 195956 131764 195968
rect 131719 195928 131764 195956
rect 131758 195916 131764 195928
rect 131816 195916 131822 195968
rect 132862 195956 132868 195968
rect 132823 195928 132868 195956
rect 132862 195916 132868 195928
rect 132920 195916 132926 195968
rect 134058 195956 134064 195968
rect 134019 195928 134064 195956
rect 134058 195916 134064 195928
rect 134116 195916 134122 195968
rect 128630 195888 128636 195900
rect 128556 195860 128636 195888
rect 128630 195848 128636 195860
rect 128688 195848 128694 195900
rect 15838 194624 15844 194676
rect 15896 194664 15902 194676
rect 130838 194664 130844 194676
rect 15896 194636 130844 194664
rect 15896 194624 15902 194636
rect 130838 194624 130844 194636
rect 130896 194624 130902 194676
rect 14458 194488 14464 194540
rect 14516 194528 14522 194540
rect 130838 194528 130844 194540
rect 14516 194500 130844 194528
rect 14516 194488 14522 194500
rect 130838 194488 130844 194500
rect 130896 194488 130902 194540
rect 5258 193128 5264 193180
rect 5316 193168 5322 193180
rect 130746 193168 130752 193180
rect 5316 193140 130752 193168
rect 5316 193128 5322 193140
rect 130746 193128 130752 193140
rect 130804 193128 130810 193180
rect 5442 193060 5448 193112
rect 5500 193100 5506 193112
rect 130838 193100 130844 193112
rect 5500 193072 130844 193100
rect 5500 193060 5506 193072
rect 130838 193060 130844 193072
rect 130896 193060 130902 193112
rect 5166 191768 5172 191820
rect 5224 191808 5230 191820
rect 130838 191808 130844 191820
rect 5224 191780 130844 191808
rect 5224 191768 5230 191780
rect 130838 191768 130844 191780
rect 130896 191768 130902 191820
rect 128630 191740 128636 191752
rect 128591 191712 128636 191740
rect 128630 191700 128636 191712
rect 128688 191700 128694 191752
rect 128998 191740 129004 191752
rect 128959 191712 129004 191740
rect 128998 191700 129004 191712
rect 129056 191700 129062 191752
rect 5074 190408 5080 190460
rect 5132 190448 5138 190460
rect 130838 190448 130844 190460
rect 5132 190420 130844 190448
rect 5132 190408 5138 190420
rect 130838 190408 130844 190420
rect 130896 190408 130902 190460
rect 3510 188980 3516 189032
rect 3568 189020 3574 189032
rect 130746 189020 130752 189032
rect 3568 188992 130752 189020
rect 3568 188980 3574 188992
rect 130746 188980 130752 188992
rect 130804 188980 130810 189032
rect 4982 188912 4988 188964
rect 5040 188952 5046 188964
rect 130838 188952 130844 188964
rect 5040 188924 130844 188952
rect 5040 188912 5046 188924
rect 130838 188912 130844 188924
rect 130896 188912 130902 188964
rect 4890 187620 4896 187672
rect 4948 187660 4954 187672
rect 130838 187660 130844 187672
rect 4948 187632 130844 187660
rect 4948 187620 4954 187632
rect 130838 187620 130844 187632
rect 130896 187620 130902 187672
rect 4798 186260 4804 186312
rect 4856 186300 4862 186312
rect 131117 186303 131175 186309
rect 4856 186272 131068 186300
rect 4856 186260 4862 186272
rect 128630 186232 128636 186244
rect 128591 186204 128636 186232
rect 128630 186192 128636 186204
rect 128688 186192 128694 186244
rect 131040 186232 131068 186272
rect 131117 186269 131129 186303
rect 131163 186300 131175 186303
rect 131206 186300 131212 186312
rect 131163 186272 131212 186300
rect 131163 186269 131175 186272
rect 131117 186263 131175 186269
rect 131206 186260 131212 186272
rect 131264 186260 131270 186312
rect 131040 186204 131252 186232
rect 131224 186176 131252 186204
rect 131206 186124 131212 186176
rect 131264 186124 131270 186176
rect 13078 184832 13084 184884
rect 13136 184872 13142 184884
rect 131206 184872 131212 184884
rect 13136 184844 131212 184872
rect 13136 184832 13142 184844
rect 131206 184832 131212 184844
rect 131264 184832 131270 184884
rect 128998 183920 129004 183932
rect 128959 183892 129004 183920
rect 128998 183880 129004 183892
rect 129056 183880 129062 183932
rect 72418 183472 72424 183524
rect 72476 183512 72482 183524
rect 131206 183512 131212 183524
rect 72476 183484 131212 183512
rect 72476 183472 72482 183484
rect 131206 183472 131212 183484
rect 131264 183472 131270 183524
rect 131117 183379 131175 183385
rect 131117 183345 131129 183379
rect 131163 183376 131175 183379
rect 131206 183376 131212 183388
rect 131163 183348 131212 183376
rect 131163 183345 131175 183348
rect 131117 183339 131175 183345
rect 131206 183336 131212 183348
rect 131264 183336 131270 183388
rect 128814 182112 128820 182164
rect 128872 182112 128878 182164
rect 128633 182087 128691 182093
rect 128633 182053 128645 182087
rect 128679 182084 128691 182087
rect 128722 182084 128728 182096
rect 128679 182056 128728 182084
rect 128679 182053 128691 182056
rect 128633 182047 128691 182053
rect 128722 182044 128728 182056
rect 128780 182044 128786 182096
rect 128832 182084 128860 182112
rect 128906 182084 128912 182096
rect 128832 182056 128912 182084
rect 128906 182044 128912 182056
rect 128964 182044 128970 182096
rect 132862 181432 132868 181484
rect 132920 181472 132926 181484
rect 133322 181472 133328 181484
rect 132920 181444 133328 181472
rect 132920 181432 132926 181444
rect 133322 181432 133328 181444
rect 133380 181432 133386 181484
rect 2866 180752 2872 180804
rect 2924 180792 2930 180804
rect 15838 180792 15844 180804
rect 2924 180764 15844 180792
rect 2924 180752 2930 180764
rect 15838 180752 15844 180764
rect 15896 180752 15902 180804
rect 133966 180384 133972 180396
rect 133927 180356 133972 180384
rect 133966 180344 133972 180356
rect 134024 180344 134030 180396
rect 133874 176604 133880 176656
rect 133932 176644 133938 176656
rect 134058 176644 134064 176656
rect 133932 176616 134064 176644
rect 133932 176604 133938 176616
rect 134058 176604 134064 176616
rect 134116 176604 134122 176656
rect 504450 173884 504456 173936
rect 504508 173924 504514 173936
rect 504634 173924 504640 173936
rect 504508 173896 504640 173924
rect 504508 173884 504514 173896
rect 504634 173884 504640 173896
rect 504692 173884 504698 173936
rect 128630 172564 128636 172576
rect 128591 172536 128636 172564
rect 128630 172524 128636 172536
rect 128688 172524 128694 172576
rect 133966 172564 133972 172576
rect 133927 172536 133972 172564
rect 133966 172524 133972 172536
rect 134024 172524 134030 172576
rect 128906 167016 128912 167068
rect 128964 167016 128970 167068
rect 128924 166932 128952 167016
rect 128906 166880 128912 166932
rect 128964 166880 128970 166932
rect 132586 164704 132592 164756
rect 132644 164744 132650 164756
rect 133322 164744 133328 164756
rect 132644 164716 133328 164744
rect 132644 164704 132650 164716
rect 133322 164704 133328 164716
rect 133380 164704 133386 164756
rect 128630 164160 128636 164212
rect 128688 164200 128694 164212
rect 128722 164200 128728 164212
rect 128688 164172 128728 164200
rect 128688 164160 128694 164172
rect 128722 164160 128728 164172
rect 128780 164160 128786 164212
rect 132586 164160 132592 164212
rect 132644 164160 132650 164212
rect 504174 164160 504180 164212
rect 504232 164200 504238 164212
rect 504358 164200 504364 164212
rect 504232 164172 504364 164200
rect 504232 164160 504238 164172
rect 504358 164160 504364 164172
rect 504416 164160 504422 164212
rect 132604 164132 132632 164160
rect 132770 164132 132776 164144
rect 132604 164104 132776 164132
rect 132770 164092 132776 164104
rect 132828 164092 132834 164144
rect 128630 162840 128636 162852
rect 128591 162812 128636 162840
rect 128630 162800 128636 162812
rect 128688 162800 128694 162852
rect 133877 162843 133935 162849
rect 133877 162809 133889 162843
rect 133923 162840 133935 162843
rect 133966 162840 133972 162852
rect 133923 162812 133972 162840
rect 133923 162809 133935 162812
rect 133877 162803 133935 162809
rect 133966 162800 133972 162812
rect 134024 162800 134030 162852
rect 436830 157360 436836 157412
rect 436888 157400 436894 157412
rect 580166 157400 580172 157412
rect 436888 157372 580172 157400
rect 436888 157360 436894 157372
rect 580166 157360 580172 157372
rect 580224 157360 580230 157412
rect 131114 156272 131120 156324
rect 131172 156312 131178 156324
rect 131172 156284 131436 156312
rect 131172 156272 131178 156284
rect 3510 156068 3516 156120
rect 3568 156108 3574 156120
rect 131298 156108 131304 156120
rect 3568 156080 131304 156108
rect 3568 156068 3574 156080
rect 131298 156068 131304 156080
rect 131356 156068 131362 156120
rect 3234 156000 3240 156052
rect 3292 156040 3298 156052
rect 131114 156040 131120 156052
rect 3292 156012 131120 156040
rect 3292 156000 3298 156012
rect 131114 156000 131120 156012
rect 131172 156000 131178 156052
rect 131298 155932 131304 155984
rect 131356 155972 131362 155984
rect 131408 155972 131436 156284
rect 131356 155944 131436 155972
rect 131356 155932 131362 155944
rect 3602 155864 3608 155916
rect 3660 155904 3666 155916
rect 131114 155904 131120 155916
rect 3660 155876 131120 155904
rect 3660 155864 3666 155876
rect 131114 155864 131120 155876
rect 131172 155864 131178 155916
rect 436094 155184 436100 155236
rect 436152 155224 436158 155236
rect 438118 155224 438124 155236
rect 436152 155196 438124 155224
rect 436152 155184 436158 155196
rect 438118 155184 438124 155196
rect 438176 155184 438182 155236
rect 131206 155048 131212 155100
rect 131264 155088 131270 155100
rect 132678 155088 132684 155100
rect 131264 155060 132684 155088
rect 131264 155048 131270 155060
rect 132678 155048 132684 155060
rect 132736 155048 132742 155100
rect 57977 154547 58035 154553
rect 57977 154544 57989 154547
rect 31680 154516 57989 154544
rect 31680 154476 31708 154516
rect 57977 154513 57989 154516
rect 58023 154513 58035 154547
rect 99285 154547 99343 154553
rect 99285 154544 99297 154547
rect 57977 154507 58035 154513
rect 89640 154516 99297 154544
rect 22112 154448 31708 154476
rect 67545 154479 67603 154485
rect 19245 154411 19303 154417
rect 19245 154377 19257 154411
rect 19291 154408 19303 154411
rect 22112 154408 22140 154448
rect 67545 154445 67557 154479
rect 67591 154476 67603 154479
rect 89640 154476 89668 154516
rect 99285 154513 99297 154516
rect 99331 154513 99343 154547
rect 99285 154507 99343 154513
rect 109037 154547 109095 154553
rect 109037 154513 109049 154547
rect 109083 154544 109095 154547
rect 118605 154547 118663 154553
rect 118605 154544 118617 154547
rect 109083 154516 118617 154544
rect 109083 154513 109095 154516
rect 109037 154507 109095 154513
rect 118605 154513 118617 154516
rect 118651 154513 118663 154547
rect 118605 154507 118663 154513
rect 67591 154448 70348 154476
rect 67591 154445 67603 154448
rect 67545 154439 67603 154445
rect 19291 154380 22140 154408
rect 70320 154408 70348 154448
rect 86880 154448 89668 154476
rect 99469 154479 99527 154485
rect 80057 154411 80115 154417
rect 80057 154408 80069 154411
rect 70320 154380 80069 154408
rect 19291 154377 19303 154380
rect 19245 154371 19303 154377
rect 80057 154377 80069 154380
rect 80103 154377 80115 154411
rect 80057 154371 80115 154377
rect 80149 154411 80207 154417
rect 80149 154377 80161 154411
rect 80195 154408 80207 154411
rect 86880 154408 86908 154448
rect 99469 154445 99481 154479
rect 99515 154476 99527 154479
rect 118789 154479 118847 154485
rect 99515 154448 108988 154476
rect 99515 154445 99527 154448
rect 99469 154439 99527 154445
rect 80195 154380 86908 154408
rect 108960 154408 108988 154448
rect 118789 154445 118801 154479
rect 118835 154476 118847 154479
rect 118835 154448 128308 154476
rect 118835 154445 118847 154448
rect 118789 154439 118847 154445
rect 109037 154411 109095 154417
rect 109037 154408 109049 154411
rect 108960 154380 109049 154408
rect 80195 154377 80207 154380
rect 80149 154371 80207 154377
rect 109037 154377 109049 154380
rect 109083 154377 109095 154411
rect 128280 154408 128308 154448
rect 131114 154408 131120 154420
rect 128280 154380 131120 154408
rect 109037 154371 109095 154377
rect 131114 154368 131120 154380
rect 131172 154368 131178 154420
rect 3326 154300 3332 154352
rect 3384 154340 3390 154352
rect 9677 154343 9735 154349
rect 9677 154340 9689 154343
rect 3384 154312 9689 154340
rect 3384 154300 3390 154312
rect 9677 154309 9689 154312
rect 9723 154309 9735 154343
rect 9677 154303 9735 154309
rect 57977 154343 58035 154349
rect 57977 154309 57989 154343
rect 58023 154340 58035 154343
rect 67545 154343 67603 154349
rect 67545 154340 67557 154343
rect 58023 154312 67557 154340
rect 58023 154309 58035 154312
rect 57977 154303 58035 154309
rect 67545 154309 67557 154312
rect 67591 154309 67603 154343
rect 67545 154303 67603 154309
rect 9677 154207 9735 154213
rect 9677 154173 9689 154207
rect 9723 154204 9735 154207
rect 19245 154207 19303 154213
rect 19245 154204 19257 154207
rect 9723 154176 19257 154204
rect 9723 154173 9735 154176
rect 9677 154167 9735 154173
rect 19245 154173 19257 154176
rect 19291 154173 19303 154207
rect 19245 154167 19303 154173
rect 128630 153252 128636 153264
rect 128591 153224 128636 153252
rect 128630 153212 128636 153224
rect 128688 153212 128694 153264
rect 4062 153144 4068 153196
rect 4120 153184 4126 153196
rect 131114 153184 131120 153196
rect 4120 153156 131120 153184
rect 4120 153144 4126 153156
rect 131114 153144 131120 153156
rect 131172 153144 131178 153196
rect 437382 153144 437388 153196
rect 437440 153184 437446 153196
rect 447778 153184 447784 153196
rect 437440 153156 447784 153184
rect 437440 153144 437446 153156
rect 447778 153144 447784 153156
rect 447836 153144 447842 153196
rect 32401 153119 32459 153125
rect 32401 153085 32413 153119
rect 32447 153116 32459 153119
rect 108945 153119 109003 153125
rect 108945 153116 108957 153119
rect 32447 153088 60780 153116
rect 32447 153085 32459 153088
rect 32401 153079 32459 153085
rect 22741 153051 22799 153057
rect 22741 153017 22753 153051
rect 22787 153048 22799 153051
rect 27617 153051 27675 153057
rect 27617 153048 27629 153051
rect 22787 153020 27629 153048
rect 22787 153017 22799 153020
rect 22741 153011 22799 153017
rect 27617 153017 27629 153020
rect 27663 153017 27675 153051
rect 60752 153048 60780 153088
rect 89640 153088 108957 153116
rect 86865 153051 86923 153057
rect 60752 153020 70348 153048
rect 27617 153011 27675 153017
rect 70320 152980 70348 153020
rect 86865 153017 86877 153051
rect 86911 153048 86923 153051
rect 89640 153048 89668 153088
rect 108945 153085 108957 153088
rect 108991 153085 109003 153119
rect 115937 153119 115995 153125
rect 115937 153116 115949 153119
rect 108945 153079 109003 153085
rect 115860 153088 115949 153116
rect 115860 153057 115888 153088
rect 115937 153085 115949 153088
rect 115983 153085 115995 153119
rect 131298 153116 131304 153128
rect 131259 153088 131304 153116
rect 115937 153079 115995 153085
rect 131298 153076 131304 153088
rect 131356 153076 131362 153128
rect 86911 153020 89668 153048
rect 115845 153051 115903 153057
rect 86911 153017 86923 153020
rect 86865 153011 86923 153017
rect 115845 153017 115857 153051
rect 115891 153017 115903 153051
rect 115845 153011 115903 153017
rect 125505 153051 125563 153057
rect 125505 153017 125517 153051
rect 125551 153048 125563 153051
rect 125551 153020 128308 153048
rect 125551 153017 125563 153020
rect 125505 153011 125563 153017
rect 77297 152983 77355 152989
rect 77297 152980 77309 152983
rect 9600 152952 9720 152980
rect 70320 152952 77309 152980
rect 3970 152872 3976 152924
rect 4028 152912 4034 152924
rect 9600 152912 9628 152952
rect 4028 152884 9628 152912
rect 9692 152912 9720 152952
rect 77297 152949 77309 152952
rect 77343 152949 77355 152983
rect 128280 152980 128308 153020
rect 131298 152980 131304 152992
rect 128280 152952 131304 152980
rect 77297 152943 77355 152949
rect 131298 152940 131304 152952
rect 131356 152940 131362 152992
rect 17957 152915 18015 152921
rect 17957 152912 17969 152915
rect 9692 152884 17969 152912
rect 4028 152872 4034 152884
rect 17957 152881 17969 152884
rect 18003 152881 18015 152915
rect 17957 152875 18015 152881
rect 27617 152915 27675 152921
rect 27617 152881 27629 152915
rect 27663 152912 27675 152915
rect 32401 152915 32459 152921
rect 32401 152912 32413 152915
rect 27663 152884 32413 152912
rect 27663 152881 27675 152884
rect 27617 152875 27675 152881
rect 32401 152881 32413 152884
rect 32447 152881 32459 152915
rect 32401 152875 32459 152881
rect 108945 152915 109003 152921
rect 108945 152881 108957 152915
rect 108991 152912 109003 152915
rect 115845 152915 115903 152921
rect 115845 152912 115857 152915
rect 108991 152884 115857 152912
rect 108991 152881 109003 152884
rect 108945 152875 109003 152881
rect 115845 152881 115857 152884
rect 115891 152881 115903 152915
rect 115845 152875 115903 152881
rect 115937 152915 115995 152921
rect 115937 152881 115949 152915
rect 115983 152912 115995 152915
rect 125505 152915 125563 152921
rect 125505 152912 125517 152915
rect 115983 152884 125517 152912
rect 115983 152881 115995 152884
rect 115937 152875 115995 152881
rect 125505 152881 125517 152884
rect 125551 152881 125563 152915
rect 125505 152875 125563 152881
rect 77297 152847 77355 152853
rect 77297 152813 77309 152847
rect 77343 152844 77355 152847
rect 86865 152847 86923 152853
rect 86865 152844 86877 152847
rect 77343 152816 86877 152844
rect 77343 152813 77355 152816
rect 77297 152807 77355 152813
rect 86865 152813 86877 152816
rect 86911 152813 86923 152847
rect 86865 152807 86923 152813
rect 17957 152779 18015 152785
rect 17957 152745 17969 152779
rect 18003 152776 18015 152779
rect 22741 152779 22799 152785
rect 22741 152776 22753 152779
rect 18003 152748 22753 152776
rect 18003 152745 18015 152748
rect 17957 152739 18015 152745
rect 22741 152745 22753 152748
rect 22787 152745 22799 152779
rect 22741 152739 22799 152745
rect 131298 151892 131304 151904
rect 131259 151864 131304 151892
rect 131298 151852 131304 151864
rect 131356 151852 131362 151904
rect 3786 151716 3792 151768
rect 3844 151756 3850 151768
rect 131114 151756 131120 151768
rect 3844 151728 131120 151756
rect 3844 151716 3850 151728
rect 131114 151716 131120 151728
rect 131172 151716 131178 151768
rect 3694 150356 3700 150408
rect 3752 150396 3758 150408
rect 131114 150396 131120 150408
rect 3752 150368 131120 150396
rect 3752 150356 3758 150368
rect 131114 150356 131120 150368
rect 131172 150356 131178 150408
rect 437382 150356 437388 150408
rect 437440 150396 437446 150408
rect 446398 150396 446404 150408
rect 437440 150368 446404 150396
rect 437440 150356 437446 150368
rect 446398 150356 446404 150368
rect 446456 150356 446462 150408
rect 28258 148996 28264 149048
rect 28316 149036 28322 149048
rect 28316 149008 131252 149036
rect 28316 148996 28322 149008
rect 31018 148928 31024 148980
rect 31076 148968 31082 148980
rect 131114 148968 131120 148980
rect 31076 148940 131120 148968
rect 31076 148928 31082 148940
rect 131114 148928 131120 148940
rect 131172 148928 131178 148980
rect 131224 148900 131252 149008
rect 436094 148996 436100 149048
rect 436152 149036 436158 149048
rect 445018 149036 445024 149048
rect 436152 149008 445024 149036
rect 436152 148996 436158 149008
rect 445018 148996 445024 149008
rect 445076 148996 445082 149048
rect 131132 148872 131252 148900
rect 131132 148640 131160 148872
rect 131114 148588 131120 148640
rect 131172 148588 131178 148640
rect 128630 147744 128636 147756
rect 128591 147716 128636 147744
rect 128630 147704 128636 147716
rect 128688 147704 128694 147756
rect 21358 147568 21364 147620
rect 21416 147608 21422 147620
rect 131206 147608 131212 147620
rect 21416 147580 131068 147608
rect 131167 147580 131212 147608
rect 21416 147568 21422 147580
rect 128630 147540 128636 147552
rect 128591 147512 128636 147540
rect 128630 147500 128636 147512
rect 128688 147500 128694 147552
rect 131040 147472 131068 147580
rect 131206 147568 131212 147580
rect 131264 147568 131270 147620
rect 131206 147472 131212 147484
rect 131040 147444 131212 147472
rect 131206 147432 131212 147444
rect 131264 147432 131270 147484
rect 19978 146208 19984 146260
rect 20036 146248 20042 146260
rect 131114 146248 131120 146260
rect 20036 146220 131120 146248
rect 20036 146208 20042 146220
rect 131114 146208 131120 146220
rect 131172 146208 131178 146260
rect 437382 146140 437388 146192
rect 437440 146180 437446 146192
rect 442258 146180 442264 146192
rect 437440 146152 442264 146180
rect 437440 146140 437446 146152
rect 442258 146140 442264 146152
rect 442316 146140 442322 146192
rect 128906 144916 128912 144968
rect 128964 144916 128970 144968
rect 67637 144891 67695 144897
rect 67637 144857 67649 144891
rect 67683 144888 67695 144891
rect 79965 144891 80023 144897
rect 79965 144888 79977 144891
rect 67683 144860 79977 144888
rect 67683 144857 67695 144860
rect 67637 144851 67695 144857
rect 79965 144857 79977 144860
rect 80011 144857 80023 144891
rect 79965 144851 80023 144857
rect 96525 144891 96583 144897
rect 96525 144857 96537 144891
rect 96571 144888 96583 144891
rect 99285 144891 99343 144897
rect 99285 144888 99297 144891
rect 96571 144860 99297 144888
rect 96571 144857 96583 144860
rect 96525 144851 96583 144857
rect 99285 144857 99297 144860
rect 99331 144857 99343 144891
rect 99285 144851 99343 144857
rect 109037 144891 109095 144897
rect 109037 144857 109049 144891
rect 109083 144888 109095 144891
rect 118605 144891 118663 144897
rect 118605 144888 118617 144891
rect 109083 144860 118617 144888
rect 109083 144857 109095 144860
rect 109037 144851 109095 144857
rect 118605 144857 118617 144860
rect 118651 144857 118663 144891
rect 118605 144851 118663 144857
rect 128814 144848 128820 144900
rect 128872 144888 128878 144900
rect 128924 144888 128952 144916
rect 128872 144860 128952 144888
rect 128872 144848 128878 144860
rect 437014 144848 437020 144900
rect 437072 144888 437078 144900
rect 514018 144888 514024 144900
rect 437072 144860 514024 144888
rect 437072 144848 437078 144860
rect 514018 144848 514024 144860
rect 514076 144848 514082 144900
rect 99469 144823 99527 144829
rect 99469 144789 99481 144823
rect 99515 144820 99527 144823
rect 99515 144792 108988 144820
rect 99515 144789 99527 144792
rect 99469 144783 99527 144789
rect 38565 144755 38623 144761
rect 38565 144721 38577 144755
rect 38611 144752 38623 144755
rect 41325 144755 41383 144761
rect 41325 144752 41337 144755
rect 38611 144724 41337 144752
rect 38611 144721 38623 144724
rect 38565 144715 38623 144721
rect 41325 144721 41337 144724
rect 41371 144721 41383 144755
rect 41325 144715 41383 144721
rect 41417 144755 41475 144761
rect 41417 144721 41429 144755
rect 41463 144752 41475 144755
rect 57885 144755 57943 144761
rect 41463 144724 42656 144752
rect 41463 144721 41475 144724
rect 41417 144715 41475 144721
rect 24762 144644 24768 144696
rect 24820 144684 24826 144696
rect 28997 144687 29055 144693
rect 28997 144684 29009 144687
rect 24820 144656 29009 144684
rect 24820 144644 24826 144656
rect 28997 144653 29009 144656
rect 29043 144653 29055 144687
rect 42628 144684 42656 144724
rect 57885 144721 57897 144755
rect 57931 144752 57943 144755
rect 60645 144755 60703 144761
rect 60645 144752 60657 144755
rect 57931 144724 60657 144752
rect 57931 144721 57943 144724
rect 57885 144715 57943 144721
rect 60645 144721 60657 144724
rect 60691 144721 60703 144755
rect 60645 144715 60703 144721
rect 60737 144755 60795 144761
rect 60737 144721 60749 144755
rect 60783 144752 60795 144755
rect 80149 144755 80207 144761
rect 60783 144724 61976 144752
rect 60783 144721 60795 144724
rect 60737 144715 60795 144721
rect 48317 144687 48375 144693
rect 48317 144684 48329 144687
rect 42628 144656 48329 144684
rect 28997 144647 29055 144653
rect 48317 144653 48329 144656
rect 48363 144653 48375 144687
rect 61948 144684 61976 144724
rect 80149 144721 80161 144755
rect 80195 144752 80207 144755
rect 86957 144755 87015 144761
rect 86957 144752 86969 144755
rect 80195 144724 86969 144752
rect 80195 144721 80207 144724
rect 80149 144715 80207 144721
rect 86957 144721 86969 144724
rect 87003 144721 87015 144755
rect 108960 144752 108988 144792
rect 109037 144755 109095 144761
rect 109037 144752 109049 144755
rect 108960 144724 109049 144752
rect 86957 144715 87015 144721
rect 109037 144721 109049 144724
rect 109083 144721 109095 144755
rect 109037 144715 109095 144721
rect 118789 144755 118847 144761
rect 118789 144721 118801 144755
rect 118835 144752 118847 144755
rect 128170 144752 128176 144764
rect 118835 144724 128176 144752
rect 118835 144721 118847 144724
rect 118789 144715 118847 144721
rect 128170 144712 128176 144724
rect 128228 144712 128234 144764
rect 67637 144687 67695 144693
rect 67637 144684 67649 144687
rect 61948 144656 67649 144684
rect 48317 144647 48375 144653
rect 67637 144653 67649 144656
rect 67683 144653 67695 144687
rect 67637 144647 67695 144653
rect 86957 144619 87015 144625
rect 86957 144585 86969 144619
rect 87003 144616 87015 144619
rect 96525 144619 96583 144625
rect 96525 144616 96537 144619
rect 87003 144588 96537 144616
rect 87003 144585 87015 144588
rect 86957 144579 87015 144585
rect 96525 144585 96537 144588
rect 96571 144585 96583 144619
rect 96525 144579 96583 144585
rect 28997 144551 29055 144557
rect 28997 144517 29009 144551
rect 29043 144548 29055 144551
rect 38565 144551 38623 144557
rect 38565 144548 38577 144551
rect 29043 144520 38577 144548
rect 29043 144517 29055 144520
rect 28997 144511 29055 144517
rect 38565 144517 38577 144520
rect 38611 144517 38623 144551
rect 38565 144511 38623 144517
rect 48317 144551 48375 144557
rect 48317 144517 48329 144551
rect 48363 144548 48375 144551
rect 57885 144551 57943 144557
rect 57885 144548 57897 144551
rect 48363 144520 57897 144548
rect 48363 144517 48375 144520
rect 48317 144511 48375 144517
rect 57885 144517 57897 144520
rect 57931 144517 57943 144551
rect 57885 144511 57943 144517
rect 126238 144372 126244 144424
rect 126296 144412 126302 144424
rect 131114 144412 131120 144424
rect 126296 144384 131120 144412
rect 126296 144372 126302 144384
rect 131114 144372 131120 144384
rect 131172 144372 131178 144424
rect 133877 143599 133935 143605
rect 133877 143565 133889 143599
rect 133923 143596 133935 143599
rect 133966 143596 133972 143608
rect 133923 143568 133972 143596
rect 133923 143565 133935 143568
rect 133877 143559 133935 143565
rect 133966 143556 133972 143568
rect 134024 143556 134030 143608
rect 132678 142100 132684 142112
rect 132639 142072 132684 142100
rect 132678 142060 132684 142072
rect 132736 142060 132742 142112
rect 436094 142060 436100 142112
rect 436152 142100 436158 142112
rect 438210 142100 438216 142112
rect 436152 142072 438216 142100
rect 436152 142060 436158 142072
rect 438210 142060 438216 142072
rect 438268 142060 438274 142112
rect 133874 138660 133880 138712
rect 133932 138700 133938 138712
rect 133932 138672 133977 138700
rect 133932 138660 133938 138672
rect 437382 137912 437388 137964
rect 437440 137952 437446 137964
rect 580534 137952 580540 137964
rect 437440 137924 580540 137952
rect 437440 137912 437446 137924
rect 580534 137912 580540 137924
rect 580592 137912 580598 137964
rect 3326 136552 3332 136604
rect 3384 136592 3390 136604
rect 17218 136592 17224 136604
rect 3384 136564 17224 136592
rect 3384 136552 3390 136564
rect 17218 136552 17224 136564
rect 17276 136552 17282 136604
rect 437014 136552 437020 136604
rect 437072 136592 437078 136604
rect 504450 136592 504456 136604
rect 437072 136564 504456 136592
rect 437072 136552 437078 136564
rect 504450 136552 504456 136564
rect 504508 136552 504514 136604
rect 132681 135235 132739 135241
rect 132681 135201 132693 135235
rect 132727 135232 132739 135235
rect 132770 135232 132776 135244
rect 132727 135204 132776 135232
rect 132727 135201 132739 135204
rect 132681 135195 132739 135201
rect 132770 135192 132776 135204
rect 132828 135192 132834 135244
rect 437382 133832 437388 133884
rect 437440 133872 437446 133884
rect 580626 133872 580632 133884
rect 437440 133844 580632 133872
rect 437440 133832 437446 133844
rect 580626 133832 580632 133844
rect 580684 133832 580690 133884
rect 128630 132812 128636 132864
rect 128688 132852 128694 132864
rect 128814 132852 128820 132864
rect 128688 132824 128820 132852
rect 128688 132812 128694 132824
rect 128814 132812 128820 132824
rect 128872 132812 128878 132864
rect 131206 132512 131212 132524
rect 131167 132484 131212 132512
rect 131206 132472 131212 132484
rect 131264 132472 131270 132524
rect 132681 132447 132739 132453
rect 132681 132413 132693 132447
rect 132727 132444 132739 132447
rect 132770 132444 132776 132456
rect 132727 132416 132776 132444
rect 132727 132413 132739 132416
rect 132681 132407 132739 132413
rect 132770 132404 132776 132416
rect 132828 132404 132834 132456
rect 437382 132404 437388 132456
rect 437440 132444 437446 132456
rect 580718 132444 580724 132456
rect 437440 132416 580724 132444
rect 437440 132404 437446 132416
rect 580718 132404 580724 132416
rect 580776 132404 580782 132456
rect 437382 129684 437388 129736
rect 437440 129724 437446 129736
rect 580810 129724 580816 129736
rect 437440 129696 580816 129724
rect 437440 129684 437446 129696
rect 580810 129684 580816 129696
rect 580868 129684 580874 129736
rect 131114 125604 131120 125656
rect 131172 125644 131178 125656
rect 131206 125644 131212 125656
rect 131172 125616 131212 125644
rect 131172 125604 131178 125616
rect 131206 125604 131212 125616
rect 131264 125604 131270 125656
rect 133874 125644 133880 125656
rect 133835 125616 133880 125644
rect 133874 125604 133880 125616
rect 133932 125604 133938 125656
rect 131114 124148 131120 124160
rect 131075 124120 131120 124148
rect 131114 124108 131120 124120
rect 131172 124108 131178 124160
rect 133874 121184 133880 121236
rect 133932 121224 133938 121236
rect 580534 121224 580540 121236
rect 133932 121196 580540 121224
rect 133932 121184 133938 121196
rect 580534 121184 580540 121196
rect 580592 121184 580598 121236
rect 132402 121116 132408 121168
rect 132460 121156 132466 121168
rect 580350 121156 580356 121168
rect 132460 121128 580356 121156
rect 132460 121116 132466 121128
rect 580350 121116 580356 121128
rect 580408 121116 580414 121168
rect 133966 121048 133972 121100
rect 134024 121088 134030 121100
rect 580258 121088 580264 121100
rect 134024 121060 580264 121088
rect 134024 121048 134030 121060
rect 580258 121048 580264 121060
rect 580316 121048 580322 121100
rect 3050 120980 3056 121032
rect 3108 121020 3114 121032
rect 436278 121020 436284 121032
rect 3108 120992 436284 121020
rect 3108 120980 3114 120992
rect 436278 120980 436284 120992
rect 436336 120980 436342 121032
rect 134058 120912 134064 120964
rect 134116 120952 134122 120964
rect 138845 120955 138903 120961
rect 138845 120952 138857 120955
rect 134116 120924 138857 120952
rect 134116 120912 134122 120924
rect 138845 120921 138857 120924
rect 138891 120921 138903 120955
rect 138845 120915 138903 120921
rect 180978 119756 180984 119808
rect 181036 119796 181042 119808
rect 182036 119796 182042 119808
rect 181036 119768 182042 119796
rect 181036 119756 181042 119768
rect 182036 119756 182042 119768
rect 182094 119756 182100 119808
rect 185118 119756 185124 119808
rect 185176 119796 185182 119808
rect 185716 119796 185722 119808
rect 185176 119768 185722 119796
rect 185176 119756 185182 119768
rect 185716 119756 185722 119768
rect 185774 119756 185780 119808
rect 138290 119348 138296 119400
rect 138348 119388 138354 119400
rect 138842 119388 138848 119400
rect 138348 119360 138848 119388
rect 138348 119348 138354 119360
rect 138842 119348 138848 119360
rect 138900 119348 138906 119400
rect 143626 119348 143632 119400
rect 143684 119388 143690 119400
rect 144362 119388 144368 119400
rect 143684 119360 144368 119388
rect 143684 119348 143690 119360
rect 144362 119348 144368 119360
rect 144420 119348 144426 119400
rect 67542 119076 67548 119128
rect 67600 119116 67606 119128
rect 70302 119116 70308 119128
rect 67600 119088 70308 119116
rect 67600 119076 67606 119088
rect 70302 119076 70308 119088
rect 70360 119116 70366 119128
rect 75825 119119 75883 119125
rect 75825 119116 75837 119119
rect 70360 119088 75837 119116
rect 70360 119076 70366 119088
rect 75825 119085 75837 119088
rect 75871 119085 75883 119119
rect 75825 119079 75883 119085
rect 130930 118872 130936 118924
rect 130988 118912 130994 118924
rect 142246 118912 142252 118924
rect 130988 118884 142252 118912
rect 130988 118872 130994 118884
rect 142246 118872 142252 118884
rect 142304 118912 142310 118924
rect 142522 118912 142528 118924
rect 142304 118884 142528 118912
rect 142304 118872 142310 118884
rect 142522 118872 142528 118884
rect 142580 118872 142586 118924
rect 129642 118804 129648 118856
rect 129700 118844 129706 118856
rect 145098 118844 145104 118856
rect 129700 118816 145104 118844
rect 129700 118804 129706 118816
rect 145098 118804 145104 118816
rect 145156 118804 145162 118856
rect 131022 118736 131028 118788
rect 131080 118776 131086 118788
rect 147766 118776 147772 118788
rect 131080 118748 147772 118776
rect 131080 118736 131086 118748
rect 147766 118736 147772 118748
rect 147824 118736 147830 118788
rect 128722 118668 128728 118720
rect 128780 118708 128786 118720
rect 128906 118708 128912 118720
rect 128780 118680 128912 118708
rect 128780 118668 128786 118680
rect 128906 118668 128912 118680
rect 128964 118668 128970 118720
rect 129550 118668 129556 118720
rect 129608 118708 129614 118720
rect 149054 118708 149060 118720
rect 129608 118680 149060 118708
rect 129608 118668 129614 118680
rect 149054 118668 149060 118680
rect 149112 118668 149118 118720
rect 248233 118711 248291 118717
rect 248233 118677 248245 118711
rect 248279 118708 248291 118711
rect 248279 118680 248552 118708
rect 248279 118677 248291 118680
rect 248233 118671 248291 118677
rect 89717 118643 89775 118649
rect 89717 118609 89729 118643
rect 89763 118640 89775 118643
rect 99285 118643 99343 118649
rect 99285 118640 99297 118643
rect 89763 118612 99297 118640
rect 89763 118609 89775 118612
rect 89717 118603 89775 118609
rect 99285 118609 99297 118612
rect 99331 118609 99343 118643
rect 99285 118603 99343 118609
rect 104161 118643 104219 118649
rect 104161 118609 104173 118643
rect 104207 118640 104219 118643
rect 113821 118643 113879 118649
rect 113821 118640 113833 118643
rect 104207 118612 113833 118640
rect 104207 118609 104219 118612
rect 104161 118603 104219 118609
rect 113821 118609 113833 118612
rect 113867 118609 113879 118643
rect 113821 118603 113879 118609
rect 122745 118643 122803 118649
rect 122745 118609 122757 118643
rect 122791 118640 122803 118643
rect 168374 118640 168380 118652
rect 122791 118612 168380 118640
rect 122791 118609 122803 118612
rect 122745 118603 122803 118609
rect 168374 118600 168380 118612
rect 168432 118600 168438 118652
rect 178678 118600 178684 118652
rect 178736 118640 178742 118652
rect 216674 118640 216680 118652
rect 178736 118612 216680 118640
rect 178736 118600 178742 118612
rect 216674 118600 216680 118612
rect 216732 118600 216738 118652
rect 217318 118600 217324 118652
rect 217376 118640 217382 118652
rect 242250 118640 242256 118652
rect 217376 118612 242256 118640
rect 217376 118600 217382 118612
rect 242250 118600 242256 118612
rect 242308 118600 242314 118652
rect 244921 118643 244979 118649
rect 244921 118640 244933 118643
rect 242360 118612 244933 118640
rect 75914 118572 75920 118584
rect 75840 118544 75920 118572
rect 75840 118513 75868 118544
rect 75914 118532 75920 118544
rect 75972 118532 75978 118584
rect 97902 118532 97908 118584
rect 97960 118572 97966 118584
rect 181070 118572 181076 118584
rect 97960 118544 181076 118572
rect 97960 118532 97966 118544
rect 181070 118532 181076 118544
rect 181128 118532 181134 118584
rect 195882 118532 195888 118584
rect 195940 118572 195946 118584
rect 234614 118572 234620 118584
rect 195940 118544 234620 118572
rect 195940 118532 195946 118544
rect 234614 118532 234620 118544
rect 234672 118532 234678 118584
rect 238389 118575 238447 118581
rect 238389 118541 238401 118575
rect 238435 118572 238447 118575
rect 242360 118572 242388 118612
rect 244921 118609 244933 118612
rect 244967 118609 244979 118643
rect 244921 118603 244979 118609
rect 245841 118643 245899 118649
rect 245841 118609 245853 118643
rect 245887 118640 245899 118643
rect 248141 118643 248199 118649
rect 248141 118640 248153 118643
rect 245887 118612 248153 118640
rect 245887 118609 245899 118612
rect 245841 118603 245899 118609
rect 248141 118609 248153 118612
rect 248187 118609 248199 118643
rect 248524 118640 248552 118680
rect 428458 118668 428464 118720
rect 428516 118708 428522 118720
rect 433337 118711 433395 118717
rect 433337 118708 433349 118711
rect 428516 118680 433349 118708
rect 428516 118668 428522 118680
rect 433337 118677 433349 118680
rect 433383 118677 433395 118711
rect 433337 118671 433395 118677
rect 258258 118640 258264 118652
rect 248524 118612 258264 118640
rect 248141 118603 248199 118609
rect 258258 118600 258264 118612
rect 258316 118600 258322 118652
rect 306006 118600 306012 118652
rect 306064 118640 306070 118652
rect 332870 118640 332876 118652
rect 306064 118612 332876 118640
rect 306064 118600 306070 118612
rect 332870 118600 332876 118612
rect 332928 118600 332934 118652
rect 339586 118640 339592 118652
rect 333716 118612 339592 118640
rect 238435 118544 242388 118572
rect 242437 118575 242495 118581
rect 238435 118541 238447 118544
rect 238389 118535 238447 118541
rect 242437 118541 242449 118575
rect 242483 118572 242495 118575
rect 249153 118575 249211 118581
rect 242483 118544 249104 118572
rect 242483 118541 242495 118544
rect 242437 118535 242495 118541
rect 75825 118507 75883 118513
rect 75825 118473 75837 118507
rect 75871 118473 75883 118507
rect 75825 118467 75883 118473
rect 81345 118507 81403 118513
rect 81345 118473 81357 118507
rect 81391 118504 81403 118507
rect 82722 118504 82728 118516
rect 81391 118476 82728 118504
rect 81391 118473 81403 118476
rect 81345 118467 81403 118473
rect 82722 118464 82728 118476
rect 82780 118504 82786 118516
rect 164510 118504 164516 118516
rect 82780 118476 164516 118504
rect 82780 118464 82786 118476
rect 164510 118464 164516 118476
rect 164568 118464 164574 118516
rect 190362 118464 190368 118516
rect 190420 118504 190426 118516
rect 231302 118504 231308 118516
rect 190420 118476 231308 118504
rect 190420 118464 190426 118476
rect 231302 118464 231308 118476
rect 231360 118464 231366 118516
rect 239401 118507 239459 118513
rect 239401 118504 239413 118507
rect 231412 118476 239413 118504
rect 85482 118396 85488 118448
rect 85540 118436 85546 118448
rect 104161 118439 104219 118445
rect 104161 118436 104173 118439
rect 85540 118408 104173 118436
rect 85540 118396 85546 118408
rect 104161 118405 104173 118408
rect 104207 118405 104219 118439
rect 113082 118436 113088 118448
rect 104161 118399 104219 118405
rect 112456 118408 113088 118436
rect 71498 118328 71504 118380
rect 71556 118368 71562 118380
rect 88334 118368 88340 118380
rect 71556 118340 88340 118368
rect 71556 118328 71562 118340
rect 88334 118328 88340 118340
rect 88392 118328 88398 118380
rect 99285 118371 99343 118377
rect 99285 118337 99297 118371
rect 99331 118368 99343 118371
rect 112456 118368 112484 118408
rect 113082 118396 113088 118408
rect 113140 118396 113146 118448
rect 122653 118439 122711 118445
rect 122653 118405 122665 118439
rect 122699 118436 122711 118439
rect 175550 118436 175556 118448
rect 122699 118408 175556 118436
rect 122699 118405 122711 118408
rect 122653 118399 122711 118405
rect 175550 118396 175556 118408
rect 175608 118396 175614 118448
rect 186222 118396 186228 118448
rect 186280 118436 186286 118448
rect 229462 118436 229468 118448
rect 186280 118408 229468 118436
rect 186280 118396 186286 118408
rect 229462 118396 229468 118408
rect 229520 118396 229526 118448
rect 230382 118396 230388 118448
rect 230440 118436 230446 118448
rect 231412 118436 231440 118476
rect 239401 118473 239413 118476
rect 239447 118473 239459 118507
rect 239401 118467 239459 118473
rect 239493 118507 239551 118513
rect 239493 118473 239505 118507
rect 239539 118504 239551 118507
rect 240873 118507 240931 118513
rect 240873 118504 240885 118507
rect 239539 118476 240885 118504
rect 239539 118473 239551 118476
rect 239493 118467 239551 118473
rect 240873 118473 240885 118476
rect 240919 118473 240931 118507
rect 248969 118507 249027 118513
rect 248969 118504 248981 118507
rect 240873 118467 240931 118473
rect 240980 118476 248981 118504
rect 230440 118408 231440 118436
rect 231489 118439 231547 118445
rect 230440 118396 230446 118408
rect 231489 118405 231501 118439
rect 231535 118436 231547 118439
rect 236178 118436 236184 118448
rect 231535 118408 236184 118436
rect 231535 118405 231547 118408
rect 231489 118399 231547 118405
rect 236178 118396 236184 118408
rect 236236 118396 236242 118448
rect 238662 118396 238668 118448
rect 238720 118436 238726 118448
rect 240980 118436 241008 118476
rect 248969 118473 248981 118476
rect 249015 118473 249027 118507
rect 249076 118504 249104 118544
rect 249153 118541 249165 118575
rect 249199 118572 249211 118575
rect 252738 118572 252744 118584
rect 249199 118544 252744 118572
rect 249199 118541 249211 118544
rect 249153 118535 249211 118541
rect 252738 118532 252744 118544
rect 252796 118532 252802 118584
rect 252833 118575 252891 118581
rect 252833 118541 252845 118575
rect 252879 118572 252891 118575
rect 257614 118572 257620 118584
rect 252879 118544 257620 118572
rect 252879 118541 252891 118544
rect 252833 118535 252891 118541
rect 257614 118532 257620 118544
rect 257672 118532 257678 118584
rect 309686 118532 309692 118584
rect 309744 118572 309750 118584
rect 333716 118572 333744 118612
rect 339586 118600 339592 118612
rect 339644 118600 339650 118652
rect 345842 118600 345848 118652
rect 345900 118640 345906 118652
rect 396718 118640 396724 118652
rect 345900 118612 396724 118640
rect 345900 118600 345906 118612
rect 396718 118600 396724 118612
rect 396776 118600 396782 118652
rect 396813 118643 396871 118649
rect 396813 118609 396825 118643
rect 396859 118640 396871 118643
rect 398745 118643 398803 118649
rect 398745 118640 398757 118643
rect 396859 118612 398757 118640
rect 396859 118609 396871 118612
rect 396813 118603 396871 118609
rect 398745 118609 398757 118612
rect 398791 118609 398803 118643
rect 398745 118603 398803 118609
rect 400858 118600 400864 118652
rect 400916 118640 400922 118652
rect 480898 118640 480904 118652
rect 400916 118612 480904 118640
rect 400916 118600 400922 118612
rect 480898 118600 480904 118612
rect 480956 118600 480962 118652
rect 338390 118572 338396 118584
rect 309744 118544 333744 118572
rect 334728 118544 338396 118572
rect 309744 118532 309750 118544
rect 255314 118504 255320 118516
rect 249076 118476 255320 118504
rect 248969 118467 249027 118473
rect 255314 118464 255320 118476
rect 255372 118464 255378 118516
rect 257338 118464 257344 118516
rect 257396 118504 257402 118516
rect 264330 118504 264336 118516
rect 257396 118476 264336 118504
rect 257396 118464 257402 118476
rect 264330 118464 264336 118476
rect 264388 118464 264394 118516
rect 310882 118464 310888 118516
rect 310940 118504 310946 118516
rect 334529 118507 334587 118513
rect 334529 118504 334541 118507
rect 310940 118476 334541 118504
rect 310940 118464 310946 118476
rect 334529 118473 334541 118476
rect 334575 118473 334587 118507
rect 334529 118467 334587 118473
rect 238720 118408 241008 118436
rect 241057 118439 241115 118445
rect 238720 118396 238726 118408
rect 241057 118405 241069 118439
rect 241103 118436 241115 118439
rect 255774 118436 255780 118448
rect 241103 118408 255780 118436
rect 241103 118405 241115 118408
rect 241057 118399 241115 118405
rect 255774 118396 255780 118408
rect 255832 118396 255838 118448
rect 308490 118396 308496 118448
rect 308548 118436 308554 118448
rect 334728 118436 334756 118544
rect 338390 118532 338396 118544
rect 338448 118532 338454 118584
rect 362310 118532 362316 118584
rect 362368 118572 362374 118584
rect 442994 118572 443000 118584
rect 362368 118544 443000 118572
rect 362368 118532 362374 118544
rect 442994 118532 443000 118544
rect 443052 118532 443058 118584
rect 444377 118575 444435 118581
rect 444377 118541 444389 118575
rect 444423 118572 444435 118575
rect 456705 118575 456763 118581
rect 456705 118572 456717 118575
rect 444423 118544 456717 118572
rect 444423 118541 444435 118544
rect 444377 118535 444435 118541
rect 456705 118541 456717 118544
rect 456751 118541 456763 118575
rect 456705 118535 456763 118541
rect 334897 118507 334955 118513
rect 334897 118473 334909 118507
rect 334943 118504 334955 118507
rect 341334 118504 341340 118516
rect 334943 118476 341340 118504
rect 334943 118473 334955 118476
rect 334897 118467 334955 118473
rect 341334 118464 341340 118476
rect 341392 118464 341398 118516
rect 347590 118464 347596 118516
rect 347648 118504 347654 118516
rect 376018 118504 376024 118516
rect 347648 118476 376024 118504
rect 347648 118464 347654 118476
rect 376018 118464 376024 118476
rect 376076 118464 376082 118516
rect 393590 118464 393596 118516
rect 393648 118504 393654 118516
rect 475378 118504 475384 118516
rect 393648 118476 475384 118504
rect 393648 118464 393654 118476
rect 475378 118464 475384 118476
rect 475436 118464 475442 118516
rect 308548 118408 334756 118436
rect 308548 118396 308554 118408
rect 334802 118396 334808 118448
rect 334860 118436 334866 118448
rect 335262 118436 335268 118448
rect 334860 118408 335268 118436
rect 334860 118396 334866 118408
rect 335262 118396 335268 118408
rect 335320 118396 335326 118448
rect 342162 118396 342168 118448
rect 342220 118436 342226 118448
rect 389818 118436 389824 118448
rect 342220 118408 389824 118436
rect 342220 118396 342226 118408
rect 389818 118396 389824 118408
rect 389876 118396 389882 118448
rect 389913 118439 389971 118445
rect 389913 118405 389925 118439
rect 389959 118436 389971 118439
rect 396813 118439 396871 118445
rect 396813 118436 396825 118439
rect 389959 118408 396825 118436
rect 389959 118405 389971 118408
rect 389913 118399 389971 118405
rect 396813 118405 396825 118408
rect 396859 118405 396871 118439
rect 396813 118399 396871 118405
rect 397270 118396 397276 118448
rect 397328 118436 397334 118448
rect 478138 118436 478144 118448
rect 397328 118408 478144 118436
rect 397328 118396 397334 118408
rect 478138 118396 478144 118408
rect 478196 118396 478202 118448
rect 99331 118340 112484 118368
rect 112533 118371 112591 118377
rect 99331 118337 99343 118340
rect 99285 118331 99343 118337
rect 112533 118337 112545 118371
rect 112579 118368 112591 118371
rect 149882 118368 149888 118380
rect 112579 118340 149888 118368
rect 112579 118337 112591 118340
rect 112533 118331 112591 118337
rect 149882 118328 149888 118340
rect 149940 118328 149946 118380
rect 194502 118328 194508 118380
rect 194560 118368 194566 118380
rect 233234 118368 233240 118380
rect 194560 118340 233240 118368
rect 194560 118328 194566 118340
rect 233234 118328 233240 118340
rect 233292 118328 233298 118380
rect 234522 118328 234528 118380
rect 234580 118368 234586 118380
rect 253934 118368 253940 118380
rect 234580 118340 253940 118368
rect 234580 118328 234586 118340
rect 253934 118328 253940 118340
rect 253992 118328 253998 118380
rect 256602 118328 256608 118380
rect 256660 118368 256666 118380
rect 265526 118368 265532 118380
rect 256660 118340 265532 118368
rect 256660 118328 256666 118340
rect 265526 118328 265532 118340
rect 265584 118328 265590 118380
rect 311526 118328 311532 118380
rect 311584 118368 311590 118380
rect 343910 118368 343916 118380
rect 311584 118340 343916 118368
rect 311584 118328 311590 118340
rect 343910 118328 343916 118340
rect 343968 118328 343974 118380
rect 365990 118328 365996 118380
rect 366048 118368 366054 118380
rect 449894 118368 449900 118380
rect 366048 118340 449900 118368
rect 366048 118328 366054 118340
rect 449894 118328 449900 118340
rect 449952 118328 449958 118380
rect 71682 118260 71688 118312
rect 71740 118300 71746 118312
rect 73890 118300 73896 118312
rect 71740 118272 73896 118300
rect 71740 118260 71746 118272
rect 73890 118260 73896 118272
rect 73948 118260 73954 118312
rect 82630 118260 82636 118312
rect 82688 118300 82694 118312
rect 89717 118303 89775 118309
rect 89717 118300 89729 118303
rect 82688 118272 89729 118300
rect 82688 118260 82694 118272
rect 89717 118269 89729 118272
rect 89763 118269 89775 118303
rect 89717 118263 89775 118269
rect 113821 118303 113879 118309
rect 113821 118269 113833 118303
rect 113867 118300 113879 118303
rect 122745 118303 122803 118309
rect 122745 118300 122757 118303
rect 113867 118272 122757 118300
rect 113867 118269 113879 118272
rect 113821 118263 113879 118269
rect 122745 118269 122757 118272
rect 122791 118269 122803 118303
rect 125870 118300 125876 118312
rect 122745 118263 122803 118269
rect 125520 118272 125876 118300
rect 31662 118192 31668 118244
rect 31720 118232 31726 118244
rect 107562 118232 107568 118244
rect 31720 118204 107568 118232
rect 31720 118192 31726 118204
rect 107562 118192 107568 118204
rect 107620 118192 107626 118244
rect 108298 118192 108304 118244
rect 108356 118232 108362 118244
rect 125520 118232 125548 118272
rect 125870 118260 125876 118272
rect 125928 118300 125934 118312
rect 126882 118300 126888 118312
rect 125928 118272 126888 118300
rect 125928 118260 125934 118272
rect 126882 118260 126888 118272
rect 126940 118260 126946 118312
rect 129274 118260 129280 118312
rect 129332 118300 129338 118312
rect 182910 118300 182916 118312
rect 129332 118272 182916 118300
rect 129332 118260 129338 118272
rect 182910 118260 182916 118272
rect 182968 118260 182974 118312
rect 184842 118260 184848 118312
rect 184900 118300 184906 118312
rect 229186 118300 229192 118312
rect 184900 118272 229192 118300
rect 184900 118260 184906 118272
rect 229186 118260 229192 118272
rect 229244 118260 229250 118312
rect 231762 118260 231768 118312
rect 231820 118300 231826 118312
rect 244921 118303 244979 118309
rect 231820 118272 244872 118300
rect 231820 118260 231826 118272
rect 108356 118204 125548 118232
rect 108356 118192 108362 118204
rect 126238 118192 126244 118244
rect 126296 118232 126302 118244
rect 126974 118232 126980 118244
rect 126296 118204 126980 118232
rect 126296 118192 126302 118204
rect 126974 118192 126980 118204
rect 127032 118192 127038 118244
rect 129182 118192 129188 118244
rect 129240 118232 129246 118244
rect 177390 118232 177396 118244
rect 129240 118204 177396 118232
rect 129240 118192 129246 118204
rect 177390 118192 177396 118204
rect 177448 118192 177454 118244
rect 180058 118192 180064 118244
rect 180116 118232 180122 118244
rect 225138 118232 225144 118244
rect 180116 118204 225144 118232
rect 180116 118192 180122 118204
rect 225138 118192 225144 118204
rect 225196 118192 225202 118244
rect 225785 118235 225843 118241
rect 225785 118201 225797 118235
rect 225831 118232 225843 118235
rect 236822 118232 236828 118244
rect 225831 118204 236828 118232
rect 225831 118201 225843 118204
rect 225785 118195 225843 118201
rect 236822 118192 236828 118204
rect 236880 118192 236886 118244
rect 237190 118192 237196 118244
rect 237248 118232 237254 118244
rect 239309 118235 239367 118241
rect 239309 118232 239321 118235
rect 237248 118204 239321 118232
rect 237248 118192 237254 118204
rect 239309 118201 239321 118204
rect 239355 118201 239367 118235
rect 239309 118195 239367 118201
rect 239401 118235 239459 118241
rect 239401 118201 239413 118235
rect 239447 118232 239459 118235
rect 244737 118235 244795 118241
rect 244737 118232 244749 118235
rect 239447 118204 244749 118232
rect 239447 118201 239459 118204
rect 239401 118195 239459 118201
rect 244737 118201 244749 118204
rect 244783 118201 244795 118235
rect 244844 118232 244872 118272
rect 244921 118269 244933 118303
rect 244967 118300 244979 118303
rect 249794 118300 249800 118312
rect 244967 118272 249800 118300
rect 244967 118269 244979 118272
rect 244921 118263 244979 118269
rect 249794 118260 249800 118272
rect 249852 118260 249858 118312
rect 249889 118303 249947 118309
rect 249889 118269 249901 118303
rect 249935 118300 249947 118303
rect 251450 118300 251456 118312
rect 249935 118272 251456 118300
rect 249935 118269 249947 118272
rect 249889 118263 249947 118269
rect 251450 118260 251456 118272
rect 251508 118260 251514 118312
rect 251542 118260 251548 118312
rect 251600 118300 251606 118312
rect 256970 118300 256976 118312
rect 251600 118272 256976 118300
rect 251600 118260 251606 118272
rect 256970 118260 256976 118272
rect 257028 118260 257034 118312
rect 257982 118260 257988 118312
rect 258040 118300 258046 118312
rect 266354 118300 266360 118312
rect 258040 118272 266360 118300
rect 258040 118260 258046 118272
rect 266354 118260 266360 118272
rect 266412 118260 266418 118312
rect 296162 118260 296168 118312
rect 296220 118300 296226 118312
rect 305638 118300 305644 118312
rect 296220 118272 305644 118300
rect 296220 118260 296226 118272
rect 305638 118260 305644 118272
rect 305696 118260 305702 118312
rect 307202 118260 307208 118312
rect 307260 118300 307266 118312
rect 334618 118300 334624 118312
rect 307260 118272 334624 118300
rect 307260 118260 307266 118272
rect 334618 118260 334624 118272
rect 334676 118260 334682 118312
rect 336642 118260 336648 118312
rect 336700 118300 336706 118312
rect 374638 118300 374644 118312
rect 336700 118272 374644 118300
rect 336700 118260 336706 118272
rect 374638 118260 374644 118272
rect 374696 118260 374702 118312
rect 377030 118260 377036 118312
rect 377088 118300 377094 118312
rect 384301 118303 384359 118309
rect 384301 118300 384313 118303
rect 377088 118272 384313 118300
rect 377088 118260 377094 118272
rect 384301 118269 384313 118272
rect 384347 118269 384359 118303
rect 384301 118263 384359 118269
rect 398745 118303 398803 118309
rect 398745 118269 398757 118303
rect 398791 118300 398803 118303
rect 469858 118300 469864 118312
rect 398791 118272 469864 118300
rect 398791 118269 398803 118272
rect 398745 118263 398803 118269
rect 469858 118260 469864 118272
rect 469916 118260 469922 118312
rect 248877 118235 248935 118241
rect 248877 118232 248889 118235
rect 244844 118204 248889 118232
rect 244737 118195 244795 118201
rect 248877 118201 248889 118204
rect 248923 118201 248935 118235
rect 248877 118195 248935 118201
rect 254670 118192 254676 118244
rect 254728 118232 254734 118244
rect 263686 118232 263692 118244
rect 254728 118204 263692 118232
rect 254728 118192 254734 118204
rect 263686 118192 263692 118204
rect 263744 118192 263750 118244
rect 293770 118192 293776 118244
rect 293828 118232 293834 118244
rect 302878 118232 302884 118244
rect 293828 118204 302884 118232
rect 293828 118192 293834 118204
rect 302878 118192 302884 118204
rect 302936 118192 302942 118244
rect 307662 118192 307668 118244
rect 307720 118232 307726 118244
rect 336918 118232 336924 118244
rect 307720 118204 336924 118232
rect 307720 118192 307726 118204
rect 336918 118192 336924 118204
rect 336976 118192 336982 118244
rect 338482 118192 338488 118244
rect 338540 118232 338546 118244
rect 384206 118232 384212 118244
rect 338540 118204 384212 118232
rect 338540 118192 338546 118204
rect 384206 118192 384212 118204
rect 384264 118192 384270 118244
rect 386230 118192 386236 118244
rect 386288 118232 386294 118244
rect 389821 118235 389879 118241
rect 389821 118232 389833 118235
rect 386288 118204 389833 118232
rect 386288 118192 386294 118204
rect 389821 118201 389833 118204
rect 389867 118201 389879 118235
rect 389821 118195 389879 118201
rect 389910 118192 389916 118244
rect 389968 118232 389974 118244
rect 473998 118232 474004 118244
rect 389968 118204 474004 118232
rect 389968 118192 389974 118204
rect 473998 118192 474004 118204
rect 474056 118192 474062 118244
rect 28902 118124 28908 118176
rect 28960 118164 28966 118176
rect 111702 118164 111708 118176
rect 28960 118136 111708 118164
rect 28960 118124 28966 118136
rect 111702 118124 111708 118136
rect 111760 118124 111766 118176
rect 133233 118167 133291 118173
rect 126164 118136 133184 118164
rect 23382 118056 23388 118108
rect 23440 118096 23446 118108
rect 110322 118096 110328 118108
rect 23440 118068 110328 118096
rect 23440 118056 23446 118068
rect 110322 118056 110328 118068
rect 110380 118056 110386 118108
rect 113082 118056 113088 118108
rect 113140 118096 113146 118108
rect 122653 118099 122711 118105
rect 122653 118096 122665 118099
rect 113140 118068 122665 118096
rect 113140 118056 113146 118068
rect 122653 118065 122665 118068
rect 122699 118065 122711 118099
rect 122653 118059 122711 118065
rect 122745 118099 122803 118105
rect 122745 118065 122757 118099
rect 122791 118096 122803 118099
rect 125686 118096 125692 118108
rect 122791 118068 125692 118096
rect 122791 118065 122803 118068
rect 122745 118059 122803 118065
rect 125686 118056 125692 118068
rect 125744 118096 125750 118108
rect 126164 118096 126192 118136
rect 125744 118068 126192 118096
rect 125744 118056 125750 118068
rect 126974 118056 126980 118108
rect 127032 118096 127038 118108
rect 129553 118099 129611 118105
rect 129553 118096 129565 118099
rect 127032 118068 129565 118096
rect 127032 118056 127038 118068
rect 129553 118065 129565 118068
rect 129599 118065 129611 118099
rect 129553 118059 129611 118065
rect 129642 118056 129648 118108
rect 129700 118096 129706 118108
rect 133049 118099 133107 118105
rect 133049 118096 133061 118099
rect 129700 118068 133061 118096
rect 129700 118056 129706 118068
rect 133049 118065 133061 118068
rect 133095 118065 133107 118099
rect 133156 118096 133184 118136
rect 133233 118133 133245 118167
rect 133279 118164 133291 118167
rect 173894 118164 173900 118176
rect 133279 118136 173900 118164
rect 133279 118133 133291 118136
rect 133233 118127 133291 118133
rect 173894 118124 173900 118136
rect 173952 118124 173958 118176
rect 174538 118124 174544 118176
rect 174596 118164 174602 118176
rect 210421 118167 210479 118173
rect 210421 118164 210433 118167
rect 174596 118136 210433 118164
rect 174596 118124 174602 118136
rect 210421 118133 210433 118136
rect 210467 118133 210479 118167
rect 210421 118127 210479 118133
rect 220078 118124 220084 118176
rect 220136 118164 220142 118176
rect 238481 118167 238539 118173
rect 238481 118164 238493 118167
rect 220136 118136 238493 118164
rect 220136 118124 220142 118136
rect 238481 118133 238493 118136
rect 238527 118133 238539 118167
rect 249245 118167 249303 118173
rect 238481 118127 238539 118133
rect 239416 118136 247356 118164
rect 170030 118096 170036 118108
rect 133156 118068 170036 118096
rect 133049 118059 133107 118065
rect 170030 118056 170036 118068
rect 170088 118056 170094 118108
rect 179322 118056 179328 118108
rect 179380 118096 179386 118108
rect 225782 118096 225788 118108
rect 179380 118068 225788 118096
rect 179380 118056 179386 118068
rect 225782 118056 225788 118068
rect 225840 118056 225846 118108
rect 227622 118056 227628 118108
rect 227680 118096 227686 118108
rect 239416 118096 239444 118136
rect 227680 118068 239444 118096
rect 239493 118099 239551 118105
rect 227680 118056 227686 118068
rect 239493 118065 239505 118099
rect 239539 118096 239551 118099
rect 247218 118096 247224 118108
rect 239539 118068 247224 118096
rect 239539 118065 239551 118068
rect 239493 118059 239551 118065
rect 247218 118056 247224 118068
rect 247276 118056 247282 118108
rect 247328 118096 247356 118136
rect 249245 118133 249257 118167
rect 249291 118164 249303 118167
rect 250165 118167 250223 118173
rect 250165 118164 250177 118167
rect 249291 118136 250177 118164
rect 249291 118133 249303 118136
rect 249245 118127 249303 118133
rect 250165 118133 250177 118136
rect 250211 118133 250223 118167
rect 260006 118164 260012 118176
rect 250165 118127 250223 118133
rect 250364 118136 260012 118164
rect 250254 118096 250260 118108
rect 247328 118068 250260 118096
rect 250254 118056 250260 118068
rect 250312 118056 250318 118108
rect 60642 117988 60648 118040
rect 60700 118028 60706 118040
rect 81345 118031 81403 118037
rect 81345 118028 81357 118031
rect 60700 118000 81357 118028
rect 60700 117988 60706 118000
rect 81345 117997 81357 118000
rect 81391 117997 81403 118031
rect 81345 117991 81403 117997
rect 88334 117988 88340 118040
rect 88392 118028 88398 118040
rect 179414 118028 179420 118040
rect 88392 118000 179420 118028
rect 88392 117988 88398 118000
rect 179414 117988 179420 118000
rect 179472 117988 179478 118040
rect 183462 117988 183468 118040
rect 183520 118028 183526 118040
rect 227714 118028 227720 118040
rect 183520 118000 227720 118028
rect 183520 117988 183526 118000
rect 227714 117988 227720 118000
rect 227772 117988 227778 118040
rect 229002 117988 229008 118040
rect 229060 118028 229066 118040
rect 229060 118000 244688 118028
rect 229060 117988 229066 118000
rect 9582 117920 9588 117972
rect 9640 117960 9646 117972
rect 70210 117960 70216 117972
rect 9640 117932 70216 117960
rect 9640 117920 9646 117932
rect 70210 117920 70216 117932
rect 70268 117920 70274 117972
rect 73890 117920 73896 117972
rect 73948 117960 73954 117972
rect 75917 117963 75975 117969
rect 75917 117960 75929 117963
rect 73948 117932 75929 117960
rect 73948 117920 73954 117932
rect 75917 117929 75929 117932
rect 75963 117929 75975 117963
rect 75917 117923 75975 117929
rect 89717 117963 89775 117969
rect 89717 117929 89729 117963
rect 89763 117960 89775 117963
rect 96617 117963 96675 117969
rect 96617 117960 96629 117963
rect 89763 117932 96629 117960
rect 89763 117929 89775 117932
rect 89717 117923 89775 117929
rect 96617 117929 96629 117932
rect 96663 117929 96675 117963
rect 96617 117923 96675 117929
rect 107562 117920 107568 117972
rect 107620 117960 107626 117972
rect 112533 117963 112591 117969
rect 112533 117960 112545 117963
rect 107620 117932 112545 117960
rect 107620 117920 107626 117932
rect 112533 117929 112545 117932
rect 112579 117929 112591 117963
rect 112533 117923 112591 117929
rect 128906 117920 128912 117972
rect 128964 117960 128970 117972
rect 129642 117960 129648 117972
rect 128964 117932 129648 117960
rect 128964 117920 128970 117932
rect 129642 117920 129648 117932
rect 129700 117920 129706 117972
rect 132405 117963 132463 117969
rect 132405 117929 132417 117963
rect 132451 117960 132463 117963
rect 141973 117963 142031 117969
rect 141973 117960 141985 117963
rect 132451 117932 141985 117960
rect 132451 117929 132463 117932
rect 132405 117923 132463 117929
rect 141973 117929 141985 117932
rect 142019 117929 142031 117963
rect 141973 117923 142031 117929
rect 142154 117920 142160 117972
rect 142212 117960 142218 117972
rect 143074 117960 143080 117972
rect 142212 117932 143080 117960
rect 142212 117920 142218 117932
rect 143074 117920 143080 117932
rect 143132 117920 143138 117972
rect 156506 117920 156512 117972
rect 156564 117960 156570 117972
rect 156874 117960 156880 117972
rect 156564 117932 156880 117960
rect 156564 117920 156570 117932
rect 156874 117920 156880 117932
rect 156932 117920 156938 117972
rect 157245 117963 157303 117969
rect 157245 117929 157257 117963
rect 157291 117960 157303 117963
rect 171870 117960 171876 117972
rect 157291 117932 171876 117960
rect 157291 117929 157303 117932
rect 157245 117923 157303 117929
rect 171870 117920 171876 117932
rect 171928 117920 171934 117972
rect 176562 117920 176568 117972
rect 176620 117960 176626 117972
rect 223942 117960 223948 117972
rect 176620 117932 223948 117960
rect 176620 117920 176626 117932
rect 223942 117920 223948 117932
rect 224000 117920 224006 117972
rect 226242 117920 226248 117972
rect 226300 117960 226306 117972
rect 238389 117963 238447 117969
rect 238389 117960 238401 117963
rect 226300 117932 238401 117960
rect 226300 117920 226306 117932
rect 238389 117929 238401 117932
rect 238435 117929 238447 117963
rect 238389 117923 238447 117929
rect 238481 117963 238539 117969
rect 238481 117929 238493 117963
rect 238527 117960 238539 117963
rect 244274 117960 244280 117972
rect 238527 117932 244280 117960
rect 238527 117929 238539 117932
rect 238481 117923 238539 117929
rect 244274 117920 244280 117932
rect 244332 117920 244338 117972
rect 85485 117895 85543 117901
rect 85485 117861 85497 117895
rect 85531 117892 85543 117895
rect 85531 117864 89668 117892
rect 85531 117861 85543 117864
rect 85485 117855 85543 117861
rect 89640 117824 89668 117864
rect 122098 117852 122104 117904
rect 122156 117892 122162 117904
rect 122558 117892 122564 117904
rect 122156 117864 122564 117892
rect 122156 117852 122162 117864
rect 122558 117852 122564 117864
rect 122616 117892 122622 117904
rect 160830 117892 160836 117904
rect 122616 117864 160836 117892
rect 122616 117852 122622 117864
rect 160830 117852 160836 117864
rect 160888 117852 160894 117904
rect 197262 117852 197268 117904
rect 197320 117892 197326 117904
rect 234982 117892 234988 117904
rect 197320 117864 234988 117892
rect 197320 117852 197326 117864
rect 234982 117852 234988 117864
rect 235040 117852 235046 117904
rect 235350 117852 235356 117904
rect 235408 117892 235414 117904
rect 244553 117895 244611 117901
rect 244553 117892 244565 117895
rect 235408 117864 244565 117892
rect 235408 117852 235414 117864
rect 244553 117861 244565 117864
rect 244599 117861 244611 117895
rect 244660 117892 244688 118000
rect 245470 117988 245476 118040
rect 245528 118028 245534 118040
rect 250364 118028 250392 118136
rect 260006 118124 260012 118136
rect 260064 118124 260070 118176
rect 295610 118124 295616 118176
rect 295668 118164 295674 118176
rect 308398 118164 308404 118176
rect 295668 118136 308404 118164
rect 295668 118124 295674 118136
rect 308398 118124 308404 118136
rect 308456 118124 308462 118176
rect 320729 118167 320787 118173
rect 320729 118133 320741 118167
rect 320775 118164 320787 118167
rect 345106 118164 345112 118176
rect 320775 118136 345112 118164
rect 320775 118133 320787 118136
rect 320729 118127 320787 118133
rect 345106 118124 345112 118136
rect 345164 118124 345170 118176
rect 349430 118124 349436 118176
rect 349488 118164 349494 118176
rect 355321 118167 355379 118173
rect 355321 118164 355333 118167
rect 349488 118136 355333 118164
rect 349488 118124 349494 118136
rect 355321 118133 355333 118136
rect 355367 118133 355379 118167
rect 355321 118127 355379 118133
rect 369670 118124 369676 118176
rect 369728 118164 369734 118176
rect 456794 118164 456800 118176
rect 369728 118136 456800 118164
rect 369728 118124 369734 118136
rect 456794 118124 456800 118136
rect 456852 118124 456858 118176
rect 250441 118099 250499 118105
rect 250441 118065 250453 118099
rect 250487 118096 250499 118099
rect 250487 118068 252232 118096
rect 250487 118065 250499 118068
rect 250441 118059 250499 118065
rect 252094 118028 252100 118040
rect 245528 118000 250392 118028
rect 250456 118000 252100 118028
rect 245528 117988 245534 118000
rect 244737 117963 244795 117969
rect 244737 117929 244749 117963
rect 244783 117960 244795 117963
rect 250456 117960 250484 118000
rect 252094 117988 252100 118000
rect 252152 117988 252158 118040
rect 252204 118028 252232 118068
rect 252462 118056 252468 118108
rect 252520 118096 252526 118108
rect 263134 118096 263140 118108
rect 252520 118068 263140 118096
rect 252520 118056 252526 118068
rect 263134 118056 263140 118068
rect 263192 118056 263198 118108
rect 263410 118056 263416 118108
rect 263468 118096 263474 118108
rect 269206 118096 269212 118108
rect 263468 118068 269212 118096
rect 263468 118056 263474 118068
rect 269206 118056 269212 118068
rect 269264 118056 269270 118108
rect 284570 118056 284576 118108
rect 284628 118096 284634 118108
rect 291378 118096 291384 118108
rect 284628 118068 291384 118096
rect 284628 118056 284634 118068
rect 291378 118056 291384 118068
rect 291436 118056 291442 118108
rect 296622 118056 296628 118108
rect 296680 118096 296686 118108
rect 314838 118096 314844 118108
rect 296680 118068 314844 118096
rect 296680 118056 296686 118068
rect 314838 118056 314844 118068
rect 314896 118056 314902 118108
rect 324869 118099 324927 118105
rect 324869 118065 324881 118099
rect 324915 118096 324927 118099
rect 354306 118096 354312 118108
rect 324915 118068 354312 118096
rect 324915 118065 324927 118068
rect 324869 118059 324927 118065
rect 354306 118056 354312 118068
rect 354364 118056 354370 118108
rect 354401 118099 354459 118105
rect 354401 118065 354413 118099
rect 354447 118096 354459 118099
rect 369210 118096 369216 118108
rect 354447 118068 369216 118096
rect 354447 118065 354459 118068
rect 354401 118059 354459 118065
rect 369210 118056 369216 118068
rect 369268 118056 369274 118108
rect 373350 118056 373356 118108
rect 373408 118096 373414 118108
rect 463694 118096 463700 118108
rect 373408 118068 463700 118096
rect 373408 118056 373414 118068
rect 463694 118056 463700 118068
rect 463752 118056 463758 118108
rect 463789 118099 463847 118105
rect 463789 118065 463801 118099
rect 463835 118096 463847 118099
rect 476025 118099 476083 118105
rect 476025 118096 476037 118099
rect 463835 118068 476037 118096
rect 463835 118065 463847 118068
rect 463789 118059 463847 118065
rect 476025 118065 476037 118068
rect 476071 118065 476083 118099
rect 476025 118059 476083 118065
rect 252833 118031 252891 118037
rect 252833 118028 252845 118031
rect 252204 118000 252845 118028
rect 252833 117997 252845 118000
rect 252879 117997 252891 118031
rect 252833 117991 252891 117997
rect 255222 117988 255228 118040
rect 255280 118028 255286 118040
rect 264974 118028 264980 118040
rect 255280 118000 264980 118028
rect 255280 117988 255286 118000
rect 264974 117988 264980 118000
rect 265032 117988 265038 118040
rect 283926 117988 283932 118040
rect 283984 118028 283990 118040
rect 290090 118028 290096 118040
rect 283984 118000 290096 118028
rect 283984 117988 283990 118000
rect 290090 117988 290096 118000
rect 290148 117988 290154 118040
rect 298646 117988 298652 118040
rect 298704 118028 298710 118040
rect 318978 118028 318984 118040
rect 298704 118000 318984 118028
rect 298704 117988 298710 118000
rect 318978 117988 318984 118000
rect 319036 117988 319042 118040
rect 321922 117988 321928 118040
rect 321980 118028 321986 118040
rect 363506 118028 363512 118040
rect 321980 118000 363512 118028
rect 321980 117988 321986 118000
rect 363506 117988 363512 118000
rect 363564 117988 363570 118040
rect 384301 118031 384359 118037
rect 384301 117997 384313 118031
rect 384347 118028 384359 118031
rect 470594 118028 470600 118040
rect 384347 118000 470600 118028
rect 384347 117997 384359 118000
rect 384301 117991 384359 117997
rect 470594 117988 470600 118000
rect 470652 117988 470658 118040
rect 244783 117932 250484 117960
rect 244783 117929 244795 117932
rect 244737 117923 244795 117929
rect 251082 117920 251088 117972
rect 251140 117960 251146 117972
rect 262490 117960 262496 117972
rect 251140 117932 262496 117960
rect 251140 117920 251146 117932
rect 262490 117920 262496 117932
rect 262548 117920 262554 117972
rect 263502 117920 263508 117972
rect 263560 117960 263566 117972
rect 268654 117960 268660 117972
rect 263560 117932 268660 117960
rect 263560 117920 263566 117932
rect 268654 117920 268660 117932
rect 268712 117920 268718 117972
rect 294322 117920 294328 117972
rect 294380 117960 294386 117972
rect 295242 117960 295248 117972
rect 294380 117932 295248 117960
rect 294380 117920 294386 117932
rect 295242 117920 295248 117932
rect 295300 117920 295306 117972
rect 297450 117920 297456 117972
rect 297508 117960 297514 117972
rect 298002 117960 298008 117972
rect 297508 117932 298008 117960
rect 297508 117920 297514 117932
rect 298002 117920 298008 117932
rect 298060 117920 298066 117972
rect 300486 117920 300492 117972
rect 300544 117960 300550 117972
rect 321738 117960 321744 117972
rect 300544 117932 321744 117960
rect 300544 117920 300550 117932
rect 321738 117920 321744 117932
rect 321796 117920 321802 117972
rect 354306 117920 354312 117972
rect 354364 117960 354370 117972
rect 358170 117960 358176 117972
rect 354364 117932 358176 117960
rect 354364 117920 354370 117932
rect 358170 117920 358176 117932
rect 358228 117920 358234 117972
rect 380710 117920 380716 117972
rect 380768 117960 380774 117972
rect 477494 117960 477500 117972
rect 380768 117932 477500 117960
rect 380768 117920 380774 117932
rect 477494 117920 477500 117932
rect 477552 117920 477558 117972
rect 249153 117895 249211 117901
rect 244660 117864 249104 117892
rect 244553 117855 244611 117861
rect 89717 117827 89775 117833
rect 89717 117824 89729 117827
rect 89640 117796 89729 117824
rect 89717 117793 89729 117796
rect 89763 117793 89775 117827
rect 89717 117787 89775 117793
rect 96617 117827 96675 117833
rect 96617 117793 96629 117827
rect 96663 117824 96675 117827
rect 115845 117827 115903 117833
rect 96663 117796 99512 117824
rect 96663 117793 96675 117796
rect 96617 117787 96675 117793
rect 75917 117759 75975 117765
rect 75917 117725 75929 117759
rect 75963 117756 75975 117759
rect 85485 117759 85543 117765
rect 85485 117756 85497 117759
rect 75963 117728 85497 117756
rect 75963 117725 75975 117728
rect 75917 117719 75975 117725
rect 85485 117725 85497 117728
rect 85531 117725 85543 117759
rect 99484 117756 99512 117796
rect 115845 117793 115857 117827
rect 115891 117824 115903 117827
rect 117317 117827 117375 117833
rect 117317 117824 117329 117827
rect 115891 117796 117329 117824
rect 115891 117793 115903 117796
rect 115845 117787 115903 117793
rect 117317 117793 117329 117796
rect 117363 117793 117375 117827
rect 162854 117824 162860 117836
rect 117317 117787 117375 117793
rect 127728 117796 162860 117824
rect 106277 117759 106335 117765
rect 106277 117756 106289 117759
rect 99484 117728 106289 117756
rect 85485 117719 85543 117725
rect 106277 117725 106289 117728
rect 106323 117725 106335 117759
rect 106277 117719 106335 117725
rect 120718 117716 120724 117768
rect 120776 117756 120782 117768
rect 122745 117759 122803 117765
rect 122745 117756 122757 117759
rect 120776 117728 122757 117756
rect 120776 117716 120782 117728
rect 122745 117725 122757 117728
rect 122791 117725 122803 117759
rect 122745 117719 122803 117725
rect 126882 117716 126888 117768
rect 126940 117756 126946 117768
rect 127728 117756 127756 117796
rect 162854 117784 162860 117796
rect 162912 117784 162918 117836
rect 201402 117784 201408 117836
rect 201460 117824 201466 117836
rect 225785 117827 225843 117833
rect 225785 117824 225797 117827
rect 201460 117796 225797 117824
rect 201460 117784 201466 117796
rect 225785 117793 225797 117796
rect 225831 117793 225843 117827
rect 225785 117787 225843 117793
rect 233878 117784 233884 117836
rect 233936 117824 233942 117836
rect 238846 117824 238852 117836
rect 233936 117796 238852 117824
rect 233936 117784 233942 117796
rect 238846 117784 238852 117796
rect 238904 117784 238910 117836
rect 240042 117784 240048 117836
rect 240100 117824 240106 117836
rect 248966 117824 248972 117836
rect 240100 117796 248972 117824
rect 240100 117784 240106 117796
rect 248966 117784 248972 117796
rect 249024 117784 249030 117836
rect 249076 117824 249104 117864
rect 249153 117861 249165 117895
rect 249199 117892 249211 117895
rect 256694 117892 256700 117904
rect 249199 117864 256700 117892
rect 249199 117861 249211 117864
rect 249153 117855 249211 117861
rect 256694 117852 256700 117864
rect 256752 117852 256758 117904
rect 262122 117852 262128 117904
rect 262180 117892 262186 117904
rect 268010 117892 268016 117904
rect 262180 117864 268016 117892
rect 262180 117852 262186 117864
rect 268010 117852 268016 117864
rect 268068 117852 268074 117904
rect 288894 117852 288900 117904
rect 288952 117892 288958 117904
rect 288952 117864 293080 117892
rect 288952 117852 288958 117864
rect 251266 117824 251272 117836
rect 249076 117796 251272 117824
rect 251266 117784 251272 117796
rect 251324 117784 251330 117836
rect 293052 117824 293080 117864
rect 293126 117852 293132 117904
rect 293184 117892 293190 117904
rect 293862 117892 293868 117904
rect 293184 117864 293868 117892
rect 293184 117852 293190 117864
rect 293862 117852 293868 117864
rect 293920 117852 293926 117904
rect 304810 117852 304816 117904
rect 304868 117892 304874 117904
rect 304868 117864 311204 117892
rect 304868 117852 304874 117864
rect 297358 117824 297364 117836
rect 293052 117796 297364 117824
rect 297358 117784 297364 117796
rect 297416 117784 297422 117836
rect 311176 117824 311204 117864
rect 311802 117852 311808 117904
rect 311860 117892 311866 117904
rect 315485 117895 315543 117901
rect 315485 117892 315497 117895
rect 311860 117864 315497 117892
rect 311860 117852 311866 117864
rect 315485 117861 315497 117864
rect 315531 117861 315543 117895
rect 315485 117855 315543 117861
rect 315577 117895 315635 117901
rect 315577 117861 315589 117895
rect 315623 117892 315635 117895
rect 333974 117892 333980 117904
rect 315623 117864 333980 117892
rect 315623 117861 315635 117864
rect 315577 117855 315635 117861
rect 333974 117852 333980 117864
rect 334032 117852 334038 117904
rect 336737 117895 336795 117901
rect 336737 117861 336749 117895
rect 336783 117892 336795 117895
rect 350445 117895 350503 117901
rect 350445 117892 350457 117895
rect 336783 117864 350457 117892
rect 336783 117861 336795 117864
rect 336737 117855 336795 117861
rect 350445 117861 350457 117864
rect 350491 117861 350503 117895
rect 350445 117855 350503 117861
rect 353110 117852 353116 117904
rect 353168 117892 353174 117904
rect 425054 117892 425060 117904
rect 353168 117864 425060 117892
rect 353168 117852 353174 117864
rect 425054 117852 425060 117864
rect 425112 117852 425118 117904
rect 425146 117852 425152 117904
rect 425204 117892 425210 117904
rect 432601 117895 432659 117901
rect 432601 117892 432613 117895
rect 425204 117864 432613 117892
rect 425204 117852 425210 117864
rect 432601 117861 432613 117864
rect 432647 117861 432659 117895
rect 432601 117855 432659 117861
rect 432693 117895 432751 117901
rect 432693 117861 432705 117895
rect 432739 117892 432751 117895
rect 511258 117892 511264 117904
rect 432739 117864 511264 117892
rect 432739 117861 432751 117864
rect 432693 117855 432751 117861
rect 511258 117852 511264 117864
rect 511316 117852 511322 117904
rect 331306 117824 331312 117836
rect 311176 117796 331312 117824
rect 331306 117784 331312 117796
rect 331364 117784 331370 117836
rect 332962 117784 332968 117836
rect 333020 117824 333026 117836
rect 333882 117824 333888 117836
rect 333020 117796 333888 117824
rect 333020 117784 333026 117796
rect 333882 117784 333888 117796
rect 333940 117784 333946 117836
rect 350537 117827 350595 117833
rect 350537 117793 350549 117827
rect 350583 117824 350595 117827
rect 354401 117827 354459 117833
rect 354401 117824 354413 117827
rect 350583 117796 354413 117824
rect 350583 117793 350595 117796
rect 350537 117787 350595 117793
rect 354401 117793 354413 117796
rect 354447 117793 354459 117827
rect 354401 117787 354459 117793
rect 355321 117827 355379 117833
rect 355321 117793 355333 117827
rect 355367 117824 355379 117827
rect 416774 117824 416780 117836
rect 355367 117796 416780 117824
rect 355367 117793 355379 117796
rect 355321 117787 355379 117793
rect 416774 117784 416780 117796
rect 416832 117784 416838 117836
rect 419258 117784 419264 117836
rect 419316 117824 419322 117836
rect 420178 117824 420184 117836
rect 419316 117796 420184 117824
rect 419316 117784 419322 117796
rect 420178 117784 420184 117796
rect 420236 117784 420242 117836
rect 420733 117827 420791 117833
rect 420733 117793 420745 117827
rect 420779 117824 420791 117827
rect 422757 117827 422815 117833
rect 422757 117824 422769 117827
rect 420779 117796 422769 117824
rect 420779 117793 420791 117796
rect 420733 117787 420791 117793
rect 422757 117793 422769 117796
rect 422803 117793 422815 117827
rect 426437 117827 426495 117833
rect 426437 117824 426449 117827
rect 422757 117787 422815 117793
rect 422864 117796 426449 117824
rect 126940 117728 127756 117756
rect 126940 117716 126946 117728
rect 129090 117716 129096 117768
rect 129148 117756 129154 117768
rect 133233 117759 133291 117765
rect 133233 117756 133245 117759
rect 129148 117728 133245 117756
rect 129148 117716 129154 117728
rect 133233 117725 133245 117728
rect 133279 117725 133291 117759
rect 133233 117719 133291 117725
rect 133325 117759 133383 117765
rect 133325 117725 133337 117759
rect 133371 117756 133383 117759
rect 166350 117756 166356 117768
rect 133371 117728 166356 117756
rect 133371 117725 133383 117728
rect 133325 117719 133383 117725
rect 166350 117716 166356 117728
rect 166408 117716 166414 117768
rect 208302 117716 208308 117768
rect 208360 117756 208366 117768
rect 240410 117756 240416 117768
rect 208360 117728 240416 117756
rect 208360 117716 208366 117728
rect 240410 117716 240416 117728
rect 240468 117716 240474 117768
rect 240505 117759 240563 117765
rect 240505 117725 240517 117759
rect 240551 117756 240563 117759
rect 243538 117756 243544 117768
rect 240551 117728 243544 117756
rect 240551 117725 240563 117728
rect 240505 117719 240563 117725
rect 243538 117716 243544 117728
rect 243596 117716 243602 117768
rect 244182 117716 244188 117768
rect 244240 117756 244246 117768
rect 258810 117756 258816 117768
rect 244240 117728 258816 117756
rect 244240 117716 244246 117728
rect 258810 117716 258816 117728
rect 258868 117716 258874 117768
rect 302142 117716 302148 117768
rect 302200 117756 302206 117768
rect 325697 117759 325755 117765
rect 325697 117756 325709 117759
rect 302200 117728 325709 117756
rect 302200 117716 302206 117728
rect 325697 117725 325709 117728
rect 325743 117725 325755 117759
rect 325697 117719 325755 117725
rect 329282 117716 329288 117768
rect 329340 117756 329346 117768
rect 340785 117759 340843 117765
rect 340785 117756 340797 117759
rect 329340 117728 340797 117756
rect 329340 117716 329346 117728
rect 340785 117725 340797 117728
rect 340831 117725 340843 117759
rect 340785 117719 340843 117725
rect 340877 117759 340935 117765
rect 340877 117725 340889 117759
rect 340923 117756 340935 117759
rect 357986 117756 357992 117768
rect 340923 117728 357992 117756
rect 340923 117725 340935 117728
rect 340877 117719 340935 117725
rect 357986 117716 357992 117728
rect 358044 117716 358050 117768
rect 364058 117716 364064 117768
rect 364116 117756 364122 117768
rect 402238 117756 402244 117768
rect 364116 117728 402244 117756
rect 364116 117716 364122 117728
rect 402238 117716 402244 117728
rect 402296 117716 402302 117768
rect 411898 117716 411904 117768
rect 411956 117756 411962 117768
rect 413373 117759 413431 117765
rect 413373 117756 413385 117759
rect 411956 117728 413385 117756
rect 411956 117716 411962 117728
rect 413373 117725 413385 117728
rect 413419 117725 413431 117759
rect 413373 117719 413431 117725
rect 415302 117716 415308 117768
rect 415360 117756 415366 117768
rect 422864 117756 422892 117796
rect 426437 117793 426449 117796
rect 426483 117793 426495 117827
rect 426437 117787 426495 117793
rect 426529 117827 426587 117833
rect 426529 117793 426541 117827
rect 426575 117824 426587 117827
rect 500218 117824 500224 117836
rect 426575 117796 500224 117824
rect 426575 117793 426587 117796
rect 426529 117787 426587 117793
rect 500218 117784 500224 117796
rect 500276 117784 500282 117836
rect 415360 117728 422892 117756
rect 415360 117716 415366 117728
rect 422938 117716 422944 117768
rect 422996 117756 423002 117768
rect 424318 117756 424324 117768
rect 422996 117728 424324 117756
rect 422996 117716 423002 117728
rect 424318 117716 424324 117728
rect 424376 117716 424382 117768
rect 426342 117716 426348 117768
rect 426400 117756 426406 117768
rect 427817 117759 427875 117765
rect 427817 117756 427829 117759
rect 426400 117728 427829 117756
rect 426400 117716 426406 117728
rect 427817 117725 427829 117728
rect 427863 117725 427875 117759
rect 427817 117719 427875 117725
rect 433521 117759 433579 117765
rect 433521 117725 433533 117759
rect 433567 117756 433579 117759
rect 507118 117756 507124 117768
rect 433567 117728 507124 117756
rect 433567 117725 433579 117728
rect 433521 117719 433579 117725
rect 507118 117716 507124 117728
rect 507176 117716 507182 117768
rect 129553 117691 129611 117697
rect 129553 117657 129565 117691
rect 129599 117688 129611 117691
rect 157334 117688 157340 117700
rect 129599 117660 157340 117688
rect 129599 117657 129611 117660
rect 129553 117651 129611 117657
rect 157334 117648 157340 117660
rect 157392 117648 157398 117700
rect 185578 117648 185584 117700
rect 185636 117688 185642 117700
rect 209222 117688 209228 117700
rect 185636 117660 209228 117688
rect 185636 117648 185642 117660
rect 209222 117648 209228 117660
rect 209280 117648 209286 117700
rect 211062 117648 211068 117700
rect 211120 117688 211126 117700
rect 241698 117688 241704 117700
rect 211120 117660 241704 117688
rect 211120 117648 211126 117660
rect 241698 117648 241704 117660
rect 241756 117648 241762 117700
rect 245562 117648 245568 117700
rect 245620 117688 245626 117700
rect 259454 117688 259460 117700
rect 245620 117660 259460 117688
rect 245620 117648 245626 117660
rect 259454 117648 259460 117660
rect 259512 117648 259518 117700
rect 304166 117648 304172 117700
rect 304224 117688 304230 117700
rect 329834 117688 329840 117700
rect 304224 117660 329840 117688
rect 304224 117648 304230 117660
rect 329834 117648 329840 117660
rect 329892 117648 329898 117700
rect 336737 117691 336795 117697
rect 336737 117688 336749 117691
rect 329944 117660 336749 117688
rect 106277 117623 106335 117629
rect 106277 117589 106289 117623
rect 106323 117620 106335 117623
rect 115845 117623 115903 117629
rect 115845 117620 115857 117623
rect 106323 117592 115857 117620
rect 106323 117589 106335 117592
rect 106277 117583 106335 117589
rect 115845 117589 115857 117592
rect 115891 117589 115903 117623
rect 115845 117583 115903 117589
rect 130378 117580 130384 117632
rect 130436 117620 130442 117632
rect 158990 117620 158996 117632
rect 130436 117592 158996 117620
rect 130436 117580 130442 117592
rect 158990 117580 158996 117592
rect 159048 117580 159054 117632
rect 192478 117580 192484 117632
rect 192536 117620 192542 117632
rect 211154 117620 211160 117632
rect 192536 117592 211160 117620
rect 192536 117580 192542 117592
rect 211154 117580 211160 117592
rect 211212 117580 211218 117632
rect 213822 117580 213828 117632
rect 213880 117620 213886 117632
rect 235077 117623 235135 117629
rect 235077 117620 235089 117623
rect 213880 117592 235089 117620
rect 213880 117580 213886 117592
rect 235077 117589 235089 117592
rect 235123 117589 235135 117623
rect 235077 117583 235135 117589
rect 235169 117623 235227 117629
rect 235169 117589 235181 117623
rect 235215 117620 235227 117623
rect 238018 117620 238024 117632
rect 235215 117592 238024 117620
rect 235215 117589 235227 117592
rect 235169 117583 235227 117589
rect 238018 117580 238024 117592
rect 238076 117580 238082 117632
rect 238864 117592 246068 117620
rect 129458 117512 129464 117564
rect 129516 117552 129522 117564
rect 151998 117552 152004 117564
rect 129516 117524 152004 117552
rect 129516 117512 129522 117524
rect 151998 117512 152004 117524
rect 152056 117552 152062 117564
rect 155310 117552 155316 117564
rect 152056 117524 155316 117552
rect 152056 117512 152062 117524
rect 155310 117512 155316 117524
rect 155368 117512 155374 117564
rect 197998 117512 198004 117564
rect 198056 117552 198062 117564
rect 209958 117552 209964 117564
rect 198056 117524 209964 117552
rect 198056 117512 198062 117524
rect 209958 117512 209964 117524
rect 210016 117512 210022 117564
rect 210421 117555 210479 117561
rect 210421 117521 210433 117555
rect 210467 117552 210479 117555
rect 220262 117552 220268 117564
rect 210467 117524 220268 117552
rect 210467 117521 210479 117524
rect 210421 117515 210479 117521
rect 220262 117512 220268 117524
rect 220320 117512 220326 117564
rect 224218 117512 224224 117564
rect 224276 117552 224282 117564
rect 238757 117555 238815 117561
rect 238757 117552 238769 117555
rect 224276 117524 238769 117552
rect 224276 117512 224282 117524
rect 238757 117521 238769 117524
rect 238803 117521 238815 117555
rect 238757 117515 238815 117521
rect 129366 117444 129372 117496
rect 129424 117484 129430 117496
rect 135438 117484 135444 117496
rect 129424 117456 135444 117484
rect 129424 117444 129430 117456
rect 135438 117444 135444 117456
rect 135496 117484 135502 117496
rect 141878 117484 141884 117496
rect 135496 117456 141884 117484
rect 135496 117444 135502 117456
rect 141878 117444 141884 117456
rect 141936 117444 141942 117496
rect 141973 117487 142031 117493
rect 141973 117453 141985 117487
rect 142019 117484 142031 117487
rect 157245 117487 157303 117493
rect 157245 117484 157257 117487
rect 142019 117456 157257 117484
rect 142019 117453 142031 117456
rect 141973 117447 142031 117453
rect 157245 117453 157257 117456
rect 157291 117453 157303 117487
rect 157245 117447 157303 117453
rect 213178 117444 213184 117496
rect 213236 117484 213242 117496
rect 226978 117484 226984 117496
rect 213236 117456 226984 117484
rect 213236 117444 213242 117456
rect 226978 117444 226984 117456
rect 227036 117444 227042 117496
rect 228358 117444 228364 117496
rect 228416 117484 228422 117496
rect 238864 117484 238892 117592
rect 239585 117555 239643 117561
rect 239585 117521 239597 117555
rect 239631 117552 239643 117555
rect 242437 117555 242495 117561
rect 242437 117552 242449 117555
rect 239631 117524 242449 117552
rect 239631 117521 239643 117524
rect 239585 117515 239643 117521
rect 242437 117521 242449 117524
rect 242483 117521 242495 117555
rect 242437 117515 242495 117521
rect 243630 117512 243636 117564
rect 243688 117552 243694 117564
rect 245841 117555 245899 117561
rect 245841 117552 245853 117555
rect 243688 117524 245853 117552
rect 243688 117512 243694 117524
rect 245841 117521 245853 117524
rect 245887 117521 245899 117555
rect 246040 117552 246068 117592
rect 247678 117580 247684 117632
rect 247736 117620 247742 117632
rect 260834 117620 260840 117632
rect 247736 117592 260840 117620
rect 247736 117580 247742 117592
rect 260834 117580 260840 117592
rect 260892 117580 260898 117632
rect 294966 117580 294972 117632
rect 295024 117620 295030 117632
rect 311894 117620 311900 117632
rect 295024 117592 311900 117620
rect 295024 117580 295030 117592
rect 311894 117580 311900 117592
rect 311952 117580 311958 117632
rect 314562 117580 314568 117632
rect 314620 117620 314626 117632
rect 315485 117623 315543 117629
rect 314620 117592 315436 117620
rect 314620 117580 314626 117592
rect 247770 117552 247776 117564
rect 246040 117524 247776 117552
rect 245841 117515 245899 117521
rect 247770 117512 247776 117524
rect 247828 117512 247834 117564
rect 249245 117555 249303 117561
rect 249245 117552 249257 117555
rect 247880 117524 249257 117552
rect 228416 117456 238892 117484
rect 238941 117487 238999 117493
rect 228416 117444 228422 117456
rect 238941 117453 238953 117487
rect 238987 117484 238999 117487
rect 245930 117484 245936 117496
rect 238987 117456 245936 117484
rect 238987 117453 238999 117456
rect 238941 117447 238999 117453
rect 245930 117444 245936 117456
rect 245988 117444 245994 117496
rect 246025 117487 246083 117493
rect 246025 117453 246037 117487
rect 246071 117484 246083 117487
rect 247880 117484 247908 117524
rect 249245 117521 249257 117524
rect 249291 117521 249303 117555
rect 249245 117515 249303 117521
rect 249702 117512 249708 117564
rect 249760 117552 249766 117564
rect 262214 117552 262220 117564
rect 249760 117524 262220 117552
rect 249760 117512 249766 117524
rect 262214 117512 262220 117524
rect 262272 117512 262278 117564
rect 266262 117512 266268 117564
rect 266320 117552 266326 117564
rect 270494 117552 270500 117564
rect 266320 117524 270500 117552
rect 266320 117512 266326 117524
rect 270494 117512 270500 117524
rect 270552 117512 270558 117564
rect 280062 117512 280068 117564
rect 280120 117552 280126 117564
rect 283098 117552 283104 117564
rect 280120 117524 283104 117552
rect 280120 117512 280126 117524
rect 283098 117512 283104 117524
rect 283156 117512 283162 117564
rect 299842 117512 299848 117564
rect 299900 117552 299906 117564
rect 315298 117552 315304 117564
rect 299900 117524 315304 117552
rect 299900 117512 299906 117524
rect 315298 117512 315304 117524
rect 315356 117512 315362 117564
rect 315408 117552 315436 117592
rect 315485 117589 315497 117623
rect 315531 117620 315543 117623
rect 320729 117623 320787 117629
rect 320729 117620 320741 117623
rect 315531 117592 320741 117620
rect 315531 117589 315543 117592
rect 315485 117583 315543 117589
rect 320729 117589 320741 117592
rect 320775 117589 320787 117623
rect 320729 117583 320787 117589
rect 325418 117580 325424 117632
rect 325476 117620 325482 117632
rect 329944 117620 329972 117660
rect 336737 117657 336749 117660
rect 336783 117657 336795 117691
rect 336737 117651 336795 117657
rect 356790 117648 356796 117700
rect 356848 117688 356854 117700
rect 393958 117688 393964 117700
rect 356848 117660 393964 117688
rect 356848 117648 356854 117660
rect 393958 117648 393964 117660
rect 394016 117648 394022 117700
rect 404262 117648 404268 117700
rect 404320 117688 404326 117700
rect 482278 117688 482284 117700
rect 404320 117660 482284 117688
rect 404320 117648 404326 117660
rect 482278 117648 482284 117660
rect 482336 117648 482342 117700
rect 492585 117691 492643 117697
rect 492585 117657 492597 117691
rect 492631 117688 492643 117691
rect 492631 117660 492720 117688
rect 492631 117657 492643 117660
rect 492585 117651 492643 117657
rect 325476 117592 329972 117620
rect 325476 117580 325482 117592
rect 330478 117580 330484 117632
rect 330536 117620 330542 117632
rect 331030 117620 331036 117632
rect 330536 117592 331036 117620
rect 330536 117580 330542 117592
rect 331030 117580 331036 117592
rect 331088 117580 331094 117632
rect 354950 117580 354956 117632
rect 355008 117620 355014 117632
rect 355008 117592 358768 117620
rect 355008 117580 355014 117592
rect 320818 117552 320824 117564
rect 315408 117524 320824 117552
rect 320818 117512 320824 117524
rect 320876 117512 320882 117564
rect 358078 117512 358084 117564
rect 358136 117552 358142 117564
rect 358630 117552 358636 117564
rect 358136 117524 358636 117552
rect 358136 117512 358142 117524
rect 358630 117512 358636 117524
rect 358688 117512 358694 117564
rect 358740 117552 358768 117592
rect 359274 117580 359280 117632
rect 359332 117620 359338 117632
rect 360102 117620 360108 117632
rect 359332 117592 360108 117620
rect 359332 117580 359338 117592
rect 360102 117580 360108 117592
rect 360160 117580 360166 117632
rect 360470 117580 360476 117632
rect 360528 117620 360534 117632
rect 398098 117620 398104 117632
rect 360528 117592 398104 117620
rect 360528 117580 360534 117592
rect 398098 117580 398104 117592
rect 398156 117580 398162 117632
rect 408218 117580 408224 117632
rect 408276 117620 408282 117632
rect 486418 117620 486424 117632
rect 408276 117592 486424 117620
rect 408276 117580 408282 117592
rect 486418 117580 486424 117592
rect 486476 117580 486482 117632
rect 492692 117629 492720 117660
rect 492677 117623 492735 117629
rect 492677 117589 492689 117623
rect 492723 117589 492735 117623
rect 492677 117583 492735 117589
rect 369118 117552 369124 117564
rect 358740 117524 369124 117552
rect 369118 117512 369124 117524
rect 369176 117512 369182 117564
rect 384390 117512 384396 117564
rect 384448 117552 384454 117564
rect 413278 117552 413284 117564
rect 384448 117524 413284 117552
rect 384448 117512 384454 117524
rect 413278 117512 413284 117524
rect 413336 117512 413342 117564
rect 413373 117555 413431 117561
rect 413373 117521 413385 117555
rect 413419 117552 413431 117555
rect 413419 117524 416176 117552
rect 413419 117521 413431 117524
rect 413373 117515 413431 117521
rect 246071 117456 247908 117484
rect 246071 117453 246083 117456
rect 246025 117447 246083 117453
rect 248322 117444 248328 117496
rect 248380 117484 248386 117496
rect 261294 117484 261300 117496
rect 248380 117456 261300 117484
rect 248380 117444 248386 117456
rect 261294 117444 261300 117456
rect 261352 117444 261358 117496
rect 267642 117444 267648 117496
rect 267700 117484 267706 117496
rect 271046 117484 271052 117496
rect 267700 117456 271052 117484
rect 267700 117444 267706 117456
rect 271046 117444 271052 117456
rect 271104 117444 271110 117496
rect 282730 117444 282736 117496
rect 282788 117484 282794 117496
rect 284938 117484 284944 117496
rect 282788 117456 284944 117484
rect 282788 117444 282794 117456
rect 284938 117444 284944 117456
rect 284996 117444 285002 117496
rect 289446 117444 289452 117496
rect 289504 117484 289510 117496
rect 294598 117484 294604 117496
rect 289504 117456 294604 117484
rect 289504 117444 289510 117456
rect 294598 117444 294604 117456
rect 294656 117444 294662 117496
rect 306650 117444 306656 117496
rect 306708 117484 306714 117496
rect 315577 117487 315635 117493
rect 315577 117484 315589 117487
rect 306708 117456 315589 117484
rect 306708 117444 306714 117456
rect 315577 117453 315589 117456
rect 315623 117453 315635 117487
rect 315577 117447 315635 117453
rect 320082 117444 320088 117496
rect 320140 117484 320146 117496
rect 324869 117487 324927 117493
rect 324869 117484 324881 117487
rect 320140 117456 324881 117484
rect 320140 117444 320146 117456
rect 324869 117453 324881 117456
rect 324915 117453 324927 117487
rect 324869 117447 324927 117453
rect 324958 117444 324964 117496
rect 325016 117484 325022 117496
rect 326338 117484 326344 117496
rect 325016 117456 326344 117484
rect 325016 117444 325022 117456
rect 326338 117444 326344 117456
rect 326396 117444 326402 117496
rect 328086 117444 328092 117496
rect 328144 117484 328150 117496
rect 328270 117484 328276 117496
rect 328144 117456 328276 117484
rect 328144 117444 328150 117456
rect 328270 117444 328276 117456
rect 328328 117444 328334 117496
rect 367830 117444 367836 117496
rect 367888 117484 367894 117496
rect 377398 117484 377404 117496
rect 367888 117456 377404 117484
rect 367888 117444 367894 117456
rect 377398 117444 377404 117456
rect 377456 117444 377462 117496
rect 399662 117444 399668 117496
rect 399720 117484 399726 117496
rect 400030 117484 400036 117496
rect 399720 117456 400036 117484
rect 399720 117444 399726 117456
rect 400030 117444 400036 117456
rect 400088 117444 400094 117496
rect 408862 117444 408868 117496
rect 408920 117484 408926 117496
rect 409690 117484 409696 117496
rect 408920 117456 409696 117484
rect 408920 117444 408926 117456
rect 409690 117444 409696 117456
rect 409748 117444 409754 117496
rect 111702 117376 111708 117428
rect 111760 117416 111766 117428
rect 148042 117416 148048 117428
rect 111760 117388 148048 117416
rect 111760 117376 111766 117388
rect 148042 117376 148048 117388
rect 148100 117376 148106 117428
rect 229738 117376 229744 117428
rect 229796 117416 229802 117428
rect 235169 117419 235227 117425
rect 235169 117416 235181 117419
rect 229796 117388 235181 117416
rect 229796 117376 229802 117388
rect 235169 117385 235181 117388
rect 235215 117385 235227 117419
rect 235169 117379 235227 117385
rect 235258 117376 235264 117428
rect 235316 117416 235322 117428
rect 244553 117419 244611 117425
rect 235316 117388 244504 117416
rect 235316 117376 235322 117388
rect 92382 117308 92388 117360
rect 92440 117348 92446 117360
rect 97902 117348 97908 117360
rect 92440 117320 97908 117348
rect 92440 117308 92446 117320
rect 97902 117308 97908 117320
rect 97960 117308 97966 117360
rect 117317 117351 117375 117357
rect 117317 117317 117329 117351
rect 117363 117348 117375 117351
rect 132405 117351 132463 117357
rect 132405 117348 132417 117351
rect 117363 117320 132417 117348
rect 117363 117317 117375 117320
rect 117317 117311 117375 117317
rect 132405 117317 132417 117320
rect 132451 117317 132463 117351
rect 132405 117311 132463 117317
rect 132681 117351 132739 117357
rect 132681 117317 132693 117351
rect 132727 117348 132739 117351
rect 133049 117351 133107 117357
rect 133049 117348 133061 117351
rect 132727 117320 133061 117348
rect 132727 117317 132739 117320
rect 132681 117311 132739 117317
rect 133049 117317 133061 117320
rect 133095 117348 133107 117351
rect 190270 117348 190276 117360
rect 133095 117320 190276 117348
rect 133095 117317 133107 117320
rect 133049 117311 133107 117317
rect 190270 117308 190276 117320
rect 190328 117308 190334 117360
rect 190546 117308 190552 117360
rect 190604 117348 190610 117360
rect 195974 117348 195980 117360
rect 190604 117320 195980 117348
rect 190604 117308 190610 117320
rect 195974 117308 195980 117320
rect 196032 117308 196038 117360
rect 225598 117308 225604 117360
rect 225656 117348 225662 117360
rect 231489 117351 231547 117357
rect 231489 117348 231501 117351
rect 225656 117320 231501 117348
rect 225656 117308 225662 117320
rect 231489 117317 231501 117320
rect 231535 117317 231547 117351
rect 231489 117311 231547 117317
rect 232406 117308 232412 117360
rect 232464 117348 232470 117360
rect 239493 117351 239551 117357
rect 239493 117348 239505 117351
rect 232464 117320 239505 117348
rect 232464 117308 232470 117320
rect 239493 117317 239505 117320
rect 239539 117317 239551 117351
rect 239493 117311 239551 117317
rect 239585 117351 239643 117357
rect 239585 117317 239597 117351
rect 239631 117317 239643 117351
rect 240505 117351 240563 117357
rect 240505 117348 240517 117351
rect 239585 117311 239643 117317
rect 239692 117320 240517 117348
rect 132954 117240 132960 117292
rect 133012 117280 133018 117292
rect 186133 117283 186191 117289
rect 186133 117280 186145 117283
rect 133012 117252 186145 117280
rect 133012 117240 133018 117252
rect 186133 117249 186145 117252
rect 186179 117249 186191 117283
rect 186133 117243 186191 117249
rect 237282 117240 237288 117292
rect 237340 117280 237346 117292
rect 239600 117280 239628 117311
rect 237340 117252 239628 117280
rect 237340 117240 237346 117252
rect 161385 117215 161443 117221
rect 161385 117181 161397 117215
rect 161431 117212 161443 117215
rect 235077 117215 235135 117221
rect 161431 117184 164096 117212
rect 161431 117181 161443 117184
rect 161385 117175 161443 117181
rect 138845 117147 138903 117153
rect 138845 117113 138857 117147
rect 138891 117144 138903 117147
rect 143537 117147 143595 117153
rect 143537 117144 143549 117147
rect 138891 117116 143549 117144
rect 138891 117113 138903 117116
rect 138845 117107 138903 117113
rect 143537 117113 143549 117116
rect 143583 117113 143595 117147
rect 143537 117107 143595 117113
rect 151817 117147 151875 117153
rect 151817 117113 151829 117147
rect 151863 117144 151875 117147
rect 161293 117147 161351 117153
rect 161293 117144 161305 117147
rect 151863 117116 161305 117144
rect 151863 117113 151875 117116
rect 151817 117107 151875 117113
rect 161293 117113 161305 117116
rect 161339 117113 161351 117147
rect 161293 117107 161351 117113
rect 164068 117076 164096 117184
rect 171152 117184 180748 117212
rect 171152 117144 171180 117184
rect 167656 117116 171180 117144
rect 180720 117144 180748 117184
rect 235077 117181 235089 117215
rect 235123 117212 235135 117215
rect 239692 117212 239720 117320
rect 240505 117317 240517 117320
rect 240551 117317 240563 117351
rect 240505 117311 240563 117317
rect 241422 117308 241428 117360
rect 241480 117348 241486 117360
rect 244476 117348 244504 117388
rect 244553 117385 244565 117419
rect 244599 117416 244611 117419
rect 253290 117416 253296 117428
rect 244599 117388 253296 117416
rect 244599 117385 244611 117388
rect 244553 117379 244611 117385
rect 253290 117376 253296 117388
rect 253348 117376 253354 117428
rect 261478 117376 261484 117428
rect 261536 117416 261542 117428
rect 267734 117416 267740 117428
rect 261536 117388 267740 117416
rect 261536 117376 261542 117388
rect 267734 117376 267740 117388
rect 267792 117376 267798 117428
rect 269758 117376 269764 117428
rect 269816 117416 269822 117428
rect 271874 117416 271880 117428
rect 269816 117388 271880 117416
rect 269816 117376 269822 117388
rect 271874 117376 271880 117388
rect 271932 117376 271938 117428
rect 272518 117376 272524 117428
rect 272576 117416 272582 117428
rect 273530 117416 273536 117428
rect 272576 117388 273536 117416
rect 272576 117376 272582 117388
rect 273530 117376 273536 117388
rect 273588 117376 273594 117428
rect 278406 117376 278412 117428
rect 278464 117416 278470 117428
rect 279142 117416 279148 117428
rect 278464 117388 279148 117416
rect 278464 117376 278470 117388
rect 279142 117376 279148 117388
rect 279200 117376 279206 117428
rect 282086 117376 282092 117428
rect 282144 117416 282150 117428
rect 283558 117416 283564 117428
rect 282144 117388 283564 117416
rect 282144 117376 282150 117388
rect 283558 117376 283564 117388
rect 283616 117376 283622 117428
rect 289998 117376 290004 117428
rect 290056 117416 290062 117428
rect 291102 117416 291108 117428
rect 290056 117388 291108 117416
rect 290056 117376 290062 117388
rect 291102 117376 291108 117388
rect 291160 117376 291166 117428
rect 316402 117376 316408 117428
rect 316460 117416 316466 117428
rect 317322 117416 317328 117428
rect 316460 117388 317328 117416
rect 316460 117376 316466 117388
rect 317322 117376 317328 117388
rect 317380 117376 317386 117428
rect 318242 117376 318248 117428
rect 318300 117416 318306 117428
rect 322198 117416 322204 117428
rect 318300 117388 322204 117416
rect 318300 117376 318306 117388
rect 322198 117376 322204 117388
rect 322256 117376 322262 117428
rect 344002 117376 344008 117428
rect 344060 117416 344066 117428
rect 344922 117416 344928 117428
rect 344060 117388 344928 117416
rect 344060 117376 344066 117388
rect 344922 117376 344928 117388
rect 344980 117376 344986 117428
rect 371510 117376 371516 117428
rect 371568 117416 371574 117428
rect 372522 117416 372528 117428
rect 371568 117388 372528 117416
rect 371568 117376 371574 117388
rect 372522 117376 372528 117388
rect 372580 117376 372586 117428
rect 405182 117376 405188 117428
rect 405240 117416 405246 117428
rect 405642 117416 405648 117428
rect 405240 117388 405648 117416
rect 405240 117376 405246 117388
rect 405642 117376 405648 117388
rect 405700 117376 405706 117428
rect 410702 117376 410708 117428
rect 410760 117416 410766 117428
rect 411162 117416 411168 117428
rect 410760 117388 411168 117416
rect 410760 117376 410766 117388
rect 411162 117376 411168 117388
rect 411220 117376 411226 117428
rect 413738 117376 413744 117428
rect 413796 117416 413802 117428
rect 416038 117416 416044 117428
rect 413796 117388 416044 117416
rect 413796 117376 413802 117388
rect 416038 117376 416044 117388
rect 416096 117376 416102 117428
rect 249889 117351 249947 117357
rect 249889 117348 249901 117351
rect 241480 117320 244412 117348
rect 244476 117320 249901 117348
rect 241480 117308 241486 117320
rect 244384 117280 244412 117320
rect 249889 117317 249901 117320
rect 249935 117317 249947 117351
rect 249889 117311 249947 117317
rect 250438 117308 250444 117360
rect 250496 117348 250502 117360
rect 254578 117348 254584 117360
rect 250496 117320 254584 117348
rect 250496 117308 250502 117320
rect 254578 117308 254584 117320
rect 254636 117308 254642 117360
rect 259362 117308 259368 117360
rect 259420 117348 259426 117360
rect 266814 117348 266820 117360
rect 259420 117320 266820 117348
rect 259420 117308 259426 117320
rect 266814 117308 266820 117320
rect 266872 117308 266878 117360
rect 268378 117308 268384 117360
rect 268436 117348 268442 117360
rect 269850 117348 269856 117360
rect 268436 117320 269856 117348
rect 268436 117308 268442 117320
rect 269850 117308 269856 117320
rect 269908 117308 269914 117360
rect 273162 117308 273168 117360
rect 273220 117348 273226 117360
rect 274174 117348 274180 117360
rect 273220 117320 274180 117348
rect 273220 117308 273226 117320
rect 274174 117308 274180 117320
rect 274232 117308 274238 117360
rect 277854 117308 277860 117360
rect 277912 117348 277918 117360
rect 278866 117348 278872 117360
rect 277912 117320 278872 117348
rect 277912 117308 277918 117320
rect 278866 117308 278872 117320
rect 278924 117308 278930 117360
rect 279050 117308 279056 117360
rect 279108 117348 279114 117360
rect 280338 117348 280344 117360
rect 279108 117320 280344 117348
rect 279108 117308 279114 117320
rect 280338 117308 280344 117320
rect 280396 117308 280402 117360
rect 280890 117308 280896 117360
rect 280948 117348 280954 117360
rect 281350 117348 281356 117360
rect 280948 117320 281356 117348
rect 280948 117308 280954 117320
rect 281350 117308 281356 117320
rect 281408 117308 281414 117360
rect 283374 117308 283380 117360
rect 283432 117348 283438 117360
rect 284202 117348 284208 117360
rect 283432 117320 284208 117348
rect 283432 117308 283438 117320
rect 284202 117308 284208 117320
rect 284260 117308 284266 117360
rect 285214 117308 285220 117360
rect 285272 117348 285278 117360
rect 285582 117348 285588 117360
rect 285272 117320 285588 117348
rect 285272 117308 285278 117320
rect 285582 117308 285588 117320
rect 285640 117308 285646 117360
rect 286410 117308 286416 117360
rect 286468 117348 286474 117360
rect 286870 117348 286876 117360
rect 286468 117320 286876 117348
rect 286468 117308 286474 117320
rect 286870 117308 286876 117320
rect 286928 117308 286934 117360
rect 287606 117308 287612 117360
rect 287664 117348 287670 117360
rect 288342 117348 288348 117360
rect 287664 117320 288348 117348
rect 287664 117308 287670 117320
rect 288342 117308 288348 117320
rect 288400 117308 288406 117360
rect 290734 117308 290740 117360
rect 290792 117348 290798 117360
rect 291010 117348 291016 117360
rect 290792 117320 291016 117348
rect 290792 117308 290798 117320
rect 291010 117308 291016 117320
rect 291068 117308 291074 117360
rect 291930 117308 291936 117360
rect 291988 117348 291994 117360
rect 292482 117348 292488 117360
rect 291988 117320 292488 117348
rect 291988 117308 291994 117320
rect 292482 117308 292488 117320
rect 292540 117308 292546 117360
rect 301130 117308 301136 117360
rect 301188 117348 301194 117360
rect 302142 117348 302148 117360
rect 301188 117320 302148 117348
rect 301188 117308 301194 117320
rect 302142 117308 302148 117320
rect 302200 117308 302206 117360
rect 302970 117308 302976 117360
rect 303028 117348 303034 117360
rect 303522 117348 303528 117360
rect 303028 117320 303528 117348
rect 303028 117308 303034 117320
rect 303522 117308 303528 117320
rect 303580 117308 303586 117360
rect 305362 117308 305368 117360
rect 305420 117348 305426 117360
rect 306282 117348 306288 117360
rect 305420 117320 306288 117348
rect 305420 117308 305426 117320
rect 306282 117308 306288 117320
rect 306340 117308 306346 117360
rect 312722 117308 312728 117360
rect 312780 117348 312786 117360
rect 313182 117348 313188 117360
rect 312780 117320 313188 117348
rect 312780 117308 312786 117320
rect 313182 117308 313188 117320
rect 313240 117308 313246 117360
rect 313918 117308 313924 117360
rect 313976 117348 313982 117360
rect 314562 117348 314568 117360
rect 313976 117320 314568 117348
rect 313976 117308 313982 117320
rect 314562 117308 314568 117320
rect 314620 117308 314626 117360
rect 315206 117308 315212 117360
rect 315264 117348 315270 117360
rect 315850 117348 315856 117360
rect 315264 117320 315856 117348
rect 315264 117308 315270 117320
rect 315850 117308 315856 117320
rect 315908 117308 315914 117360
rect 317046 117308 317052 117360
rect 317104 117348 317110 117360
rect 317230 117348 317236 117360
rect 317104 117320 317236 117348
rect 317104 117308 317110 117320
rect 317230 117308 317236 117320
rect 317288 117308 317294 117360
rect 319438 117308 319444 117360
rect 319496 117348 319502 117360
rect 320082 117348 320088 117360
rect 319496 117320 320088 117348
rect 319496 117308 319502 117320
rect 320082 117308 320088 117320
rect 320140 117308 320146 117360
rect 320726 117308 320732 117360
rect 320784 117348 320790 117360
rect 321370 117348 321376 117360
rect 320784 117320 321376 117348
rect 320784 117308 320790 117320
rect 321370 117308 321376 117320
rect 321428 117308 321434 117360
rect 323762 117308 323768 117360
rect 323820 117348 323826 117360
rect 324222 117348 324228 117360
rect 323820 117320 324228 117348
rect 323820 117308 323826 117320
rect 324222 117308 324228 117320
rect 324280 117308 324286 117360
rect 326246 117308 326252 117360
rect 326304 117348 326310 117360
rect 326982 117348 326988 117360
rect 326304 117320 326988 117348
rect 326304 117308 326310 117320
rect 326982 117308 326988 117320
rect 327040 117308 327046 117360
rect 327442 117308 327448 117360
rect 327500 117348 327506 117360
rect 328362 117348 328368 117360
rect 327500 117320 328368 117348
rect 327500 117308 327506 117320
rect 328362 117308 328368 117320
rect 328420 117308 328426 117360
rect 331674 117308 331680 117360
rect 331732 117348 331738 117360
rect 332502 117348 332508 117360
rect 331732 117320 332508 117348
rect 331732 117308 331738 117320
rect 332502 117308 332508 117320
rect 332560 117308 332566 117360
rect 333514 117308 333520 117360
rect 333572 117348 333578 117360
rect 333790 117348 333796 117360
rect 333572 117320 333796 117348
rect 333572 117308 333578 117320
rect 333790 117308 333796 117320
rect 333848 117308 333854 117360
rect 335998 117308 336004 117360
rect 336056 117348 336062 117360
rect 336642 117348 336648 117360
rect 336056 117320 336648 117348
rect 336056 117308 336062 117320
rect 336642 117308 336648 117320
rect 336700 117308 336706 117360
rect 337194 117308 337200 117360
rect 337252 117348 337258 117360
rect 338022 117348 338028 117360
rect 337252 117320 338028 117348
rect 337252 117308 337258 117320
rect 338022 117308 338028 117320
rect 338080 117308 338086 117360
rect 339034 117308 339040 117360
rect 339092 117348 339098 117360
rect 339402 117348 339408 117360
rect 339092 117320 339408 117348
rect 339092 117308 339098 117320
rect 339402 117308 339408 117320
rect 339460 117308 339466 117360
rect 340322 117308 340328 117360
rect 340380 117348 340386 117360
rect 340782 117348 340788 117360
rect 340380 117320 340788 117348
rect 340380 117308 340386 117320
rect 340782 117308 340788 117320
rect 340840 117308 340846 117360
rect 341518 117308 341524 117360
rect 341576 117348 341582 117360
rect 342162 117348 342168 117360
rect 341576 117320 342168 117348
rect 341576 117308 341582 117320
rect 342162 117308 342168 117320
rect 342220 117308 342226 117360
rect 342714 117308 342720 117360
rect 342772 117348 342778 117360
rect 343542 117348 343548 117360
rect 342772 117320 343548 117348
rect 342772 117308 342778 117320
rect 343542 117308 343548 117320
rect 343600 117308 343606 117360
rect 344554 117308 344560 117360
rect 344612 117348 344618 117360
rect 344830 117348 344836 117360
rect 344612 117320 344836 117348
rect 344612 117308 344618 117320
rect 344830 117308 344836 117320
rect 344888 117308 344894 117360
rect 347038 117308 347044 117360
rect 347096 117348 347102 117360
rect 347682 117348 347688 117360
rect 347096 117320 347688 117348
rect 347096 117308 347102 117320
rect 347682 117308 347688 117320
rect 347740 117308 347746 117360
rect 348234 117308 348240 117360
rect 348292 117348 348298 117360
rect 349062 117348 349068 117360
rect 348292 117320 349068 117348
rect 348292 117308 348298 117320
rect 349062 117308 349068 117320
rect 349120 117308 349126 117360
rect 350074 117308 350080 117360
rect 350132 117348 350138 117360
rect 350442 117348 350448 117360
rect 350132 117320 350448 117348
rect 350132 117308 350138 117320
rect 350442 117308 350448 117320
rect 350500 117308 350506 117360
rect 351270 117308 351276 117360
rect 351328 117348 351334 117360
rect 351822 117348 351828 117360
rect 351328 117320 351828 117348
rect 351328 117308 351334 117320
rect 351822 117308 351828 117320
rect 351880 117308 351886 117360
rect 352558 117308 352564 117360
rect 352616 117348 352622 117360
rect 353202 117348 353208 117360
rect 352616 117320 353208 117348
rect 352616 117308 352622 117320
rect 353202 117308 353208 117320
rect 353260 117308 353266 117360
rect 353754 117308 353760 117360
rect 353812 117348 353818 117360
rect 354582 117348 354588 117360
rect 353812 117320 354588 117348
rect 353812 117308 353818 117320
rect 354582 117308 354588 117320
rect 354640 117308 354646 117360
rect 355594 117308 355600 117360
rect 355652 117348 355658 117360
rect 355962 117348 355968 117360
rect 355652 117320 355968 117348
rect 355652 117308 355658 117320
rect 355962 117308 355968 117320
rect 356020 117308 356026 117360
rect 361114 117308 361120 117360
rect 361172 117348 361178 117360
rect 361482 117348 361488 117360
rect 361172 117320 361488 117348
rect 361172 117308 361178 117320
rect 361482 117308 361488 117320
rect 361540 117308 361546 117360
rect 363598 117308 363604 117360
rect 363656 117348 363662 117360
rect 364242 117348 364248 117360
rect 363656 117320 364248 117348
rect 363656 117308 363662 117320
rect 364242 117308 364248 117320
rect 364300 117308 364306 117360
rect 364794 117308 364800 117360
rect 364852 117348 364858 117360
rect 365622 117348 365628 117360
rect 364852 117320 365628 117348
rect 364852 117308 364858 117320
rect 365622 117308 365628 117320
rect 365680 117308 365686 117360
rect 366634 117308 366640 117360
rect 366692 117348 366698 117360
rect 367002 117348 367008 117360
rect 366692 117320 367008 117348
rect 366692 117308 366698 117320
rect 367002 117308 367008 117320
rect 367060 117308 367066 117360
rect 369026 117308 369032 117360
rect 369084 117348 369090 117360
rect 369762 117348 369768 117360
rect 369084 117320 369768 117348
rect 369084 117308 369090 117320
rect 369762 117308 369768 117320
rect 369820 117308 369826 117360
rect 370314 117308 370320 117360
rect 370372 117348 370378 117360
rect 371142 117348 371148 117360
rect 370372 117320 371148 117348
rect 370372 117308 370378 117320
rect 371142 117308 371148 117320
rect 371200 117308 371206 117360
rect 372154 117308 372160 117360
rect 372212 117348 372218 117360
rect 372430 117348 372436 117360
rect 372212 117320 372436 117348
rect 372212 117308 372218 117320
rect 372430 117308 372436 117320
rect 372488 117308 372494 117360
rect 374546 117308 374552 117360
rect 374604 117348 374610 117360
rect 375190 117348 375196 117360
rect 374604 117320 375196 117348
rect 374604 117308 374610 117320
rect 375190 117308 375196 117320
rect 375248 117308 375254 117360
rect 375834 117308 375840 117360
rect 375892 117348 375898 117360
rect 376662 117348 376668 117360
rect 375892 117320 376668 117348
rect 375892 117308 375898 117320
rect 376662 117308 376668 117320
rect 376720 117308 376726 117360
rect 377674 117308 377680 117360
rect 377732 117348 377738 117360
rect 378042 117348 378048 117360
rect 377732 117320 378048 117348
rect 377732 117308 377738 117320
rect 378042 117308 378048 117320
rect 378100 117308 378106 117360
rect 378870 117308 378876 117360
rect 378928 117348 378934 117360
rect 379422 117348 379428 117360
rect 378928 117320 379428 117348
rect 378928 117308 378934 117320
rect 379422 117308 379428 117320
rect 379480 117308 379486 117360
rect 380066 117308 380072 117360
rect 380124 117348 380130 117360
rect 380802 117348 380808 117360
rect 380124 117320 380808 117348
rect 380124 117308 380130 117320
rect 380802 117308 380808 117320
rect 380860 117308 380866 117360
rect 381354 117308 381360 117360
rect 381412 117348 381418 117360
rect 382182 117348 382188 117360
rect 381412 117320 382188 117348
rect 381412 117308 381418 117320
rect 382182 117308 382188 117320
rect 382240 117308 382246 117360
rect 382550 117308 382556 117360
rect 382608 117348 382614 117360
rect 383562 117348 383568 117360
rect 382608 117320 383568 117348
rect 382608 117308 382614 117320
rect 383562 117308 383568 117320
rect 383620 117308 383626 117360
rect 385586 117308 385592 117360
rect 385644 117348 385650 117360
rect 386322 117348 386328 117360
rect 385644 117320 386328 117348
rect 385644 117308 385650 117320
rect 386322 117308 386328 117320
rect 386380 117308 386386 117360
rect 386782 117308 386788 117360
rect 386840 117348 386846 117360
rect 387610 117348 387616 117360
rect 386840 117320 387616 117348
rect 386840 117308 386846 117320
rect 387610 117308 387616 117320
rect 387668 117308 387674 117360
rect 388070 117308 388076 117360
rect 388128 117348 388134 117360
rect 389082 117348 389088 117360
rect 388128 117320 389088 117348
rect 388128 117308 388134 117320
rect 389082 117308 389088 117320
rect 389140 117308 389146 117360
rect 391106 117308 391112 117360
rect 391164 117348 391170 117360
rect 391750 117348 391756 117360
rect 391164 117320 391756 117348
rect 391164 117308 391170 117320
rect 391750 117308 391756 117320
rect 391808 117308 391814 117360
rect 392302 117308 392308 117360
rect 392360 117348 392366 117360
rect 393130 117348 393136 117360
rect 392360 117320 393136 117348
rect 392360 117308 392366 117320
rect 393130 117308 393136 117320
rect 393188 117308 393194 117360
rect 395430 117308 395436 117360
rect 395488 117348 395494 117360
rect 395982 117348 395988 117360
rect 395488 117320 395988 117348
rect 395488 117308 395494 117320
rect 395982 117308 395988 117320
rect 396040 117308 396046 117360
rect 396626 117308 396632 117360
rect 396684 117348 396690 117360
rect 397362 117348 397368 117360
rect 396684 117320 397368 117348
rect 396684 117308 396690 117320
rect 397362 117308 397368 117320
rect 397420 117308 397426 117360
rect 397822 117308 397828 117360
rect 397880 117348 397886 117360
rect 398742 117348 398748 117360
rect 397880 117320 398748 117348
rect 397880 117308 397886 117320
rect 398742 117308 398748 117320
rect 398800 117308 398806 117360
rect 399110 117308 399116 117360
rect 399168 117348 399174 117360
rect 400122 117348 400128 117360
rect 399168 117320 400128 117348
rect 399168 117308 399174 117320
rect 400122 117308 400128 117320
rect 400180 117308 400186 117360
rect 402146 117308 402152 117360
rect 402204 117348 402210 117360
rect 402790 117348 402796 117360
rect 402204 117320 402796 117348
rect 402204 117308 402210 117320
rect 402790 117308 402796 117320
rect 402848 117308 402854 117360
rect 403342 117308 403348 117360
rect 403400 117348 403406 117360
rect 404262 117348 404268 117360
rect 403400 117320 404268 117348
rect 403400 117308 403406 117320
rect 404262 117308 404268 117320
rect 404320 117308 404326 117360
rect 406378 117308 406384 117360
rect 406436 117348 406442 117360
rect 407022 117348 407028 117360
rect 406436 117320 407028 117348
rect 406436 117308 406442 117320
rect 407022 117308 407028 117320
rect 407080 117308 407086 117360
rect 407666 117308 407672 117360
rect 407724 117348 407730 117360
rect 408402 117348 408408 117360
rect 407724 117320 408408 117348
rect 407724 117308 407730 117320
rect 408402 117308 408408 117320
rect 408460 117308 408466 117360
rect 413186 117308 413192 117360
rect 413244 117348 413250 117360
rect 413922 117348 413928 117360
rect 413244 117320 413928 117348
rect 413244 117308 413250 117320
rect 413922 117308 413928 117320
rect 413980 117308 413986 117360
rect 414382 117308 414388 117360
rect 414440 117348 414446 117360
rect 415302 117348 415308 117360
rect 414440 117320 415308 117348
rect 414440 117308 414446 117320
rect 415302 117308 415308 117320
rect 415360 117308 415366 117360
rect 416148 117348 416176 117524
rect 417418 117512 417424 117564
rect 417476 117552 417482 117564
rect 420733 117555 420791 117561
rect 420733 117552 420745 117555
rect 417476 117524 420745 117552
rect 417476 117512 417482 117524
rect 420733 117521 420745 117524
rect 420779 117521 420791 117555
rect 420733 117515 420791 117521
rect 420822 117512 420828 117564
rect 420880 117552 420886 117564
rect 426529 117555 426587 117561
rect 426529 117552 426541 117555
rect 420880 117524 426541 117552
rect 420880 117512 420886 117524
rect 426529 117521 426541 117524
rect 426575 117521 426587 117555
rect 426529 117515 426587 117521
rect 427262 117512 427268 117564
rect 427320 117552 427326 117564
rect 427722 117552 427728 117564
rect 427320 117524 427728 117552
rect 427320 117512 427326 117524
rect 427722 117512 427728 117524
rect 427780 117512 427786 117564
rect 427817 117555 427875 117561
rect 427817 117521 427829 117555
rect 427863 117552 427875 117555
rect 429838 117552 429844 117564
rect 427863 117524 429844 117552
rect 427863 117521 427875 117524
rect 427817 117515 427875 117521
rect 429838 117512 429844 117524
rect 429896 117512 429902 117564
rect 430298 117512 430304 117564
rect 430356 117552 430362 117564
rect 431218 117552 431224 117564
rect 430356 117524 431224 117552
rect 430356 117512 430362 117524
rect 431218 117512 431224 117524
rect 431276 117512 431282 117564
rect 431770 117512 431776 117564
rect 431828 117552 431834 117564
rect 432601 117555 432659 117561
rect 431828 117524 432000 117552
rect 431828 117512 431834 117524
rect 422680 117456 425376 117484
rect 416222 117376 416228 117428
rect 416280 117416 416286 117428
rect 416682 117416 416688 117428
rect 416280 117388 416688 117416
rect 416280 117376 416286 117388
rect 416682 117376 416688 117388
rect 416740 117376 416746 117428
rect 418614 117376 418620 117428
rect 418672 117416 418678 117428
rect 419442 117416 419448 117428
rect 418672 117388 419448 117416
rect 418672 117376 418678 117388
rect 419442 117376 419448 117388
rect 419500 117376 419506 117428
rect 419902 117376 419908 117428
rect 419960 117416 419966 117428
rect 420822 117416 420828 117428
rect 419960 117388 420828 117416
rect 419960 117376 419966 117388
rect 420822 117376 420828 117388
rect 420880 117376 420886 117428
rect 421742 117376 421748 117428
rect 421800 117416 421806 117428
rect 422202 117416 422208 117428
rect 421800 117388 422208 117416
rect 421800 117376 421806 117388
rect 422202 117376 422208 117388
rect 422260 117376 422266 117428
rect 422680 117348 422708 117456
rect 422757 117419 422815 117425
rect 422757 117385 422769 117419
rect 422803 117416 422815 117419
rect 422803 117388 424088 117416
rect 422803 117385 422815 117388
rect 422757 117379 422815 117385
rect 416148 117320 422708 117348
rect 246025 117283 246083 117289
rect 246025 117280 246037 117283
rect 244384 117252 246037 117280
rect 246025 117249 246037 117252
rect 246071 117249 246083 117283
rect 424060 117280 424088 117388
rect 424134 117376 424140 117428
rect 424192 117416 424198 117428
rect 424962 117416 424968 117428
rect 424192 117388 424968 117416
rect 424192 117376 424198 117388
rect 424962 117376 424968 117388
rect 425020 117376 425026 117428
rect 425348 117348 425376 117456
rect 429654 117444 429660 117496
rect 429712 117484 429718 117496
rect 430482 117484 430488 117496
rect 429712 117456 430488 117484
rect 429712 117444 429718 117456
rect 430482 117444 430488 117456
rect 430540 117444 430546 117496
rect 430942 117444 430948 117496
rect 431000 117484 431006 117496
rect 431862 117484 431868 117496
rect 431000 117456 431868 117484
rect 431000 117444 431006 117456
rect 431862 117444 431868 117456
rect 431920 117444 431926 117496
rect 431972 117484 432000 117524
rect 432601 117521 432613 117555
rect 432647 117552 432659 117555
rect 495345 117555 495403 117561
rect 495345 117552 495357 117555
rect 432647 117524 495357 117552
rect 432647 117521 432659 117524
rect 432601 117515 432659 117521
rect 495345 117521 495357 117524
rect 495391 117521 495403 117555
rect 495345 117515 495403 117521
rect 495437 117555 495495 117561
rect 495437 117521 495449 117555
rect 495483 117552 495495 117555
rect 502978 117552 502984 117564
rect 495483 117524 502984 117552
rect 495483 117521 495495 117524
rect 495437 117515 495495 117521
rect 502978 117512 502984 117524
rect 503036 117512 503042 117564
rect 432693 117487 432751 117493
rect 432693 117484 432705 117487
rect 431972 117456 432705 117484
rect 432693 117453 432705 117456
rect 432739 117453 432751 117487
rect 432693 117447 432751 117453
rect 432782 117444 432788 117496
rect 432840 117484 432846 117496
rect 433242 117484 433248 117496
rect 432840 117456 433248 117484
rect 432840 117444 432846 117456
rect 433242 117444 433248 117456
rect 433300 117444 433306 117496
rect 434625 117487 434683 117493
rect 434625 117453 434637 117487
rect 434671 117484 434683 117487
rect 444377 117487 444435 117493
rect 444377 117484 444389 117487
rect 434671 117456 444389 117484
rect 434671 117453 434683 117456
rect 434625 117447 434683 117453
rect 444377 117453 444389 117456
rect 444423 117453 444435 117487
rect 444377 117447 444435 117453
rect 456705 117487 456763 117493
rect 456705 117453 456717 117487
rect 456751 117484 456763 117487
rect 463697 117487 463755 117493
rect 463697 117484 463709 117487
rect 456751 117456 463709 117484
rect 456751 117453 456763 117456
rect 456705 117447 456763 117453
rect 463697 117453 463709 117456
rect 463743 117453 463755 117487
rect 463697 117447 463755 117453
rect 476025 117487 476083 117493
rect 476025 117453 476037 117487
rect 476071 117484 476083 117487
rect 492585 117487 492643 117493
rect 492585 117484 492597 117487
rect 476071 117456 492597 117484
rect 476071 117453 476083 117456
rect 476025 117447 476083 117453
rect 492585 117453 492597 117456
rect 492631 117453 492643 117487
rect 492585 117447 492643 117453
rect 425422 117376 425428 117428
rect 425480 117416 425486 117428
rect 426342 117416 426348 117428
rect 425480 117388 426348 117416
rect 425480 117376 425486 117388
rect 426342 117376 426348 117388
rect 426400 117376 426406 117428
rect 426437 117419 426495 117425
rect 426437 117385 426449 117419
rect 426483 117416 426495 117419
rect 493318 117416 493324 117428
rect 426483 117388 493324 117416
rect 426483 117385 426495 117388
rect 426437 117379 426495 117385
rect 493318 117376 493324 117388
rect 493376 117376 493382 117428
rect 489178 117348 489184 117360
rect 425348 117320 489184 117348
rect 489178 117308 489184 117320
rect 489236 117308 489242 117360
rect 425057 117283 425115 117289
rect 425057 117280 425069 117283
rect 424060 117252 425069 117280
rect 246025 117243 246083 117249
rect 425057 117249 425069 117252
rect 425103 117249 425115 117283
rect 425057 117243 425115 117249
rect 235123 117184 239720 117212
rect 235123 117181 235135 117184
rect 235077 117175 235135 117181
rect 186133 117147 186191 117153
rect 180720 117116 180794 117144
rect 167656 117076 167684 117116
rect 164068 117048 167684 117076
rect 143537 117011 143595 117017
rect 143537 116977 143549 117011
rect 143583 117008 143595 117011
rect 151817 117011 151875 117017
rect 151817 117008 151829 117011
rect 143583 116980 151829 117008
rect 143583 116977 143595 116980
rect 143537 116971 143595 116977
rect 151817 116977 151829 116980
rect 151863 116977 151875 117011
rect 180766 117008 180794 117116
rect 186133 117113 186145 117147
rect 186179 117144 186191 117147
rect 192018 117144 192024 117156
rect 186179 117116 192024 117144
rect 186179 117113 186191 117116
rect 186133 117107 186191 117113
rect 192018 117104 192024 117116
rect 192076 117104 192082 117156
rect 425057 117147 425115 117153
rect 425057 117113 425069 117147
rect 425103 117144 425115 117147
rect 434625 117147 434683 117153
rect 434625 117144 434637 117147
rect 425103 117116 434637 117144
rect 425103 117113 425115 117116
rect 425057 117107 425115 117113
rect 434625 117113 434637 117116
rect 434671 117113 434683 117147
rect 434625 117107 434683 117113
rect 180766 116980 190408 117008
rect 151817 116971 151875 116977
rect 190380 116804 190408 116980
rect 492677 116943 492735 116949
rect 492677 116909 492689 116943
rect 492723 116940 492735 116943
rect 496078 116940 496084 116952
rect 492723 116912 496084 116940
rect 492723 116909 492735 116912
rect 492677 116903 492735 116909
rect 496078 116900 496084 116912
rect 496136 116900 496142 116952
rect 190546 116804 190552 116816
rect 190380 116776 190552 116804
rect 190546 116764 190552 116776
rect 190604 116764 190610 116816
rect 202966 116628 202972 116680
rect 203024 116668 203030 116680
rect 203150 116668 203156 116680
rect 203024 116640 203156 116668
rect 203024 116628 203030 116640
rect 203150 116628 203156 116640
rect 203208 116628 203214 116680
rect 197354 116560 197360 116612
rect 197412 116600 197418 116612
rect 198182 116600 198188 116612
rect 197412 116572 198188 116600
rect 197412 116560 197418 116572
rect 198182 116560 198188 116572
rect 198240 116560 198246 116612
rect 198734 116560 198740 116612
rect 198792 116600 198798 116612
rect 199470 116600 199476 116612
rect 198792 116572 199476 116600
rect 198792 116560 198798 116572
rect 199470 116560 199476 116572
rect 199528 116560 199534 116612
rect 201494 116560 201500 116612
rect 201552 116600 201558 116612
rect 201862 116600 201868 116612
rect 201552 116572 201868 116600
rect 201552 116560 201558 116572
rect 201862 116560 201868 116572
rect 201920 116560 201926 116612
rect 202874 116560 202880 116612
rect 202932 116600 202938 116612
rect 203702 116600 203708 116612
rect 202932 116572 203708 116600
rect 202932 116560 202938 116572
rect 203702 116560 203708 116572
rect 203760 116560 203766 116612
rect 204254 116560 204260 116612
rect 204312 116600 204318 116612
rect 204898 116600 204904 116612
rect 204312 116572 204904 116600
rect 204312 116560 204318 116572
rect 204898 116560 204904 116572
rect 204956 116560 204962 116612
rect 403710 116016 403716 116068
rect 403768 116056 403774 116068
rect 403986 116056 403992 116068
rect 403768 116028 403992 116056
rect 403768 116016 403774 116028
rect 403986 116016 403992 116028
rect 404044 116016 404050 116068
rect 221458 115948 221464 116000
rect 221516 115988 221522 116000
rect 221642 115988 221648 116000
rect 221516 115960 221648 115988
rect 221516 115948 221522 115960
rect 221642 115948 221648 115960
rect 221700 115948 221706 116000
rect 272242 115948 272248 116000
rect 272300 115988 272306 116000
rect 272426 115988 272432 116000
rect 272300 115960 272432 115988
rect 272300 115948 272306 115960
rect 272426 115948 272432 115960
rect 272484 115948 272490 116000
rect 301406 115948 301412 116000
rect 301464 115988 301470 116000
rect 301590 115988 301596 116000
rect 301464 115960 301596 115988
rect 301464 115948 301470 115960
rect 301590 115948 301596 115960
rect 301648 115948 301654 116000
rect 322382 115948 322388 116000
rect 322440 115988 322446 116000
rect 322566 115988 322572 116000
rect 322440 115960 322572 115988
rect 322440 115948 322446 115960
rect 322566 115948 322572 115960
rect 322624 115948 322630 116000
rect 382918 115948 382924 116000
rect 382976 115988 382982 116000
rect 383102 115988 383108 116000
rect 382976 115960 383108 115988
rect 382976 115948 382982 115960
rect 383102 115948 383108 115960
rect 383160 115948 383166 116000
rect 420270 115948 420276 116000
rect 420328 115988 420334 116000
rect 420454 115988 420460 116000
rect 420328 115960 420460 115988
rect 420328 115948 420334 115960
rect 420454 115948 420460 115960
rect 420512 115948 420518 116000
rect 425882 115948 425888 116000
rect 425940 115988 425946 116000
rect 425974 115988 425980 116000
rect 425940 115960 425980 115988
rect 425940 115948 425946 115960
rect 425974 115948 425980 115960
rect 426032 115948 426038 116000
rect 431310 115948 431316 116000
rect 431368 115988 431374 116000
rect 431494 115988 431500 116000
rect 431368 115960 431500 115988
rect 431368 115948 431374 115960
rect 431494 115948 431500 115960
rect 431552 115948 431558 116000
rect 73890 115920 73896 115932
rect 73851 115892 73896 115920
rect 73890 115880 73896 115892
rect 73948 115880 73954 115932
rect 133046 115920 133052 115932
rect 133007 115892 133052 115920
rect 133046 115880 133052 115892
rect 133104 115880 133110 115932
rect 183738 115880 183744 115932
rect 183796 115920 183802 115932
rect 183922 115920 183928 115932
rect 183796 115892 183928 115920
rect 183796 115880 183802 115892
rect 183922 115880 183928 115892
rect 183980 115880 183986 115932
rect 184750 115880 184756 115932
rect 184808 115920 184814 115932
rect 185026 115920 185032 115932
rect 184808 115892 185032 115920
rect 184808 115880 184814 115892
rect 185026 115880 185032 115892
rect 185084 115880 185090 115932
rect 233418 115880 233424 115932
rect 233476 115920 233482 115932
rect 233602 115920 233608 115932
rect 233476 115892 233608 115920
rect 233476 115880 233482 115892
rect 233602 115880 233608 115892
rect 233660 115880 233666 115932
rect 243630 115880 243636 115932
rect 243688 115920 243694 115932
rect 243906 115920 243912 115932
rect 243688 115892 243912 115920
rect 243688 115880 243694 115892
rect 243906 115880 243912 115892
rect 243964 115880 243970 115932
rect 248322 115920 248328 115932
rect 248283 115892 248328 115920
rect 248322 115880 248328 115892
rect 248380 115880 248386 115932
rect 341058 115880 341064 115932
rect 341116 115920 341122 115932
rect 341334 115920 341340 115932
rect 341116 115892 341340 115920
rect 341116 115880 341122 115892
rect 341334 115880 341340 115892
rect 341392 115880 341398 115932
rect 388714 115880 388720 115932
rect 388772 115920 388778 115932
rect 388898 115920 388904 115932
rect 388772 115892 388904 115920
rect 388772 115880 388778 115892
rect 388898 115880 388904 115892
rect 388956 115880 388962 115932
rect 403897 115923 403955 115929
rect 403897 115889 403909 115923
rect 403943 115920 403955 115923
rect 403986 115920 403992 115932
rect 403943 115892 403992 115920
rect 403943 115889 403955 115892
rect 403897 115883 403955 115889
rect 403986 115880 403992 115892
rect 404044 115880 404050 115932
rect 414842 115880 414848 115932
rect 414900 115920 414906 115932
rect 414934 115920 414940 115932
rect 414900 115892 414940 115920
rect 414900 115880 414906 115892
rect 414934 115880 414940 115892
rect 414992 115880 414998 115932
rect 420454 115852 420460 115864
rect 420415 115824 420460 115852
rect 420454 115812 420460 115824
rect 420512 115812 420518 115864
rect 131117 114563 131175 114569
rect 131117 114529 131129 114563
rect 131163 114560 131175 114563
rect 131206 114560 131212 114572
rect 131163 114532 131212 114560
rect 131163 114529 131175 114532
rect 131117 114523 131175 114529
rect 131206 114520 131212 114532
rect 131264 114520 131270 114572
rect 150894 114520 150900 114572
rect 150952 114560 150958 114572
rect 151170 114560 151176 114572
rect 150952 114532 151176 114560
rect 150952 114520 150958 114532
rect 151170 114520 151176 114532
rect 151228 114520 151234 114572
rect 157426 114520 157432 114572
rect 157484 114560 157490 114572
rect 157794 114560 157800 114572
rect 157484 114532 157800 114560
rect 157484 114520 157490 114532
rect 157794 114520 157800 114532
rect 157852 114520 157858 114572
rect 325694 114560 325700 114572
rect 325655 114532 325700 114560
rect 325694 114520 325700 114532
rect 325752 114520 325758 114572
rect 243725 114495 243783 114501
rect 243725 114461 243737 114495
rect 243771 114492 243783 114495
rect 243906 114492 243912 114504
rect 243771 114464 243912 114492
rect 243771 114461 243783 114464
rect 243725 114455 243783 114461
rect 243906 114452 243912 114464
rect 243964 114452 243970 114504
rect 272242 114492 272248 114504
rect 272203 114464 272248 114492
rect 272242 114452 272248 114464
rect 272300 114452 272306 114504
rect 213914 113976 213920 114028
rect 213972 114016 213978 114028
rect 214190 114016 214196 114028
rect 213972 113988 214196 114016
rect 213972 113976 213978 113988
rect 214190 113976 214196 113988
rect 214248 113976 214254 114028
rect 133874 113840 133880 113892
rect 133932 113880 133938 113892
rect 134518 113880 134524 113892
rect 133932 113852 134524 113880
rect 133932 113840 133938 113852
rect 134518 113840 134524 113852
rect 134576 113840 134582 113892
rect 135254 113840 135260 113892
rect 135312 113880 135318 113892
rect 135714 113880 135720 113892
rect 135312 113852 135720 113880
rect 135312 113840 135318 113852
rect 135714 113840 135720 113852
rect 135772 113840 135778 113892
rect 136726 113840 136732 113892
rect 136784 113880 136790 113892
rect 137554 113880 137560 113892
rect 136784 113852 137560 113880
rect 136784 113840 136790 113852
rect 137554 113840 137560 113852
rect 137612 113840 137618 113892
rect 139486 113840 139492 113892
rect 139544 113880 139550 113892
rect 140038 113880 140044 113892
rect 139544 113852 140044 113880
rect 139544 113840 139550 113852
rect 140038 113840 140044 113852
rect 140096 113840 140102 113892
rect 140774 113840 140780 113892
rect 140832 113880 140838 113892
rect 141234 113880 141240 113892
rect 140832 113852 141240 113880
rect 140832 113840 140838 113852
rect 141234 113840 141240 113852
rect 141292 113840 141298 113892
rect 146294 113840 146300 113892
rect 146352 113880 146358 113892
rect 146754 113880 146760 113892
rect 146352 113852 146760 113880
rect 146352 113840 146358 113852
rect 146754 113840 146760 113852
rect 146812 113840 146818 113892
rect 153194 113840 153200 113892
rect 153252 113880 153258 113892
rect 154114 113880 154120 113892
rect 153252 113852 154120 113880
rect 153252 113840 153258 113852
rect 154114 113840 154120 113852
rect 154172 113840 154178 113892
rect 161474 113840 161480 113892
rect 161532 113880 161538 113892
rect 162118 113880 162124 113892
rect 161532 113852 162124 113880
rect 161532 113840 161538 113852
rect 162118 113840 162124 113852
rect 162176 113840 162182 113892
rect 166994 113840 167000 113892
rect 167052 113880 167058 113892
rect 167638 113880 167644 113892
rect 167052 113852 167644 113880
rect 167052 113840 167058 113852
rect 167638 113840 167644 113852
rect 167696 113840 167702 113892
rect 169846 113840 169852 113892
rect 169904 113880 169910 113892
rect 170674 113880 170680 113892
rect 169904 113852 170680 113880
rect 169904 113840 169910 113852
rect 170674 113840 170680 113852
rect 170732 113840 170738 113892
rect 189166 113840 189172 113892
rect 189224 113880 189230 113892
rect 189626 113880 189632 113892
rect 189224 113852 189632 113880
rect 189224 113840 189230 113852
rect 189626 113840 189632 113852
rect 189684 113840 189690 113892
rect 191834 113840 191840 113892
rect 191892 113880 191898 113892
rect 192662 113880 192668 113892
rect 191892 113852 192668 113880
rect 191892 113840 191898 113852
rect 192662 113840 192668 113852
rect 192720 113840 192726 113892
rect 213914 113840 213920 113892
rect 213972 113880 213978 113892
rect 214098 113880 214104 113892
rect 213972 113852 214104 113880
rect 213972 113840 213978 113852
rect 214098 113840 214104 113852
rect 214156 113840 214162 113892
rect 215294 113840 215300 113892
rect 215352 113880 215358 113892
rect 215938 113880 215944 113892
rect 215352 113852 215944 113880
rect 215352 113840 215358 113852
rect 215938 113840 215944 113852
rect 215996 113840 216002 113892
rect 218054 113840 218060 113892
rect 218112 113880 218118 113892
rect 218422 113880 218428 113892
rect 218112 113852 218428 113880
rect 218112 113840 218118 113852
rect 218422 113840 218428 113852
rect 218480 113840 218486 113892
rect 219526 113840 219532 113892
rect 219584 113880 219590 113892
rect 219710 113880 219716 113892
rect 219584 113852 219716 113880
rect 219584 113840 219590 113852
rect 219710 113840 219716 113852
rect 219768 113840 219774 113892
rect 222194 113840 222200 113892
rect 222252 113880 222258 113892
rect 222654 113880 222660 113892
rect 222252 113852 222660 113880
rect 222252 113840 222258 113852
rect 222654 113840 222660 113852
rect 222712 113840 222718 113892
rect 231854 113840 231860 113892
rect 231912 113880 231918 113892
rect 232498 113880 232504 113892
rect 231912 113852 232504 113880
rect 231912 113840 231918 113852
rect 232498 113840 232504 113852
rect 232556 113840 232562 113892
rect 248506 113840 248512 113892
rect 248564 113880 248570 113892
rect 249058 113880 249064 113892
rect 248564 113852 249064 113880
rect 248564 113840 248570 113852
rect 249058 113840 249064 113852
rect 249116 113840 249122 113892
rect 173894 113160 173900 113212
rect 173952 113200 173958 113212
rect 174354 113200 174360 113212
rect 173952 113172 174360 113200
rect 173952 113160 173958 113172
rect 174354 113160 174360 113172
rect 174412 113160 174418 113212
rect 175550 113160 175556 113212
rect 175608 113200 175614 113212
rect 176194 113200 176200 113212
rect 175608 113172 176200 113200
rect 175608 113160 175614 113172
rect 176194 113160 176200 113172
rect 176252 113160 176258 113212
rect 178126 113160 178132 113212
rect 178184 113200 178190 113212
rect 178586 113200 178592 113212
rect 178184 113172 178592 113200
rect 178184 113160 178190 113172
rect 178586 113160 178592 113172
rect 178644 113160 178650 113212
rect 179414 113160 179420 113212
rect 179472 113200 179478 113212
rect 179874 113200 179880 113212
rect 179472 113172 179880 113200
rect 179472 113160 179478 113172
rect 179874 113160 179880 113172
rect 179932 113160 179938 113212
rect 180978 113132 180984 113144
rect 180939 113104 180984 113132
rect 180978 113092 180984 113104
rect 181036 113092 181042 113144
rect 200206 113092 200212 113144
rect 200264 113132 200270 113144
rect 200390 113132 200396 113144
rect 200264 113104 200396 113132
rect 200264 113092 200270 113104
rect 200390 113092 200396 113104
rect 200448 113092 200454 113144
rect 436922 111732 436928 111784
rect 436980 111772 436986 111784
rect 579798 111772 579804 111784
rect 436980 111744 579804 111772
rect 436980 111732 436986 111744
rect 579798 111732 579804 111744
rect 579856 111732 579862 111784
rect 172514 111596 172520 111648
rect 172572 111636 172578 111648
rect 173066 111636 173072 111648
rect 172572 111608 173072 111636
rect 172572 111596 172578 111608
rect 173066 111596 173072 111608
rect 173124 111596 173130 111648
rect 212626 110412 212632 110424
rect 212587 110384 212632 110412
rect 212626 110372 212632 110384
rect 212684 110372 212690 110424
rect 194689 109735 194747 109741
rect 194689 109701 194701 109735
rect 194735 109732 194747 109735
rect 194778 109732 194784 109744
rect 194735 109704 194784 109732
rect 194735 109701 194747 109704
rect 194689 109695 194747 109701
rect 194778 109692 194784 109704
rect 194836 109692 194842 109744
rect 205910 109080 205916 109132
rect 205968 109080 205974 109132
rect 207106 109080 207112 109132
rect 207164 109080 207170 109132
rect 205928 108996 205956 109080
rect 207124 108996 207152 109080
rect 214098 109012 214104 109064
rect 214156 109052 214162 109064
rect 214558 109052 214564 109064
rect 214156 109024 214564 109052
rect 214156 109012 214162 109024
rect 214558 109012 214564 109024
rect 214616 109012 214622 109064
rect 234706 109012 234712 109064
rect 234764 109052 234770 109064
rect 235442 109052 235448 109064
rect 234764 109024 235448 109052
rect 234764 109012 234770 109024
rect 235442 109012 235448 109024
rect 235500 109012 235506 109064
rect 387518 109012 387524 109064
rect 387576 109052 387582 109064
rect 387702 109052 387708 109064
rect 387576 109024 387708 109052
rect 387576 109012 387582 109024
rect 387702 109012 387708 109024
rect 387760 109012 387766 109064
rect 393038 109012 393044 109064
rect 393096 109052 393102 109064
rect 393222 109052 393228 109064
rect 393096 109024 393228 109052
rect 393096 109012 393102 109024
rect 393222 109012 393228 109024
rect 393280 109012 393286 109064
rect 73890 108984 73896 108996
rect 73851 108956 73896 108984
rect 73890 108944 73896 108956
rect 73948 108944 73954 108996
rect 205910 108944 205916 108996
rect 205968 108944 205974 108996
rect 207106 108944 207112 108996
rect 207164 108944 207170 108996
rect 420457 108987 420515 108993
rect 420457 108953 420469 108987
rect 420503 108984 420515 108987
rect 420638 108984 420644 108996
rect 420503 108956 420644 108984
rect 420503 108953 420515 108956
rect 420457 108947 420515 108953
rect 420638 108944 420644 108956
rect 420696 108944 420702 108996
rect 238846 106292 238852 106344
rect 238904 106332 238910 106344
rect 238938 106332 238944 106344
rect 238904 106304 238944 106332
rect 238904 106292 238910 106304
rect 238938 106292 238944 106304
rect 238996 106292 239002 106344
rect 248322 106332 248328 106344
rect 248283 106304 248328 106332
rect 248322 106292 248328 106304
rect 248380 106292 248386 106344
rect 403894 106332 403900 106344
rect 403855 106304 403900 106332
rect 403894 106292 403900 106304
rect 403952 106292 403958 106344
rect 131298 106264 131304 106276
rect 131259 106236 131304 106264
rect 131298 106224 131304 106236
rect 131356 106224 131362 106276
rect 301958 106264 301964 106276
rect 301919 106236 301964 106264
rect 301958 106224 301964 106236
rect 302016 106224 302022 106276
rect 322658 106264 322664 106276
rect 322619 106236 322664 106264
rect 322658 106224 322664 106236
rect 322716 106224 322722 106276
rect 388714 106224 388720 106276
rect 388772 106264 388778 106276
rect 388806 106264 388812 106276
rect 388772 106236 388812 106264
rect 388772 106224 388778 106236
rect 388806 106224 388812 106236
rect 388864 106224 388870 106276
rect 394418 106264 394424 106276
rect 394379 106236 394424 106264
rect 394418 106224 394424 106236
rect 394476 106224 394482 106276
rect 431678 106264 431684 106276
rect 431639 106236 431684 106264
rect 431678 106224 431684 106236
rect 431736 106224 431742 106276
rect 183646 106156 183652 106208
rect 183704 106196 183710 106208
rect 183922 106196 183928 106208
rect 183704 106168 183928 106196
rect 183704 106156 183710 106168
rect 183922 106156 183928 106168
rect 183980 106156 183986 106208
rect 148226 104864 148232 104916
rect 148284 104904 148290 104916
rect 148502 104904 148508 104916
rect 148284 104876 148508 104904
rect 148284 104864 148290 104876
rect 148502 104864 148508 104876
rect 148560 104864 148566 104916
rect 194686 104904 194692 104916
rect 194647 104876 194692 104904
rect 194686 104864 194692 104876
rect 194744 104864 194750 104916
rect 243722 104904 243728 104916
rect 243683 104876 243728 104904
rect 243722 104864 243728 104876
rect 243780 104864 243786 104916
rect 274910 104864 274916 104916
rect 274968 104904 274974 104916
rect 275370 104904 275376 104916
rect 274968 104876 275376 104904
rect 274968 104864 274974 104876
rect 275370 104864 275376 104876
rect 275428 104864 275434 104916
rect 133141 104839 133199 104845
rect 133141 104805 133153 104839
rect 133187 104836 133199 104839
rect 133414 104836 133420 104848
rect 133187 104808 133420 104836
rect 133187 104805 133199 104808
rect 133141 104799 133199 104805
rect 133414 104796 133420 104808
rect 133472 104796 133478 104848
rect 233418 104836 233424 104848
rect 233379 104808 233424 104836
rect 233418 104796 233424 104808
rect 233476 104796 233482 104848
rect 248233 104839 248291 104845
rect 248233 104805 248245 104839
rect 248279 104836 248291 104839
rect 248322 104836 248328 104848
rect 248279 104808 248328 104836
rect 248279 104805 248291 104808
rect 248233 104799 248291 104805
rect 248322 104796 248328 104808
rect 248380 104796 248386 104848
rect 325694 104836 325700 104848
rect 325655 104808 325700 104836
rect 325694 104796 325700 104808
rect 325752 104796 325758 104848
rect 415026 104836 415032 104848
rect 414987 104808 415032 104836
rect 415026 104796 415032 104808
rect 415084 104796 415090 104848
rect 420638 104836 420644 104848
rect 420599 104808 420644 104836
rect 420638 104796 420644 104808
rect 420696 104796 420702 104848
rect 180981 104771 181039 104777
rect 180981 104737 180993 104771
rect 181027 104768 181039 104771
rect 181070 104768 181076 104780
rect 181027 104740 181076 104768
rect 181027 104737 181039 104740
rect 180981 104731 181039 104737
rect 181070 104728 181076 104740
rect 181128 104728 181134 104780
rect 157242 103504 157248 103556
rect 157300 103544 157306 103556
rect 157426 103544 157432 103556
rect 157300 103516 157432 103544
rect 157300 103504 157306 103516
rect 157426 103504 157432 103516
rect 157484 103504 157490 103556
rect 272058 103504 272064 103556
rect 272116 103544 272122 103556
rect 272245 103547 272303 103553
rect 272245 103544 272257 103547
rect 272116 103516 272257 103544
rect 272116 103504 272122 103516
rect 272245 103513 272257 103516
rect 272291 103513 272303 103547
rect 272245 103507 272303 103513
rect 173894 103436 173900 103488
rect 173952 103436 173958 103488
rect 178126 103436 178132 103488
rect 178184 103476 178190 103488
rect 178310 103476 178316 103488
rect 178184 103448 178316 103476
rect 178184 103436 178190 103448
rect 178310 103436 178316 103448
rect 178368 103436 178374 103488
rect 179414 103436 179420 103488
rect 179472 103436 179478 103488
rect 279786 103436 279792 103488
rect 279844 103476 279850 103488
rect 279970 103476 279976 103488
rect 279844 103448 279976 103476
rect 279844 103436 279850 103448
rect 279970 103436 279976 103448
rect 280028 103436 280034 103488
rect 173912 103408 173940 103436
rect 173986 103408 173992 103420
rect 173912 103380 173992 103408
rect 173986 103368 173992 103380
rect 174044 103368 174050 103420
rect 179432 103408 179460 103436
rect 179506 103408 179512 103420
rect 179432 103380 179512 103408
rect 179506 103368 179512 103380
rect 179564 103368 179570 103420
rect 212629 100759 212687 100765
rect 212629 100725 212641 100759
rect 212675 100756 212687 100759
rect 212718 100756 212724 100768
rect 212675 100728 212724 100756
rect 212675 100725 212687 100728
rect 212629 100719 212687 100725
rect 212718 100716 212724 100728
rect 212776 100716 212782 100768
rect 221090 100076 221096 100088
rect 221051 100048 221096 100076
rect 221090 100036 221096 100048
rect 221148 100036 221154 100088
rect 150710 99464 150716 99476
rect 150636 99436 150716 99464
rect 73798 99356 73804 99408
rect 73856 99396 73862 99408
rect 73982 99396 73988 99408
rect 73856 99368 73988 99396
rect 73856 99356 73862 99368
rect 73982 99356 73988 99368
rect 74040 99356 74046 99408
rect 150636 99340 150664 99436
rect 150710 99424 150716 99436
rect 150768 99424 150774 99476
rect 209866 99424 209872 99476
rect 209924 99424 209930 99476
rect 229186 99424 229192 99476
rect 229244 99424 229250 99476
rect 234706 99424 234712 99476
rect 234764 99424 234770 99476
rect 240226 99424 240232 99476
rect 240284 99424 240290 99476
rect 272058 99464 272064 99476
rect 271984 99436 272064 99464
rect 209884 99340 209912 99424
rect 216677 99399 216735 99405
rect 216677 99365 216689 99399
rect 216723 99396 216735 99399
rect 216766 99396 216772 99408
rect 216723 99368 216772 99396
rect 216723 99365 216735 99368
rect 216677 99359 216735 99365
rect 216766 99356 216772 99368
rect 216824 99356 216830 99408
rect 229204 99340 229232 99424
rect 234724 99340 234752 99424
rect 240244 99340 240272 99424
rect 243630 99356 243636 99408
rect 243688 99396 243694 99408
rect 243725 99399 243783 99405
rect 243725 99396 243737 99399
rect 243688 99368 243737 99396
rect 243688 99356 243694 99368
rect 243725 99365 243737 99368
rect 243771 99365 243783 99399
rect 243725 99359 243783 99365
rect 244366 99356 244372 99408
rect 244424 99396 244430 99408
rect 244550 99396 244556 99408
rect 244424 99368 244556 99396
rect 244424 99356 244430 99368
rect 244550 99356 244556 99368
rect 244608 99356 244614 99408
rect 245838 99356 245844 99408
rect 245896 99396 245902 99408
rect 246022 99396 246028 99408
rect 245896 99368 246028 99396
rect 245896 99356 245902 99368
rect 246022 99356 246028 99368
rect 246080 99356 246086 99408
rect 271984 99340 272012 99436
rect 272058 99424 272064 99436
rect 272116 99424 272122 99476
rect 383286 99464 383292 99476
rect 383212 99436 383292 99464
rect 341242 99356 341248 99408
rect 341300 99356 341306 99408
rect 131298 99328 131304 99340
rect 131259 99300 131304 99328
rect 131298 99288 131304 99300
rect 131356 99288 131362 99340
rect 150618 99288 150624 99340
rect 150676 99288 150682 99340
rect 209866 99288 209872 99340
rect 209924 99288 209930 99340
rect 229186 99288 229192 99340
rect 229244 99288 229250 99340
rect 234706 99288 234712 99340
rect 234764 99288 234770 99340
rect 240226 99288 240232 99340
rect 240284 99288 240290 99340
rect 271966 99288 271972 99340
rect 272024 99288 272030 99340
rect 301958 99328 301964 99340
rect 301919 99300 301964 99328
rect 301958 99288 301964 99300
rect 302016 99288 302022 99340
rect 322658 99328 322664 99340
rect 322619 99300 322664 99328
rect 322658 99288 322664 99300
rect 322716 99288 322722 99340
rect 341260 99328 341288 99356
rect 383212 99340 383240 99436
rect 383286 99424 383292 99436
rect 383344 99424 383350 99476
rect 403894 99356 403900 99408
rect 403952 99356 403958 99408
rect 341334 99328 341340 99340
rect 341260 99300 341340 99328
rect 341334 99288 341340 99300
rect 341392 99288 341398 99340
rect 383194 99288 383200 99340
rect 383252 99288 383258 99340
rect 394418 99328 394424 99340
rect 394379 99300 394424 99328
rect 394418 99288 394424 99300
rect 394476 99288 394482 99340
rect 403912 99328 403940 99356
rect 403986 99328 403992 99340
rect 403912 99300 403992 99328
rect 403986 99288 403992 99300
rect 404044 99288 404050 99340
rect 431678 99328 431684 99340
rect 431639 99300 431684 99328
rect 431678 99288 431684 99300
rect 431736 99288 431742 99340
rect 227714 96608 227720 96620
rect 227675 96580 227720 96608
rect 227714 96568 227720 96580
rect 227772 96568 227778 96620
rect 238846 96608 238852 96620
rect 238807 96580 238852 96608
rect 238846 96568 238852 96580
rect 238904 96568 238910 96620
rect 341058 96568 341064 96620
rect 341116 96608 341122 96620
rect 341334 96608 341340 96620
rect 341116 96580 341340 96608
rect 341116 96568 341122 96580
rect 341334 96568 341340 96580
rect 341392 96568 341398 96620
rect 383105 96611 383163 96617
rect 383105 96577 383117 96611
rect 383151 96608 383163 96611
rect 383194 96608 383200 96620
rect 383151 96580 383200 96608
rect 383151 96577 383163 96580
rect 383105 96571 383163 96577
rect 383194 96568 383200 96580
rect 383252 96568 383258 96620
rect 388625 96611 388683 96617
rect 388625 96577 388637 96611
rect 388671 96608 388683 96611
rect 388714 96608 388720 96620
rect 388671 96580 388720 96608
rect 388671 96577 388683 96580
rect 388625 96571 388683 96577
rect 388714 96568 388720 96580
rect 388772 96568 388778 96620
rect 403897 96611 403955 96617
rect 403897 96577 403909 96611
rect 403943 96608 403955 96611
rect 403986 96608 403992 96620
rect 403943 96580 403992 96608
rect 403943 96577 403955 96580
rect 403897 96571 403955 96577
rect 403986 96568 403992 96580
rect 404044 96568 404050 96620
rect 145098 95344 145104 95396
rect 145156 95344 145162 95396
rect 145116 95260 145144 95344
rect 133138 95248 133144 95260
rect 133099 95220 133144 95248
rect 133138 95208 133144 95220
rect 133196 95208 133202 95260
rect 145098 95208 145104 95260
rect 145156 95208 145162 95260
rect 147950 95208 147956 95260
rect 148008 95248 148014 95260
rect 148226 95248 148232 95260
rect 148008 95220 148232 95248
rect 148008 95208 148014 95220
rect 148226 95208 148232 95220
rect 148284 95208 148290 95260
rect 181070 95208 181076 95260
rect 181128 95208 181134 95260
rect 221093 95251 221151 95257
rect 221093 95217 221105 95251
rect 221139 95248 221151 95251
rect 221182 95248 221188 95260
rect 221139 95220 221188 95248
rect 221139 95217 221151 95220
rect 221093 95211 221151 95217
rect 221182 95208 221188 95220
rect 221240 95208 221246 95260
rect 233421 95251 233479 95257
rect 233421 95217 233433 95251
rect 233467 95248 233479 95251
rect 233510 95248 233516 95260
rect 233467 95220 233516 95248
rect 233467 95217 233479 95220
rect 233421 95211 233479 95217
rect 233510 95208 233516 95220
rect 233568 95208 233574 95260
rect 243722 95248 243728 95260
rect 243683 95220 243728 95248
rect 243722 95208 243728 95220
rect 243780 95208 243786 95260
rect 248230 95248 248236 95260
rect 248191 95220 248236 95248
rect 248230 95208 248236 95220
rect 248288 95208 248294 95260
rect 325694 95248 325700 95260
rect 325655 95220 325700 95248
rect 325694 95208 325700 95220
rect 325752 95208 325758 95260
rect 415029 95251 415087 95257
rect 415029 95217 415041 95251
rect 415075 95248 415087 95251
rect 415210 95248 415216 95260
rect 415075 95220 415216 95248
rect 415075 95217 415087 95220
rect 415029 95211 415087 95217
rect 415210 95208 415216 95220
rect 415268 95208 415274 95260
rect 420638 95248 420644 95260
rect 420599 95220 420644 95248
rect 420638 95208 420644 95220
rect 420696 95208 420702 95260
rect 181088 95112 181116 95208
rect 426161 95183 426219 95189
rect 426161 95149 426173 95183
rect 426207 95180 426219 95183
rect 426250 95180 426256 95192
rect 426207 95152 426256 95180
rect 426207 95149 426219 95152
rect 426161 95143 426219 95149
rect 426250 95140 426256 95152
rect 426308 95140 426314 95192
rect 181162 95112 181168 95124
rect 181088 95084 181168 95112
rect 181162 95072 181168 95084
rect 181220 95072 181226 95124
rect 206002 93956 206008 93968
rect 205928 93928 206008 93956
rect 162854 93848 162860 93900
rect 162912 93888 162918 93900
rect 163038 93888 163044 93900
rect 162912 93860 163044 93888
rect 162912 93848 162918 93860
rect 163038 93848 163044 93860
rect 163096 93848 163102 93900
rect 205928 93832 205956 93928
rect 206002 93916 206008 93928
rect 206060 93916 206066 93968
rect 156046 93820 156052 93832
rect 156007 93792 156052 93820
rect 156046 93780 156052 93792
rect 156104 93780 156110 93832
rect 205910 93780 205916 93832
rect 205968 93780 205974 93832
rect 279694 93820 279700 93832
rect 279655 93792 279700 93820
rect 279694 93780 279700 93792
rect 279752 93780 279758 93832
rect 2774 93304 2780 93356
rect 2832 93344 2838 93356
rect 5350 93344 5356 93356
rect 2832 93316 5356 93344
rect 2832 93304 2838 93316
rect 5350 93304 5356 93316
rect 5408 93304 5414 93356
rect 181162 92460 181168 92472
rect 181123 92432 181168 92460
rect 181162 92420 181168 92432
rect 181220 92420 181226 92472
rect 212718 91060 212724 91112
rect 212776 91100 212782 91112
rect 212902 91100 212908 91112
rect 212776 91072 212908 91100
rect 212776 91060 212782 91072
rect 212902 91060 212908 91072
rect 212960 91060 212966 91112
rect 216674 91060 216680 91112
rect 216732 91100 216738 91112
rect 216732 91072 216777 91100
rect 216732 91060 216738 91072
rect 207106 91032 207112 91044
rect 207067 91004 207112 91032
rect 207106 90992 207112 91004
rect 207164 90992 207170 91044
rect 144917 90423 144975 90429
rect 144917 90389 144929 90423
rect 144963 90420 144975 90423
rect 145098 90420 145104 90432
rect 144963 90392 145104 90420
rect 144963 90389 144975 90392
rect 144917 90383 144975 90389
rect 145098 90380 145104 90392
rect 145156 90380 145162 90432
rect 73709 89879 73767 89885
rect 73709 89845 73721 89879
rect 73755 89876 73767 89879
rect 73798 89876 73804 89888
rect 73755 89848 73804 89876
rect 73755 89845 73767 89848
rect 73709 89839 73767 89845
rect 73798 89836 73804 89848
rect 73856 89836 73862 89888
rect 415210 89808 415216 89820
rect 415136 89780 415216 89808
rect 194778 89700 194784 89752
rect 194836 89700 194842 89752
rect 243722 89700 243728 89752
rect 243780 89700 243786 89752
rect 322566 89700 322572 89752
rect 322624 89740 322630 89752
rect 322750 89740 322756 89752
rect 322624 89712 322756 89740
rect 322624 89700 322630 89712
rect 322750 89700 322756 89712
rect 322808 89700 322814 89752
rect 394326 89700 394332 89752
rect 394384 89740 394390 89752
rect 394510 89740 394516 89752
rect 394384 89712 394516 89740
rect 394384 89700 394390 89712
rect 394510 89700 394516 89712
rect 394568 89700 394574 89752
rect 194796 89604 194824 89700
rect 227717 89675 227775 89681
rect 227717 89641 227729 89675
rect 227763 89672 227775 89675
rect 227806 89672 227812 89684
rect 227763 89644 227812 89672
rect 227763 89641 227775 89644
rect 227717 89635 227775 89641
rect 227806 89632 227812 89644
rect 227864 89632 227870 89684
rect 238846 89672 238852 89684
rect 238807 89644 238852 89672
rect 238846 89632 238852 89644
rect 238904 89632 238910 89684
rect 243740 89616 243768 89700
rect 415136 89684 415164 89780
rect 415210 89768 415216 89780
rect 415268 89768 415274 89820
rect 420638 89700 420644 89752
rect 420696 89700 420702 89752
rect 415118 89632 415124 89684
rect 415176 89632 415182 89684
rect 420656 89616 420684 89700
rect 194870 89604 194876 89616
rect 194796 89576 194876 89604
rect 194870 89564 194876 89576
rect 194928 89564 194934 89616
rect 243722 89564 243728 89616
rect 243780 89564 243786 89616
rect 420638 89564 420644 89616
rect 420696 89564 420702 89616
rect 179506 88992 179512 89004
rect 179467 88964 179512 88992
rect 179506 88952 179512 88964
rect 179564 88952 179570 89004
rect 131390 88272 131396 88324
rect 131448 88312 131454 88324
rect 580166 88312 580172 88324
rect 131448 88284 580172 88312
rect 131448 88272 131454 88284
rect 580166 88272 580172 88284
rect 580224 88272 580230 88324
rect 248230 87116 248236 87168
rect 248288 87156 248294 87168
rect 248288 87128 248368 87156
rect 248288 87116 248294 87128
rect 248340 87032 248368 87128
rect 73706 87020 73712 87032
rect 73667 86992 73712 87020
rect 73706 86980 73712 86992
rect 73764 86980 73770 87032
rect 233418 86980 233424 87032
rect 233476 87020 233482 87032
rect 233510 87020 233516 87032
rect 233476 86992 233516 87020
rect 233476 86980 233482 86992
rect 233510 86980 233516 86992
rect 233568 86980 233574 87032
rect 248322 86980 248328 87032
rect 248380 86980 248386 87032
rect 271874 86980 271880 87032
rect 271932 86980 271938 87032
rect 383102 87020 383108 87032
rect 383063 86992 383108 87020
rect 383102 86980 383108 86992
rect 383160 86980 383166 87032
rect 388622 87020 388628 87032
rect 388583 86992 388628 87020
rect 388622 86980 388628 86992
rect 388680 86980 388686 87032
rect 403894 87020 403900 87032
rect 403855 86992 403900 87020
rect 403894 86980 403900 86992
rect 403952 86980 403958 87032
rect 183738 86912 183744 86964
rect 183796 86952 183802 86964
rect 183922 86952 183928 86964
rect 183796 86924 183928 86952
rect 183796 86912 183802 86924
rect 183922 86912 183928 86924
rect 183980 86912 183986 86964
rect 190730 86952 190736 86964
rect 190691 86924 190736 86952
rect 190730 86912 190736 86924
rect 190788 86912 190794 86964
rect 243722 86952 243728 86964
rect 243683 86924 243728 86952
rect 243722 86912 243728 86924
rect 243780 86912 243786 86964
rect 245749 86955 245807 86961
rect 245749 86921 245761 86955
rect 245795 86952 245807 86955
rect 245930 86952 245936 86964
rect 245795 86924 245936 86952
rect 245795 86921 245807 86924
rect 245749 86915 245807 86921
rect 245930 86912 245936 86924
rect 245988 86912 245994 86964
rect 271892 86896 271920 86980
rect 274821 86955 274879 86961
rect 274821 86921 274833 86955
rect 274867 86952 274879 86955
rect 274910 86952 274916 86964
rect 274867 86924 274916 86952
rect 274867 86921 274879 86924
rect 274821 86915 274879 86921
rect 274910 86912 274916 86924
rect 274968 86912 274974 86964
rect 322658 86952 322664 86964
rect 322619 86924 322664 86952
rect 322658 86912 322664 86924
rect 322716 86912 322722 86964
rect 394418 86952 394424 86964
rect 394379 86924 394424 86952
rect 394418 86912 394424 86924
rect 394476 86912 394482 86964
rect 233418 86884 233424 86896
rect 233379 86856 233424 86884
rect 233418 86844 233424 86856
rect 233476 86844 233482 86896
rect 271874 86844 271880 86896
rect 271932 86844 271938 86896
rect 150618 85660 150624 85672
rect 150544 85632 150624 85660
rect 150544 85604 150572 85632
rect 150618 85620 150624 85632
rect 150676 85620 150682 85672
rect 144914 85592 144920 85604
rect 144875 85564 144920 85592
rect 144914 85552 144920 85564
rect 144972 85552 144978 85604
rect 150526 85552 150532 85604
rect 150584 85552 150590 85604
rect 426158 85592 426164 85604
rect 426119 85564 426164 85592
rect 426158 85552 426164 85564
rect 426216 85552 426222 85604
rect 194870 85524 194876 85536
rect 194831 85496 194876 85524
rect 194870 85484 194876 85496
rect 194928 85484 194934 85536
rect 200298 85524 200304 85536
rect 200259 85496 200304 85524
rect 200298 85484 200304 85496
rect 200356 85484 200362 85536
rect 248322 85524 248328 85536
rect 248283 85496 248328 85524
rect 248322 85484 248328 85496
rect 248380 85484 248386 85536
rect 325694 85524 325700 85536
rect 325655 85496 325700 85524
rect 325694 85484 325700 85496
rect 325752 85484 325758 85536
rect 279694 84300 279700 84312
rect 279655 84272 279700 84300
rect 279694 84260 279700 84272
rect 279752 84260 279758 84312
rect 156049 84235 156107 84241
rect 156049 84201 156061 84235
rect 156095 84232 156107 84235
rect 156138 84232 156144 84244
rect 156095 84204 156144 84232
rect 156095 84201 156107 84204
rect 156049 84195 156107 84201
rect 156138 84192 156144 84204
rect 156196 84192 156202 84244
rect 179509 84235 179567 84241
rect 179509 84201 179521 84235
rect 179555 84232 179567 84235
rect 179598 84232 179604 84244
rect 179555 84204 179604 84232
rect 179555 84201 179567 84204
rect 179509 84195 179567 84201
rect 179598 84192 179604 84204
rect 179656 84192 179662 84244
rect 162854 84164 162860 84176
rect 162815 84136 162860 84164
rect 162854 84124 162860 84136
rect 162912 84124 162918 84176
rect 279694 84164 279700 84176
rect 279655 84136 279700 84164
rect 279694 84124 279700 84136
rect 279752 84124 279758 84176
rect 426069 84167 426127 84173
rect 426069 84133 426081 84167
rect 426115 84164 426127 84167
rect 426158 84164 426164 84176
rect 426115 84136 426164 84164
rect 426115 84133 426127 84136
rect 426069 84127 426127 84133
rect 426158 84124 426164 84136
rect 426216 84124 426222 84176
rect 181165 82875 181223 82881
rect 181165 82841 181177 82875
rect 181211 82872 181223 82875
rect 181254 82872 181260 82884
rect 181211 82844 181260 82872
rect 181211 82841 181223 82844
rect 181165 82835 181223 82841
rect 181254 82832 181260 82844
rect 181312 82832 181318 82884
rect 227898 82124 227904 82136
rect 227859 82096 227904 82124
rect 227898 82084 227904 82096
rect 227956 82084 227962 82136
rect 420270 82084 420276 82136
rect 420328 82124 420334 82136
rect 420638 82124 420644 82136
rect 420328 82096 420644 82124
rect 420328 82084 420334 82096
rect 420638 82084 420644 82096
rect 420696 82084 420702 82136
rect 205910 81404 205916 81456
rect 205968 81444 205974 81456
rect 206094 81444 206100 81456
rect 205968 81416 206100 81444
rect 205968 81404 205974 81416
rect 206094 81404 206100 81416
rect 206152 81404 206158 81456
rect 207109 81447 207167 81453
rect 207109 81413 207121 81447
rect 207155 81444 207167 81447
rect 207198 81444 207204 81456
rect 207155 81416 207204 81444
rect 207155 81413 207167 81416
rect 207109 81407 207167 81413
rect 207198 81404 207204 81416
rect 207256 81404 207262 81456
rect 211338 81404 211344 81456
rect 211396 81444 211402 81456
rect 211430 81444 211436 81456
rect 211396 81416 211436 81444
rect 211396 81404 211402 81416
rect 211430 81404 211436 81416
rect 211488 81404 211494 81456
rect 238938 81444 238944 81456
rect 238899 81416 238944 81444
rect 238938 81404 238944 81416
rect 238996 81404 239002 81456
rect 150526 80724 150532 80776
rect 150584 80764 150590 80776
rect 150710 80764 150716 80776
rect 150584 80736 150716 80764
rect 150584 80724 150590 80736
rect 150710 80724 150716 80736
rect 150768 80724 150774 80776
rect 205910 80152 205916 80164
rect 205871 80124 205916 80152
rect 205910 80112 205916 80124
rect 205968 80112 205974 80164
rect 207198 80152 207204 80164
rect 207159 80124 207204 80152
rect 207198 80112 207204 80124
rect 207256 80112 207262 80164
rect 221001 80155 221059 80161
rect 221001 80121 221013 80155
rect 221047 80152 221059 80155
rect 221090 80152 221096 80164
rect 221047 80124 221096 80152
rect 221047 80121 221059 80124
rect 221001 80115 221059 80121
rect 221090 80112 221096 80124
rect 221148 80112 221154 80164
rect 229278 80152 229284 80164
rect 229204 80124 229284 80152
rect 229204 80096 229232 80124
rect 229278 80112 229284 80124
rect 229336 80112 229342 80164
rect 357986 80152 357992 80164
rect 357947 80124 357992 80152
rect 357986 80112 357992 80124
rect 358044 80112 358050 80164
rect 229186 80044 229192 80096
rect 229244 80044 229250 80096
rect 431586 80044 431592 80096
rect 431644 80084 431650 80096
rect 431770 80084 431776 80096
rect 431644 80056 431776 80084
rect 431644 80044 431650 80056
rect 431770 80044 431776 80056
rect 431828 80044 431834 80096
rect 3234 79976 3240 80028
rect 3292 80016 3298 80028
rect 434990 80016 434996 80028
rect 3292 79988 434996 80016
rect 3292 79976 3298 79988
rect 434990 79976 434996 79988
rect 435048 79976 435054 80028
rect 220998 79948 221004 79960
rect 220959 79920 221004 79948
rect 220998 79908 221004 79920
rect 221056 79908 221062 79960
rect 357986 79948 357992 79960
rect 357947 79920 357992 79948
rect 357986 79908 357992 79920
rect 358044 79908 358050 79960
rect 184842 77364 184848 77376
rect 184803 77336 184848 77364
rect 184842 77324 184848 77336
rect 184900 77324 184906 77376
rect 301866 77324 301872 77376
rect 301924 77364 301930 77376
rect 302050 77364 302056 77376
rect 301924 77336 302056 77364
rect 301924 77324 301930 77336
rect 302050 77324 302056 77336
rect 302108 77324 302114 77376
rect 128814 77256 128820 77308
rect 128872 77296 128878 77308
rect 128998 77296 129004 77308
rect 128872 77268 129004 77296
rect 128872 77256 128878 77268
rect 128998 77256 129004 77268
rect 129056 77256 129062 77308
rect 190733 77299 190791 77305
rect 190733 77265 190745 77299
rect 190779 77296 190791 77299
rect 190822 77296 190828 77308
rect 190779 77268 190828 77296
rect 190779 77265 190791 77268
rect 190733 77259 190791 77265
rect 190822 77256 190828 77268
rect 190880 77256 190886 77308
rect 227901 77299 227959 77305
rect 227901 77265 227913 77299
rect 227947 77296 227959 77299
rect 227990 77296 227996 77308
rect 227947 77268 227996 77296
rect 227947 77265 227959 77268
rect 227901 77259 227959 77265
rect 227990 77256 227996 77268
rect 228048 77256 228054 77308
rect 233418 77296 233424 77308
rect 233379 77268 233424 77296
rect 233418 77256 233424 77268
rect 233476 77256 233482 77308
rect 238938 77296 238944 77308
rect 238899 77268 238944 77296
rect 238938 77256 238944 77268
rect 238996 77256 239002 77308
rect 243722 77296 243728 77308
rect 243683 77268 243728 77296
rect 243722 77256 243728 77268
rect 243780 77256 243786 77308
rect 245746 77296 245752 77308
rect 245707 77268 245752 77296
rect 245746 77256 245752 77268
rect 245804 77256 245810 77308
rect 274818 77296 274824 77308
rect 274779 77268 274824 77296
rect 274818 77256 274824 77268
rect 274876 77256 274882 77308
rect 322661 77299 322719 77305
rect 322661 77265 322673 77299
rect 322707 77296 322719 77299
rect 322750 77296 322756 77308
rect 322707 77268 322756 77296
rect 322707 77265 322719 77268
rect 322661 77259 322719 77265
rect 322750 77256 322756 77268
rect 322808 77256 322814 77308
rect 394421 77299 394479 77305
rect 394421 77265 394433 77299
rect 394467 77296 394479 77299
rect 394510 77296 394516 77308
rect 394467 77268 394516 77296
rect 394467 77265 394479 77268
rect 394421 77259 394479 77265
rect 394510 77256 394516 77268
rect 394568 77256 394574 77308
rect 132126 77188 132132 77240
rect 132184 77228 132190 77240
rect 580166 77228 580172 77240
rect 132184 77200 580172 77228
rect 132184 77188 132190 77200
rect 580166 77188 580172 77200
rect 580224 77188 580230 77240
rect 184842 77160 184848 77172
rect 184803 77132 184848 77160
rect 184842 77120 184848 77132
rect 184900 77120 184906 77172
rect 301961 77163 302019 77169
rect 301961 77129 301973 77163
rect 302007 77160 302019 77163
rect 302050 77160 302056 77172
rect 302007 77132 302056 77160
rect 302007 77129 302019 77132
rect 301961 77123 302019 77129
rect 302050 77120 302056 77132
rect 302108 77120 302114 77172
rect 341334 77160 341340 77172
rect 341295 77132 341340 77160
rect 341334 77120 341340 77132
rect 341392 77120 341398 77172
rect 383194 77160 383200 77172
rect 383155 77132 383200 77160
rect 383194 77120 383200 77132
rect 383252 77120 383258 77172
rect 388714 77160 388720 77172
rect 388675 77132 388720 77160
rect 388714 77120 388720 77132
rect 388772 77120 388778 77172
rect 403986 77160 403992 77172
rect 403947 77132 403992 77160
rect 403986 77120 403992 77132
rect 404044 77120 404050 77172
rect 184750 77052 184756 77104
rect 184808 77092 184814 77104
rect 185026 77092 185032 77104
rect 184808 77064 185032 77092
rect 184808 77052 184814 77064
rect 185026 77052 185032 77064
rect 185084 77052 185090 77104
rect 207198 76616 207204 76628
rect 207159 76588 207204 76616
rect 207198 76576 207204 76588
rect 207256 76576 207262 76628
rect 181254 76004 181260 76016
rect 181088 75976 181260 76004
rect 173986 75896 173992 75948
rect 174044 75936 174050 75948
rect 174078 75936 174084 75948
rect 174044 75908 174084 75936
rect 174044 75896 174050 75908
rect 174078 75896 174084 75908
rect 174136 75896 174142 75948
rect 181088 75880 181116 75976
rect 181254 75964 181260 75976
rect 181312 75964 181318 76016
rect 194870 75936 194876 75948
rect 194831 75908 194876 75936
rect 194870 75896 194876 75908
rect 194928 75896 194934 75948
rect 200298 75936 200304 75948
rect 200259 75908 200304 75936
rect 200298 75896 200304 75908
rect 200356 75896 200362 75948
rect 248322 75936 248328 75948
rect 248283 75908 248328 75936
rect 248322 75896 248328 75908
rect 248380 75896 248386 75948
rect 325694 75936 325700 75948
rect 325655 75908 325700 75936
rect 325694 75896 325700 75908
rect 325752 75896 325758 75948
rect 415026 75896 415032 75948
rect 415084 75936 415090 75948
rect 415118 75936 415124 75948
rect 415084 75908 415124 75936
rect 415084 75896 415090 75908
rect 415118 75896 415124 75908
rect 415176 75896 415182 75948
rect 157426 75868 157432 75880
rect 157387 75840 157432 75868
rect 157426 75828 157432 75840
rect 157484 75828 157490 75880
rect 178126 75828 178132 75880
rect 178184 75868 178190 75880
rect 178310 75868 178316 75880
rect 178184 75840 178316 75868
rect 178184 75828 178190 75840
rect 178310 75828 178316 75840
rect 178368 75828 178374 75880
rect 181070 75828 181076 75880
rect 181128 75828 181134 75880
rect 183741 75871 183799 75877
rect 183741 75837 183753 75871
rect 183787 75868 183799 75871
rect 183922 75868 183928 75880
rect 183787 75840 183928 75868
rect 183787 75837 183799 75840
rect 183741 75831 183799 75837
rect 183922 75828 183928 75840
rect 183980 75828 183986 75880
rect 211249 75871 211307 75877
rect 211249 75837 211261 75871
rect 211295 75868 211307 75871
rect 211338 75868 211344 75880
rect 211295 75840 211344 75868
rect 211295 75837 211307 75840
rect 211249 75831 211307 75837
rect 211338 75828 211344 75840
rect 211396 75828 211402 75880
rect 244274 75868 244280 75880
rect 244235 75840 244280 75868
rect 244274 75828 244280 75840
rect 244332 75828 244338 75880
rect 245746 75868 245752 75880
rect 245707 75840 245752 75868
rect 245746 75828 245752 75840
rect 245804 75828 245810 75880
rect 271874 75868 271880 75880
rect 271835 75840 271880 75868
rect 271874 75828 271880 75840
rect 271932 75828 271938 75880
rect 431586 75868 431592 75880
rect 431547 75840 431592 75868
rect 431586 75828 431592 75840
rect 431644 75828 431650 75880
rect 156046 74536 156052 74588
rect 156104 74576 156110 74588
rect 156230 74576 156236 74588
rect 156104 74548 156236 74576
rect 156104 74536 156110 74548
rect 156230 74536 156236 74548
rect 156288 74536 156294 74588
rect 162854 74576 162860 74588
rect 162815 74548 162860 74576
rect 162854 74536 162860 74548
rect 162912 74536 162918 74588
rect 279697 74579 279755 74585
rect 279697 74545 279709 74579
rect 279743 74576 279755 74579
rect 279786 74576 279792 74588
rect 279743 74548 279792 74576
rect 279743 74545 279755 74548
rect 279697 74539 279755 74545
rect 279786 74536 279792 74548
rect 279844 74536 279850 74588
rect 173989 74511 174047 74517
rect 173989 74477 174001 74511
rect 174035 74508 174047 74511
rect 174078 74508 174084 74520
rect 174035 74480 174084 74508
rect 174035 74477 174047 74480
rect 173989 74471 174047 74477
rect 174078 74468 174084 74480
rect 174136 74468 174142 74520
rect 205910 74100 205916 74112
rect 205871 74072 205916 74100
rect 205910 74060 205916 74072
rect 205968 74060 205974 74112
rect 212810 73284 212816 73296
rect 212736 73256 212816 73284
rect 212736 73228 212764 73256
rect 212810 73244 212816 73256
rect 212868 73244 212874 73296
rect 212718 73176 212724 73228
rect 212776 73176 212782 73228
rect 181070 73148 181076 73160
rect 181031 73120 181076 73148
rect 181070 73108 181076 73120
rect 181128 73108 181134 73160
rect 150710 70496 150716 70508
rect 150636 70468 150716 70496
rect 150636 70372 150664 70468
rect 150710 70456 150716 70468
rect 150768 70456 150774 70508
rect 194870 70496 194876 70508
rect 194796 70468 194876 70496
rect 194796 70372 194824 70468
rect 194870 70456 194876 70468
rect 194928 70456 194934 70508
rect 209866 70496 209872 70508
rect 209827 70468 209872 70496
rect 209866 70456 209872 70468
rect 209924 70456 209930 70508
rect 240226 70496 240232 70508
rect 240187 70468 240232 70496
rect 240226 70456 240232 70468
rect 240284 70456 240290 70508
rect 279786 70388 279792 70440
rect 279844 70388 279850 70440
rect 150618 70320 150624 70372
rect 150676 70320 150682 70372
rect 194778 70320 194784 70372
rect 194836 70320 194842 70372
rect 279804 70304 279832 70388
rect 271877 70295 271935 70301
rect 271877 70261 271889 70295
rect 271923 70292 271935 70295
rect 271966 70292 271972 70304
rect 271923 70264 271972 70292
rect 271923 70261 271935 70264
rect 271877 70255 271935 70261
rect 271966 70252 271972 70264
rect 272024 70252 272030 70304
rect 279786 70252 279792 70304
rect 279844 70252 279850 70304
rect 426066 69680 426072 69692
rect 426027 69652 426072 69680
rect 426066 69640 426072 69652
rect 426124 69640 426130 69692
rect 212718 68388 212724 68400
rect 212679 68360 212724 68388
rect 212718 68348 212724 68360
rect 212776 68348 212782 68400
rect 128722 67668 128728 67720
rect 128780 67668 128786 67720
rect 190822 67708 190828 67720
rect 190748 67680 190828 67708
rect 128740 67640 128768 67668
rect 190748 67652 190776 67680
rect 190822 67668 190828 67680
rect 190880 67668 190886 67720
rect 234706 67708 234712 67720
rect 234667 67680 234712 67708
rect 234706 67668 234712 67680
rect 234764 67668 234770 67720
rect 128906 67640 128912 67652
rect 128740 67612 128912 67640
rect 128906 67600 128912 67612
rect 128964 67600 128970 67652
rect 184750 67600 184756 67652
rect 184808 67640 184814 67652
rect 184934 67640 184940 67652
rect 184808 67612 184940 67640
rect 184808 67600 184814 67612
rect 184934 67600 184940 67612
rect 184992 67600 184998 67652
rect 190730 67600 190736 67652
rect 190788 67600 190794 67652
rect 200298 67600 200304 67652
rect 200356 67640 200362 67652
rect 200390 67640 200396 67652
rect 200356 67612 200396 67640
rect 200356 67600 200362 67612
rect 200390 67600 200396 67612
rect 200448 67600 200454 67652
rect 209866 67640 209872 67652
rect 209827 67612 209872 67640
rect 209866 67600 209872 67612
rect 209924 67600 209930 67652
rect 240226 67640 240232 67652
rect 240187 67612 240232 67640
rect 240226 67600 240232 67612
rect 240284 67600 240290 67652
rect 301958 67640 301964 67652
rect 301919 67612 301964 67640
rect 301958 67600 301964 67612
rect 302016 67600 302022 67652
rect 341337 67643 341395 67649
rect 341337 67609 341349 67643
rect 341383 67640 341395 67643
rect 341426 67640 341432 67652
rect 341383 67612 341432 67640
rect 341383 67609 341395 67612
rect 341337 67603 341395 67609
rect 341426 67600 341432 67612
rect 341484 67600 341490 67652
rect 383197 67643 383255 67649
rect 383197 67609 383209 67643
rect 383243 67640 383255 67643
rect 383286 67640 383292 67652
rect 383243 67612 383292 67640
rect 383243 67609 383255 67612
rect 383197 67603 383255 67609
rect 383286 67600 383292 67612
rect 383344 67600 383350 67652
rect 388717 67643 388775 67649
rect 388717 67609 388729 67643
rect 388763 67640 388775 67643
rect 388806 67640 388812 67652
rect 388763 67612 388812 67640
rect 388763 67609 388775 67612
rect 388717 67603 388775 67609
rect 388806 67600 388812 67612
rect 388864 67600 388870 67652
rect 394418 67600 394424 67652
rect 394476 67640 394482 67652
rect 394510 67640 394516 67652
rect 394476 67612 394516 67640
rect 394476 67600 394482 67612
rect 394510 67600 394516 67612
rect 394568 67600 394574 67652
rect 403989 67643 404047 67649
rect 403989 67609 404001 67643
rect 404035 67640 404047 67643
rect 404078 67640 404084 67652
rect 404035 67612 404084 67640
rect 404035 67609 404047 67612
rect 403989 67603 404047 67609
rect 404078 67600 404084 67612
rect 404136 67600 404142 67652
rect 233418 67572 233424 67584
rect 233379 67544 233424 67572
rect 233418 67532 233424 67544
rect 233476 67532 233482 67584
rect 145098 66308 145104 66360
rect 145156 66348 145162 66360
rect 145282 66348 145288 66360
rect 145156 66320 145288 66348
rect 145156 66308 145162 66320
rect 145282 66308 145288 66320
rect 145340 66308 145346 66360
rect 183738 66348 183744 66360
rect 183699 66320 183744 66348
rect 183738 66308 183744 66320
rect 183796 66308 183802 66360
rect 73798 66240 73804 66292
rect 73856 66280 73862 66292
rect 73890 66280 73896 66292
rect 73856 66252 73896 66280
rect 73856 66240 73862 66252
rect 73890 66240 73896 66252
rect 73948 66240 73954 66292
rect 157426 66280 157432 66292
rect 157387 66252 157432 66280
rect 157426 66240 157432 66252
rect 157484 66240 157490 66292
rect 179506 66240 179512 66292
rect 179564 66280 179570 66292
rect 179598 66280 179604 66292
rect 179564 66252 179604 66280
rect 179564 66240 179570 66252
rect 179598 66240 179604 66252
rect 179656 66240 179662 66292
rect 211246 66280 211252 66292
rect 211207 66252 211252 66280
rect 211246 66240 211252 66252
rect 211304 66240 211310 66292
rect 234706 66280 234712 66292
rect 234667 66252 234712 66280
rect 234706 66240 234712 66252
rect 234764 66240 234770 66292
rect 244277 66283 244335 66289
rect 244277 66249 244289 66283
rect 244323 66280 244335 66283
rect 244366 66280 244372 66292
rect 244323 66252 244372 66280
rect 244323 66249 244335 66252
rect 244277 66243 244335 66249
rect 244366 66240 244372 66252
rect 244424 66240 244430 66292
rect 245749 66283 245807 66289
rect 245749 66249 245761 66283
rect 245795 66280 245807 66283
rect 245838 66280 245844 66292
rect 245795 66252 245844 66280
rect 245795 66249 245807 66252
rect 245749 66243 245807 66249
rect 245838 66240 245844 66252
rect 245896 66240 245902 66292
rect 322658 66240 322664 66292
rect 322716 66280 322722 66292
rect 322750 66280 322756 66292
rect 322716 66252 322756 66280
rect 322716 66240 322722 66252
rect 322750 66240 322756 66252
rect 322808 66240 322814 66292
rect 420454 66240 420460 66292
rect 420512 66280 420518 66292
rect 420546 66280 420552 66292
rect 420512 66252 420552 66280
rect 420512 66240 420518 66252
rect 420546 66240 420552 66252
rect 420604 66240 420610 66292
rect 431586 66280 431592 66292
rect 431547 66252 431592 66280
rect 431586 66240 431592 66252
rect 431644 66240 431650 66292
rect 128906 66212 128912 66224
rect 128867 66184 128912 66212
rect 128906 66172 128912 66184
rect 128964 66172 128970 66224
rect 183738 66212 183744 66224
rect 183699 66184 183744 66212
rect 183738 66172 183744 66184
rect 183796 66172 183802 66224
rect 190730 66172 190736 66224
rect 190788 66212 190794 66224
rect 190822 66212 190828 66224
rect 190788 66184 190828 66212
rect 190788 66172 190794 66184
rect 190822 66172 190828 66184
rect 190880 66172 190886 66224
rect 194778 66172 194784 66224
rect 194836 66212 194842 66224
rect 195149 66215 195207 66221
rect 195149 66212 195161 66215
rect 194836 66184 195161 66212
rect 194836 66172 194842 66184
rect 195149 66181 195161 66184
rect 195195 66181 195207 66215
rect 195149 66175 195207 66181
rect 207109 66215 207167 66221
rect 207109 66181 207121 66215
rect 207155 66212 207167 66215
rect 207198 66212 207204 66224
rect 207155 66184 207204 66212
rect 207155 66181 207167 66184
rect 207109 66175 207167 66181
rect 207198 66172 207204 66184
rect 207256 66172 207262 66224
rect 248322 66212 248328 66224
rect 248283 66184 248328 66212
rect 248322 66172 248328 66184
rect 248380 66172 248386 66224
rect 325513 66215 325571 66221
rect 325513 66181 325525 66215
rect 325559 66212 325571 66215
rect 325694 66212 325700 66224
rect 325559 66184 325700 66212
rect 325559 66181 325571 66184
rect 325513 66175 325571 66181
rect 325694 66172 325700 66184
rect 325752 66172 325758 66224
rect 415026 66212 415032 66224
rect 414987 66184 415032 66212
rect 415026 66172 415032 66184
rect 415084 66172 415090 66224
rect 420454 66104 420460 66156
rect 420512 66144 420518 66156
rect 420638 66144 420644 66156
rect 420512 66116 420644 66144
rect 420512 66104 420518 66116
rect 420638 66104 420644 66116
rect 420696 66104 420702 66156
rect 173986 64920 173992 64932
rect 173947 64892 173992 64920
rect 173986 64880 173992 64892
rect 174044 64880 174050 64932
rect 3326 64812 3332 64864
rect 3384 64852 3390 64864
rect 131666 64852 131672 64864
rect 3384 64824 131672 64852
rect 3384 64812 3390 64824
rect 131666 64812 131672 64824
rect 131724 64812 131730 64864
rect 145098 64852 145104 64864
rect 145059 64824 145104 64852
rect 145098 64812 145104 64824
rect 145156 64812 145162 64864
rect 147950 64852 147956 64864
rect 147911 64824 147956 64852
rect 147950 64812 147956 64824
rect 148008 64812 148014 64864
rect 159082 64852 159088 64864
rect 159043 64824 159088 64852
rect 159082 64812 159088 64824
rect 159140 64812 159146 64864
rect 162854 64812 162860 64864
rect 162912 64852 162918 64864
rect 163130 64852 163136 64864
rect 162912 64824 163136 64852
rect 162912 64812 162918 64824
rect 163130 64812 163136 64824
rect 163188 64812 163194 64864
rect 178126 64812 178132 64864
rect 178184 64852 178190 64864
rect 178310 64852 178316 64864
rect 178184 64824 178316 64852
rect 178184 64812 178190 64824
rect 178310 64812 178316 64824
rect 178368 64812 178374 64864
rect 436830 64812 436836 64864
rect 436888 64852 436894 64864
rect 579798 64852 579804 64864
rect 436888 64824 579804 64852
rect 436888 64812 436894 64824
rect 579798 64812 579804 64824
rect 579856 64812 579862 64864
rect 181070 63560 181076 63572
rect 181031 63532 181076 63560
rect 181070 63520 181076 63532
rect 181128 63520 181134 63572
rect 233418 62812 233424 62824
rect 233379 62784 233424 62812
rect 233418 62772 233424 62784
rect 233476 62772 233482 62824
rect 181070 61004 181076 61056
rect 181128 61044 181134 61056
rect 181165 61047 181223 61053
rect 181165 61044 181177 61047
rect 181128 61016 181177 61044
rect 181128 61004 181134 61016
rect 181165 61013 181177 61016
rect 181211 61013 181223 61047
rect 181165 61007 181223 61013
rect 184934 60840 184940 60852
rect 184895 60812 184940 60840
rect 184934 60800 184940 60812
rect 184992 60800 184998 60852
rect 205821 60843 205879 60849
rect 205821 60809 205833 60843
rect 205867 60840 205879 60843
rect 205910 60840 205916 60852
rect 205867 60812 205916 60840
rect 205867 60809 205879 60812
rect 205821 60803 205879 60809
rect 205910 60800 205916 60812
rect 205968 60800 205974 60852
rect 227990 60840 227996 60852
rect 227916 60812 227996 60840
rect 227916 60784 227944 60812
rect 227990 60800 227996 60812
rect 228048 60800 228054 60852
rect 243722 60800 243728 60852
rect 243780 60800 243786 60852
rect 383286 60840 383292 60852
rect 383212 60812 383292 60840
rect 227898 60732 227904 60784
rect 227956 60732 227962 60784
rect 150526 60664 150532 60716
rect 150584 60704 150590 60716
rect 150710 60704 150716 60716
rect 150584 60676 150716 60704
rect 150584 60664 150590 60676
rect 150710 60664 150716 60676
rect 150768 60664 150774 60716
rect 156046 60664 156052 60716
rect 156104 60704 156110 60716
rect 156230 60704 156236 60716
rect 156104 60676 156236 60704
rect 156104 60664 156110 60676
rect 156230 60664 156236 60676
rect 156288 60664 156294 60716
rect 216766 60664 216772 60716
rect 216824 60704 216830 60716
rect 216950 60704 216956 60716
rect 216824 60676 216956 60704
rect 216824 60664 216830 60676
rect 216950 60664 216956 60676
rect 217008 60664 217014 60716
rect 220998 60664 221004 60716
rect 221056 60704 221062 60716
rect 221182 60704 221188 60716
rect 221056 60676 221188 60704
rect 221056 60664 221062 60676
rect 221182 60664 221188 60676
rect 221240 60664 221246 60716
rect 243740 60648 243768 60800
rect 383212 60716 383240 60812
rect 383286 60800 383292 60812
rect 383344 60800 383350 60852
rect 388806 60840 388812 60852
rect 388732 60812 388812 60840
rect 388732 60716 388760 60812
rect 388806 60800 388812 60812
rect 388864 60800 388870 60852
rect 404078 60840 404084 60852
rect 404004 60812 404084 60840
rect 404004 60716 404032 60812
rect 404078 60800 404084 60812
rect 404136 60800 404142 60852
rect 244366 60664 244372 60716
rect 244424 60704 244430 60716
rect 244550 60704 244556 60716
rect 244424 60676 244556 60704
rect 244424 60664 244430 60676
rect 244550 60664 244556 60676
rect 244608 60664 244614 60716
rect 245838 60664 245844 60716
rect 245896 60704 245902 60716
rect 246022 60704 246028 60716
rect 245896 60676 246028 60704
rect 245896 60664 245902 60676
rect 246022 60664 246028 60676
rect 246080 60664 246086 60716
rect 271966 60664 271972 60716
rect 272024 60704 272030 60716
rect 272150 60704 272156 60716
rect 272024 60676 272156 60704
rect 272024 60664 272030 60676
rect 272150 60664 272156 60676
rect 272208 60664 272214 60716
rect 279878 60664 279884 60716
rect 279936 60704 279942 60716
rect 280062 60704 280068 60716
rect 279936 60676 280068 60704
rect 279936 60664 279942 60676
rect 280062 60664 280068 60676
rect 280120 60664 280126 60716
rect 383194 60664 383200 60716
rect 383252 60664 383258 60716
rect 388714 60664 388720 60716
rect 388772 60664 388778 60716
rect 403986 60664 403992 60716
rect 404044 60664 404050 60716
rect 243722 60596 243728 60648
rect 243780 60596 243786 60648
rect 178218 59848 178224 59900
rect 178276 59888 178282 59900
rect 178310 59888 178316 59900
rect 178276 59860 178316 59888
rect 178276 59848 178282 59860
rect 178310 59848 178316 59860
rect 178368 59848 178374 59900
rect 240137 58055 240195 58061
rect 240137 58021 240149 58055
rect 240183 58052 240195 58055
rect 240226 58052 240232 58064
rect 240183 58024 240232 58052
rect 240183 58021 240195 58024
rect 240137 58015 240195 58021
rect 240226 58012 240232 58024
rect 240284 58012 240290 58064
rect 73890 57944 73896 57996
rect 73948 57984 73954 57996
rect 205818 57984 205824 57996
rect 73948 57956 74028 57984
rect 205779 57956 205824 57984
rect 73948 57944 73954 57956
rect 74000 57860 74028 57956
rect 205818 57944 205824 57956
rect 205876 57944 205882 57996
rect 133141 57919 133199 57925
rect 133141 57885 133153 57919
rect 133187 57916 133199 57919
rect 133230 57916 133236 57928
rect 133187 57888 133236 57916
rect 133187 57885 133199 57888
rect 133141 57879 133199 57885
rect 133230 57876 133236 57888
rect 133288 57876 133294 57928
rect 150710 57916 150716 57928
rect 150671 57888 150716 57916
rect 150710 57876 150716 57888
rect 150768 57876 150774 57928
rect 184934 57916 184940 57928
rect 184895 57888 184940 57916
rect 184934 57876 184940 57888
rect 184992 57876 184998 57928
rect 200301 57919 200359 57925
rect 200301 57885 200313 57919
rect 200347 57916 200359 57919
rect 200390 57916 200396 57928
rect 200347 57888 200396 57916
rect 200347 57885 200359 57888
rect 200301 57879 200359 57885
rect 200390 57876 200396 57888
rect 200448 57876 200454 57928
rect 212534 57876 212540 57928
rect 212592 57916 212598 57928
rect 212718 57916 212724 57928
rect 212592 57888 212637 57916
rect 212679 57888 212724 57916
rect 212592 57876 212598 57888
rect 212718 57876 212724 57888
rect 212776 57876 212782 57928
rect 216861 57919 216919 57925
rect 216861 57885 216873 57919
rect 216907 57916 216919 57919
rect 216950 57916 216956 57928
rect 216907 57888 216956 57916
rect 216907 57885 216919 57888
rect 216861 57879 216919 57885
rect 216950 57876 216956 57888
rect 217008 57876 217014 57928
rect 276106 57876 276112 57928
rect 276164 57916 276170 57928
rect 276290 57916 276296 57928
rect 276164 57888 276296 57916
rect 276164 57876 276170 57888
rect 276290 57876 276296 57888
rect 276348 57876 276354 57928
rect 279881 57919 279939 57925
rect 279881 57885 279893 57919
rect 279927 57916 279939 57919
rect 280062 57916 280068 57928
rect 279927 57888 280068 57916
rect 279927 57885 279939 57888
rect 279881 57879 279939 57885
rect 280062 57876 280068 57888
rect 280120 57876 280126 57928
rect 301774 57916 301780 57928
rect 301735 57888 301780 57916
rect 301774 57876 301780 57888
rect 301832 57876 301838 57928
rect 322661 57919 322719 57925
rect 322661 57885 322673 57919
rect 322707 57916 322719 57919
rect 322750 57916 322756 57928
rect 322707 57888 322756 57916
rect 322707 57885 322719 57888
rect 322661 57879 322719 57885
rect 322750 57876 322756 57888
rect 322808 57876 322814 57928
rect 383194 57916 383200 57928
rect 383155 57888 383200 57916
rect 383194 57876 383200 57888
rect 383252 57876 383258 57928
rect 388714 57916 388720 57928
rect 388675 57888 388720 57916
rect 388714 57876 388720 57888
rect 388772 57876 388778 57928
rect 403986 57916 403992 57928
rect 403947 57888 403992 57916
rect 403986 57876 403992 57888
rect 404044 57876 404050 57928
rect 73982 57808 73988 57860
rect 74040 57808 74046 57860
rect 128909 57851 128967 57857
rect 128909 57817 128921 57851
rect 128955 57848 128967 57851
rect 128998 57848 129004 57860
rect 128955 57820 129004 57848
rect 128955 57817 128967 57820
rect 128909 57811 128967 57817
rect 128998 57808 129004 57820
rect 129056 57808 129062 57860
rect 183738 56624 183744 56636
rect 183699 56596 183744 56624
rect 183738 56584 183744 56596
rect 183796 56584 183802 56636
rect 195146 56584 195152 56636
rect 195204 56624 195210 56636
rect 207106 56624 207112 56636
rect 195204 56596 195249 56624
rect 207067 56596 207112 56624
rect 195204 56584 195210 56596
rect 207106 56584 207112 56596
rect 207164 56584 207170 56636
rect 240134 56584 240140 56636
rect 240192 56624 240198 56636
rect 248322 56624 248328 56636
rect 240192 56596 240237 56624
rect 248283 56596 248328 56624
rect 240192 56584 240198 56596
rect 248322 56584 248328 56596
rect 248380 56584 248386 56636
rect 325510 56624 325516 56636
rect 325471 56596 325516 56624
rect 325510 56584 325516 56596
rect 325568 56584 325574 56636
rect 415026 56624 415032 56636
rect 414987 56596 415032 56624
rect 415026 56584 415032 56596
rect 415084 56584 415090 56636
rect 145098 56556 145104 56568
rect 145059 56528 145104 56556
rect 145098 56516 145104 56528
rect 145156 56516 145162 56568
rect 234706 56556 234712 56568
rect 234667 56528 234712 56556
rect 234706 56516 234712 56528
rect 234764 56516 234770 56568
rect 431586 56516 431592 56568
rect 431644 56556 431650 56568
rect 431770 56556 431776 56568
rect 431644 56528 431776 56556
rect 431644 56516 431650 56528
rect 431770 56516 431776 56528
rect 431828 56516 431834 56568
rect 147950 55264 147956 55276
rect 147911 55236 147956 55264
rect 147950 55224 147956 55236
rect 148008 55224 148014 55276
rect 159082 55264 159088 55276
rect 159043 55236 159088 55264
rect 159082 55224 159088 55236
rect 159140 55224 159146 55276
rect 173986 55224 173992 55276
rect 174044 55264 174050 55276
rect 174078 55264 174084 55276
rect 174044 55236 174084 55264
rect 174044 55224 174050 55236
rect 174078 55224 174084 55236
rect 174136 55224 174142 55276
rect 175642 55224 175648 55276
rect 175700 55264 175706 55276
rect 175826 55264 175832 55276
rect 175700 55236 175832 55264
rect 175700 55224 175706 55236
rect 175826 55224 175832 55236
rect 175884 55224 175890 55276
rect 227898 53156 227904 53168
rect 227859 53128 227904 53156
rect 227898 53116 227904 53128
rect 227956 53116 227962 53168
rect 238846 53116 238852 53168
rect 238904 53156 238910 53168
rect 239030 53156 239036 53168
rect 238904 53128 239036 53156
rect 238904 53116 238910 53128
rect 239030 53116 239036 53128
rect 239088 53116 239094 53168
rect 243446 53116 243452 53168
rect 243504 53156 243510 53168
rect 243722 53156 243728 53168
rect 243504 53128 243728 53156
rect 243504 53116 243510 53128
rect 243722 53116 243728 53128
rect 243780 53116 243786 53168
rect 426066 53116 426072 53168
rect 426124 53156 426130 53168
rect 426250 53156 426256 53168
rect 426124 53128 426256 53156
rect 426124 53116 426130 53128
rect 426250 53116 426256 53128
rect 426308 53116 426314 53168
rect 147950 51756 147956 51808
rect 148008 51796 148014 51808
rect 148134 51796 148140 51808
rect 148008 51768 148140 51796
rect 148008 51756 148014 51768
rect 148134 51756 148140 51768
rect 148192 51756 148198 51808
rect 415026 51280 415032 51332
rect 415084 51320 415090 51332
rect 415210 51320 415216 51332
rect 415084 51292 415216 51320
rect 415084 51280 415090 51292
rect 415210 51280 415216 51292
rect 415268 51280 415274 51332
rect 209866 51184 209872 51196
rect 209827 51156 209872 51184
rect 209866 51144 209872 51156
rect 209924 51144 209930 51196
rect 341518 51184 341524 51196
rect 341479 51156 341524 51184
rect 341518 51144 341524 51156
rect 341576 51144 341582 51196
rect 159082 51076 159088 51128
rect 159140 51076 159146 51128
rect 179506 51116 179512 51128
rect 179432 51088 179512 51116
rect 159100 50992 159128 51076
rect 179432 51060 179460 51088
rect 179506 51076 179512 51088
rect 179564 51076 179570 51128
rect 184934 51116 184940 51128
rect 184895 51088 184940 51116
rect 184934 51076 184940 51088
rect 184992 51076 184998 51128
rect 212534 51076 212540 51128
rect 212592 51116 212598 51128
rect 221182 51116 221188 51128
rect 212592 51088 212637 51116
rect 221108 51088 221188 51116
rect 212592 51076 212598 51088
rect 221108 51060 221136 51088
rect 221182 51076 221188 51088
rect 221240 51076 221246 51128
rect 244550 51116 244556 51128
rect 244476 51088 244556 51116
rect 244476 51060 244504 51088
rect 244550 51076 244556 51088
rect 244608 51076 244614 51128
rect 272150 51116 272156 51128
rect 272076 51088 272156 51116
rect 272076 51060 272104 51088
rect 272150 51076 272156 51088
rect 272208 51076 272214 51128
rect 179414 51008 179420 51060
rect 179472 51008 179478 51060
rect 221090 51008 221096 51060
rect 221148 51008 221154 51060
rect 244458 51008 244464 51060
rect 244516 51008 244522 51060
rect 272058 51008 272064 51060
rect 272116 51008 272122 51060
rect 357894 51008 357900 51060
rect 357952 51048 357958 51060
rect 358078 51048 358084 51060
rect 357952 51020 358084 51048
rect 357952 51008 357958 51020
rect 358078 51008 358084 51020
rect 358136 51008 358142 51060
rect 159082 50940 159088 50992
rect 159140 50940 159146 50992
rect 181162 50640 181168 50652
rect 181123 50612 181168 50640
rect 181162 50600 181168 50612
rect 181220 50600 181226 50652
rect 133138 48328 133144 48340
rect 133099 48300 133144 48328
rect 133138 48288 133144 48300
rect 133196 48288 133202 48340
rect 150713 48331 150771 48337
rect 150713 48297 150725 48331
rect 150759 48328 150771 48331
rect 150802 48328 150808 48340
rect 150759 48300 150808 48328
rect 150759 48297 150771 48300
rect 150713 48291 150771 48297
rect 150802 48288 150808 48300
rect 150860 48288 150866 48340
rect 184934 48328 184940 48340
rect 184895 48300 184940 48328
rect 184934 48288 184940 48300
rect 184992 48288 184998 48340
rect 200298 48328 200304 48340
rect 200259 48300 200304 48328
rect 200298 48288 200304 48300
rect 200356 48288 200362 48340
rect 216858 48328 216864 48340
rect 216819 48300 216864 48328
rect 216858 48288 216864 48300
rect 216916 48288 216922 48340
rect 227901 48331 227959 48337
rect 227901 48297 227913 48331
rect 227947 48328 227959 48331
rect 227990 48328 227996 48340
rect 227947 48300 227996 48328
rect 227947 48297 227959 48300
rect 227901 48291 227959 48297
rect 227990 48288 227996 48300
rect 228048 48288 228054 48340
rect 240134 48288 240140 48340
rect 240192 48328 240198 48340
rect 240226 48328 240232 48340
rect 240192 48300 240232 48328
rect 240192 48288 240198 48300
rect 240226 48288 240232 48300
rect 240284 48288 240290 48340
rect 248322 48328 248328 48340
rect 248283 48300 248328 48328
rect 248322 48288 248328 48300
rect 248380 48288 248386 48340
rect 279878 48328 279884 48340
rect 279839 48300 279884 48328
rect 279878 48288 279884 48300
rect 279936 48288 279942 48340
rect 301777 48331 301835 48337
rect 301777 48297 301789 48331
rect 301823 48328 301835 48331
rect 301866 48328 301872 48340
rect 301823 48300 301872 48328
rect 301823 48297 301835 48300
rect 301777 48291 301835 48297
rect 301866 48288 301872 48300
rect 301924 48288 301930 48340
rect 322658 48328 322664 48340
rect 322619 48300 322664 48328
rect 322658 48288 322664 48300
rect 322716 48288 322722 48340
rect 383197 48331 383255 48337
rect 383197 48297 383209 48331
rect 383243 48328 383255 48331
rect 383286 48328 383292 48340
rect 383243 48300 383292 48328
rect 383243 48297 383255 48300
rect 383197 48291 383255 48297
rect 383286 48288 383292 48300
rect 383344 48288 383350 48340
rect 388717 48331 388775 48337
rect 388717 48297 388729 48331
rect 388763 48328 388775 48331
rect 388806 48328 388812 48340
rect 388763 48300 388812 48328
rect 388763 48297 388775 48300
rect 388717 48291 388775 48297
rect 388806 48288 388812 48300
rect 388864 48288 388870 48340
rect 394418 48288 394424 48340
rect 394476 48328 394482 48340
rect 394510 48328 394516 48340
rect 394476 48300 394516 48328
rect 394476 48288 394482 48300
rect 394510 48288 394516 48300
rect 394568 48288 394574 48340
rect 403989 48331 404047 48337
rect 403989 48297 404001 48331
rect 404035 48328 404047 48331
rect 404078 48328 404084 48340
rect 404035 48300 404084 48328
rect 404035 48297 404047 48300
rect 403989 48291 404047 48297
rect 404078 48288 404084 48300
rect 404136 48288 404142 48340
rect 73614 48220 73620 48272
rect 73672 48260 73678 48272
rect 73801 48263 73859 48269
rect 73801 48260 73813 48263
rect 73672 48232 73813 48260
rect 73672 48220 73678 48232
rect 73801 48229 73813 48232
rect 73847 48229 73859 48263
rect 73801 48223 73859 48229
rect 357989 48263 358047 48269
rect 357989 48229 358001 48263
rect 358035 48260 358047 48263
rect 358078 48260 358084 48272
rect 358035 48232 358084 48260
rect 358035 48229 358047 48232
rect 357989 48223 358047 48229
rect 358078 48220 358084 48232
rect 358136 48220 358142 48272
rect 178218 47608 178224 47660
rect 178276 47648 178282 47660
rect 178402 47648 178408 47660
rect 178276 47620 178408 47648
rect 178276 47608 178282 47620
rect 178402 47608 178408 47620
rect 178460 47608 178466 47660
rect 207106 46996 207112 47048
rect 207164 46996 207170 47048
rect 207124 46968 207152 46996
rect 207198 46968 207204 46980
rect 207124 46940 207204 46968
rect 207198 46928 207204 46940
rect 207256 46928 207262 46980
rect 209866 46968 209872 46980
rect 209827 46940 209872 46968
rect 209866 46928 209872 46940
rect 209924 46928 209930 46980
rect 211246 46968 211252 46980
rect 211207 46940 211252 46968
rect 211246 46928 211252 46940
rect 211304 46928 211310 46980
rect 234706 46968 234712 46980
rect 234667 46940 234712 46968
rect 234706 46928 234712 46940
rect 234764 46928 234770 46980
rect 248322 46968 248328 46980
rect 248283 46940 248328 46968
rect 248322 46928 248328 46940
rect 248380 46928 248386 46980
rect 157337 46903 157395 46909
rect 157337 46869 157349 46903
rect 157383 46900 157395 46903
rect 157426 46900 157432 46912
rect 157383 46872 157432 46900
rect 157383 46869 157395 46872
rect 157337 46863 157395 46869
rect 157426 46860 157432 46872
rect 157484 46860 157490 46912
rect 190733 46903 190791 46909
rect 190733 46869 190745 46903
rect 190779 46900 190791 46903
rect 190822 46900 190828 46912
rect 190779 46872 190828 46900
rect 190779 46869 190791 46872
rect 190733 46863 190791 46869
rect 190822 46860 190828 46872
rect 190880 46860 190886 46912
rect 194689 46903 194747 46909
rect 194689 46869 194701 46903
rect 194735 46900 194747 46903
rect 194962 46900 194968 46912
rect 194735 46872 194968 46900
rect 194735 46869 194747 46872
rect 194689 46863 194747 46869
rect 194962 46860 194968 46872
rect 195020 46860 195026 46912
rect 276106 46900 276112 46912
rect 276067 46872 276112 46900
rect 276106 46860 276112 46872
rect 276164 46860 276170 46912
rect 325694 46900 325700 46912
rect 325655 46872 325700 46900
rect 325694 46860 325700 46872
rect 325752 46860 325758 46912
rect 420454 46860 420460 46912
rect 420512 46900 420518 46912
rect 420638 46900 420644 46912
rect 420512 46872 420644 46900
rect 420512 46860 420518 46872
rect 420638 46860 420644 46872
rect 420696 46860 420702 46912
rect 425974 46900 425980 46912
rect 425935 46872 425980 46900
rect 425974 46860 425980 46872
rect 426032 46860 426038 46912
rect 431586 46900 431592 46912
rect 431547 46872 431592 46900
rect 431586 46860 431592 46872
rect 431644 46860 431650 46912
rect 238846 45880 238852 45892
rect 238807 45852 238852 45880
rect 238846 45840 238852 45852
rect 238904 45840 238910 45892
rect 211246 45608 211252 45620
rect 211207 45580 211252 45608
rect 211246 45568 211252 45580
rect 211304 45568 211310 45620
rect 341518 45608 341524 45620
rect 341479 45580 341524 45608
rect 341518 45568 341524 45580
rect 341576 45568 341582 45620
rect 207198 45540 207204 45552
rect 207159 45512 207204 45540
rect 207198 45500 207204 45512
rect 207256 45500 207262 45552
rect 414934 45540 414940 45552
rect 414895 45512 414940 45540
rect 414934 45500 414940 45512
rect 414992 45500 414998 45552
rect 341429 45475 341487 45481
rect 341429 45441 341441 45475
rect 341475 45472 341487 45475
rect 341518 45472 341524 45484
rect 341475 45444 341524 45472
rect 341475 45441 341487 45444
rect 341429 45435 341487 45441
rect 341518 45432 341524 45444
rect 341576 45432 341582 45484
rect 181162 44112 181168 44124
rect 181123 44084 181168 44112
rect 181162 44072 181168 44084
rect 181220 44072 181226 44124
rect 147858 42032 147864 42084
rect 147916 42072 147922 42084
rect 148134 42072 148140 42084
rect 147916 42044 148140 42072
rect 147916 42032 147922 42044
rect 148134 42032 148140 42044
rect 148192 42032 148198 42084
rect 243446 41828 243452 41880
rect 243504 41868 243510 41880
rect 243814 41868 243820 41880
rect 243504 41840 243820 41868
rect 243504 41828 243510 41840
rect 243814 41828 243820 41840
rect 243872 41828 243878 41880
rect 150802 41460 150808 41472
rect 150763 41432 150808 41460
rect 150802 41420 150808 41432
rect 150860 41420 150866 41472
rect 133598 41352 133604 41404
rect 133656 41392 133662 41404
rect 580166 41392 580172 41404
rect 133656 41364 580172 41392
rect 133656 41352 133662 41364
rect 580166 41352 580172 41364
rect 580224 41352 580230 41404
rect 238849 41327 238907 41333
rect 238849 41293 238861 41327
rect 238895 41324 238907 41327
rect 238938 41324 238944 41336
rect 238895 41296 238944 41324
rect 238895 41293 238907 41296
rect 238849 41287 238907 41293
rect 238938 41284 238944 41296
rect 238996 41284 239002 41336
rect 211338 40672 211344 40724
rect 211396 40712 211402 40724
rect 211522 40712 211528 40724
rect 211396 40684 211528 40712
rect 211396 40672 211402 40684
rect 211522 40672 211528 40684
rect 211580 40672 211586 40724
rect 173894 39312 173900 39364
rect 173952 39352 173958 39364
rect 174078 39352 174084 39364
rect 173952 39324 174084 39352
rect 173952 39312 173958 39324
rect 174078 39312 174084 39324
rect 174136 39312 174142 39364
rect 212626 38632 212632 38684
rect 212684 38672 212690 38684
rect 212718 38672 212724 38684
rect 212684 38644 212724 38672
rect 212684 38632 212690 38644
rect 212718 38632 212724 38644
rect 212776 38632 212782 38684
rect 216674 38632 216680 38684
rect 216732 38672 216738 38684
rect 216766 38672 216772 38684
rect 216732 38644 216772 38672
rect 216732 38632 216738 38644
rect 216766 38632 216772 38644
rect 216824 38632 216830 38684
rect 220906 38632 220912 38684
rect 220964 38672 220970 38684
rect 221090 38672 221096 38684
rect 220964 38644 221096 38672
rect 220964 38632 220970 38644
rect 221090 38632 221096 38644
rect 221148 38632 221154 38684
rect 244274 38632 244280 38684
rect 244332 38672 244338 38684
rect 244366 38672 244372 38684
rect 244332 38644 244372 38672
rect 244332 38632 244338 38644
rect 244366 38632 244372 38644
rect 244424 38632 244430 38684
rect 245746 38632 245752 38684
rect 245804 38672 245810 38684
rect 245838 38672 245844 38684
rect 245804 38644 245844 38672
rect 245804 38632 245810 38644
rect 245838 38632 245844 38644
rect 245896 38632 245902 38684
rect 357986 38672 357992 38684
rect 357947 38644 357992 38672
rect 357986 38632 357992 38644
rect 358044 38632 358050 38684
rect 128909 38607 128967 38613
rect 128909 38573 128921 38607
rect 128955 38604 128967 38607
rect 128998 38604 129004 38616
rect 128955 38576 129004 38604
rect 128955 38573 128967 38576
rect 128909 38567 128967 38573
rect 128998 38564 129004 38576
rect 129056 38564 129062 38616
rect 133141 38607 133199 38613
rect 133141 38573 133153 38607
rect 133187 38604 133199 38607
rect 133230 38604 133236 38616
rect 133187 38576 133236 38604
rect 133187 38573 133199 38576
rect 133141 38567 133199 38573
rect 133230 38564 133236 38576
rect 133288 38564 133294 38616
rect 150802 38604 150808 38616
rect 150763 38576 150808 38604
rect 150802 38564 150808 38576
rect 150860 38564 150866 38616
rect 200393 38607 200451 38613
rect 200393 38573 200405 38607
rect 200439 38604 200451 38607
rect 200482 38604 200488 38616
rect 200439 38576 200488 38604
rect 200439 38573 200451 38576
rect 200393 38567 200451 38573
rect 200482 38564 200488 38576
rect 200540 38564 200546 38616
rect 322661 38607 322719 38613
rect 322661 38573 322673 38607
rect 322707 38604 322719 38607
rect 322750 38604 322756 38616
rect 322707 38576 322756 38604
rect 322707 38573 322719 38576
rect 322661 38567 322719 38573
rect 322750 38564 322756 38576
rect 322808 38564 322814 38616
rect 383194 38604 383200 38616
rect 383155 38576 383200 38604
rect 383194 38564 383200 38576
rect 383252 38564 383258 38616
rect 403986 38604 403992 38616
rect 403947 38576 403992 38604
rect 403986 38564 403992 38576
rect 404044 38564 404050 38616
rect 341426 38264 341432 38276
rect 341387 38236 341432 38264
rect 341426 38224 341432 38236
rect 341484 38224 341490 38276
rect 157334 37312 157340 37324
rect 157295 37284 157340 37312
rect 157334 37272 157340 37284
rect 157392 37272 157398 37324
rect 194686 37312 194692 37324
rect 194647 37284 194692 37312
rect 194686 37272 194692 37284
rect 194744 37272 194750 37324
rect 276106 37312 276112 37324
rect 276067 37284 276112 37312
rect 276106 37272 276112 37284
rect 276164 37272 276170 37324
rect 425977 37315 426035 37321
rect 425977 37281 425989 37315
rect 426023 37312 426035 37315
rect 426066 37312 426072 37324
rect 426023 37284 426072 37312
rect 426023 37281 426035 37284
rect 425977 37275 426035 37281
rect 426066 37272 426072 37284
rect 426124 37272 426130 37324
rect 431586 37312 431592 37324
rect 431547 37284 431592 37312
rect 431586 37272 431592 37284
rect 431644 37272 431650 37324
rect 150713 37247 150771 37253
rect 150713 37213 150725 37247
rect 150759 37244 150771 37247
rect 150802 37244 150808 37256
rect 150759 37216 150808 37244
rect 150759 37213 150771 37216
rect 150713 37207 150771 37213
rect 150802 37204 150808 37216
rect 150860 37204 150866 37256
rect 234706 37244 234712 37256
rect 234667 37216 234712 37244
rect 234706 37204 234712 37216
rect 234764 37204 234770 37256
rect 238849 37247 238907 37253
rect 238849 37213 238861 37247
rect 238895 37244 238907 37247
rect 238938 37244 238944 37256
rect 238895 37216 238944 37244
rect 238895 37213 238907 37216
rect 238849 37207 238907 37213
rect 238938 37204 238944 37216
rect 238996 37204 239002 37256
rect 244274 37244 244280 37256
rect 244235 37216 244280 37244
rect 244274 37204 244280 37216
rect 244332 37204 244338 37256
rect 245746 37244 245752 37256
rect 245707 37216 245752 37244
rect 245746 37204 245752 37216
rect 245804 37204 245810 37256
rect 248322 37244 248328 37256
rect 248283 37216 248328 37244
rect 248322 37204 248328 37216
rect 248380 37204 248386 37256
rect 271874 37244 271880 37256
rect 271835 37216 271880 37244
rect 271874 37204 271880 37216
rect 271932 37204 271938 37256
rect 431586 37176 431592 37188
rect 431547 37148 431592 37176
rect 431586 37136 431592 37148
rect 431644 37136 431650 37188
rect 207198 35952 207204 35964
rect 207159 35924 207204 35952
rect 207198 35912 207204 35924
rect 207256 35912 207262 35964
rect 414937 35955 414995 35961
rect 414937 35921 414949 35955
rect 414983 35952 414995 35955
rect 415026 35952 415032 35964
rect 414983 35924 415032 35952
rect 414983 35921 414995 35924
rect 414937 35915 414995 35921
rect 415026 35912 415032 35924
rect 415084 35912 415090 35964
rect 3418 35844 3424 35896
rect 3476 35884 3482 35896
rect 436186 35884 436192 35896
rect 3476 35856 180840 35884
rect 3476 35844 3482 35856
rect 180812 35816 180840 35856
rect 183296 35856 436192 35884
rect 183296 35816 183324 35856
rect 436186 35844 436192 35856
rect 436244 35844 436250 35896
rect 180812 35788 183324 35816
rect 73798 35340 73804 35352
rect 73759 35312 73804 35340
rect 73798 35300 73804 35312
rect 73856 35300 73862 35352
rect 229186 31872 229192 31884
rect 229147 31844 229192 31872
rect 229186 31832 229192 31844
rect 229244 31832 229250 31884
rect 301958 31832 301964 31884
rect 302016 31832 302022 31884
rect 145006 31764 145012 31816
rect 145064 31804 145070 31816
rect 145190 31804 145196 31816
rect 145064 31776 145196 31804
rect 145064 31764 145070 31776
rect 145190 31764 145196 31776
rect 145248 31764 145254 31816
rect 178218 31696 178224 31748
rect 178276 31736 178282 31748
rect 178402 31736 178408 31748
rect 178276 31708 178408 31736
rect 178276 31696 178282 31708
rect 178402 31696 178408 31708
rect 178460 31696 178466 31748
rect 245749 31739 245807 31745
rect 245749 31705 245761 31739
rect 245795 31736 245807 31739
rect 245838 31736 245844 31748
rect 245795 31708 245844 31736
rect 245795 31705 245807 31708
rect 245749 31699 245807 31705
rect 245838 31696 245844 31708
rect 245896 31696 245902 31748
rect 279878 31696 279884 31748
rect 279936 31736 279942 31748
rect 280062 31736 280068 31748
rect 279936 31708 280068 31736
rect 279936 31696 279942 31708
rect 280062 31696 280068 31708
rect 280120 31696 280126 31748
rect 301976 31736 302004 31832
rect 302050 31736 302056 31748
rect 301976 31708 302056 31736
rect 302050 31696 302056 31708
rect 302108 31696 302114 31748
rect 388714 31696 388720 31748
rect 388772 31736 388778 31748
rect 388898 31736 388904 31748
rect 388772 31708 388904 31736
rect 388772 31696 388778 31708
rect 388898 31696 388904 31708
rect 388956 31696 388962 31748
rect 181162 31668 181168 31680
rect 181123 31640 181168 31668
rect 181162 31628 181168 31640
rect 181220 31628 181226 31680
rect 244277 31671 244335 31677
rect 244277 31637 244289 31671
rect 244323 31668 244335 31671
rect 244366 31668 244372 31680
rect 244323 31640 244372 31668
rect 244323 31637 244335 31640
rect 244277 31631 244335 31637
rect 244366 31628 244372 31640
rect 244424 31628 244430 31680
rect 341426 31628 341432 31680
rect 341484 31668 341490 31680
rect 341518 31668 341524 31680
rect 341484 31640 341524 31668
rect 341484 31628 341490 31640
rect 341518 31628 341524 31640
rect 341576 31628 341582 31680
rect 431589 31671 431647 31677
rect 431589 31637 431601 31671
rect 431635 31668 431647 31671
rect 431678 31668 431684 31680
rect 431635 31640 431684 31668
rect 431635 31637 431647 31640
rect 431589 31631 431647 31637
rect 431678 31628 431684 31640
rect 431736 31628 431742 31680
rect 133138 31056 133144 31068
rect 133099 31028 133144 31056
rect 133138 31016 133144 31028
rect 133196 31016 133202 31068
rect 132402 30268 132408 30320
rect 132460 30308 132466 30320
rect 580166 30308 580172 30320
rect 132460 30280 580172 30308
rect 132460 30268 132466 30280
rect 580166 30268 580172 30280
rect 580224 30268 580230 30320
rect 325694 29084 325700 29096
rect 325655 29056 325700 29084
rect 325694 29044 325700 29056
rect 325752 29044 325758 29096
rect 357713 29087 357771 29093
rect 357713 29053 357725 29087
rect 357759 29084 357771 29087
rect 357986 29084 357992 29096
rect 357759 29056 357992 29084
rect 357759 29053 357771 29056
rect 357713 29047 357771 29053
rect 357986 29044 357992 29056
rect 358044 29044 358050 29096
rect 128906 29016 128912 29028
rect 128867 28988 128912 29016
rect 128906 28976 128912 28988
rect 128964 28976 128970 29028
rect 157334 28976 157340 29028
rect 157392 29016 157398 29028
rect 157426 29016 157432 29028
rect 157392 28988 157432 29016
rect 157392 28976 157398 28988
rect 157426 28976 157432 28988
rect 157484 28976 157490 29028
rect 159082 28976 159088 29028
rect 159140 29016 159146 29028
rect 159266 29016 159272 29028
rect 159140 28988 159272 29016
rect 159140 28976 159146 28988
rect 159266 28976 159272 28988
rect 159324 28976 159330 29028
rect 190730 29016 190736 29028
rect 190691 28988 190736 29016
rect 190730 28976 190736 28988
rect 190788 28976 190794 29028
rect 200390 29016 200396 29028
rect 200351 28988 200396 29016
rect 200390 28976 200396 28988
rect 200448 28976 200454 29028
rect 229186 29016 229192 29028
rect 229147 28988 229192 29016
rect 229186 28976 229192 28988
rect 229244 28976 229250 29028
rect 322658 29016 322664 29028
rect 322619 28988 322664 29016
rect 322658 28976 322664 28988
rect 322716 28976 322722 29028
rect 383197 29019 383255 29025
rect 383197 28985 383209 29019
rect 383243 29016 383255 29019
rect 383286 29016 383292 29028
rect 383243 28988 383292 29016
rect 383243 28985 383255 28988
rect 383197 28979 383255 28985
rect 383286 28976 383292 28988
rect 383344 28976 383350 29028
rect 394418 28976 394424 29028
rect 394476 29016 394482 29028
rect 394510 29016 394516 29028
rect 394476 28988 394516 29016
rect 394476 28976 394482 28988
rect 394510 28976 394516 28988
rect 394568 28976 394574 29028
rect 403989 29019 404047 29025
rect 403989 28985 404001 29019
rect 404035 29016 404047 29019
rect 404078 29016 404084 29028
rect 404035 28988 404084 29016
rect 404035 28985 404047 28988
rect 403989 28979 404047 28985
rect 404078 28976 404084 28988
rect 404136 28976 404142 29028
rect 183738 28908 183744 28960
rect 183796 28908 183802 28960
rect 184937 28951 184995 28957
rect 184937 28917 184949 28951
rect 184983 28948 184995 28951
rect 185026 28948 185032 28960
rect 184983 28920 185032 28948
rect 184983 28917 184995 28920
rect 184937 28911 184995 28917
rect 185026 28908 185032 28920
rect 185084 28908 185090 28960
rect 207198 28908 207204 28960
rect 207256 28948 207262 28960
rect 207290 28948 207296 28960
rect 207256 28920 207296 28948
rect 207256 28908 207262 28920
rect 207290 28908 207296 28920
rect 207348 28908 207354 28960
rect 279973 28951 280031 28957
rect 279973 28917 279985 28951
rect 280019 28948 280031 28951
rect 280062 28948 280068 28960
rect 280019 28920 280068 28948
rect 280019 28917 280031 28920
rect 279973 28911 280031 28917
rect 280062 28908 280068 28920
rect 280120 28908 280126 28960
rect 183756 28824 183784 28908
rect 183738 28772 183744 28824
rect 183796 28772 183802 28824
rect 388714 28772 388720 28824
rect 388772 28812 388778 28824
rect 388898 28812 388904 28824
rect 388772 28784 388904 28812
rect 388772 28772 388778 28784
rect 388898 28772 388904 28784
rect 388956 28772 388962 28824
rect 150710 27656 150716 27668
rect 150671 27628 150716 27656
rect 150710 27616 150716 27628
rect 150768 27616 150774 27668
rect 211154 27616 211160 27668
rect 211212 27656 211218 27668
rect 211338 27656 211344 27668
rect 211212 27628 211344 27656
rect 211212 27616 211218 27628
rect 211338 27616 211344 27628
rect 211396 27616 211402 27668
rect 234706 27656 234712 27668
rect 234667 27628 234712 27656
rect 234706 27616 234712 27628
rect 234764 27616 234770 27668
rect 238846 27656 238852 27668
rect 238807 27628 238852 27656
rect 238846 27616 238852 27628
rect 238904 27616 238910 27668
rect 243722 27656 243728 27668
rect 243683 27628 243728 27656
rect 243722 27616 243728 27628
rect 243780 27616 243786 27668
rect 248322 27656 248328 27668
rect 248283 27628 248328 27656
rect 248322 27616 248328 27628
rect 248380 27616 248386 27668
rect 271877 27659 271935 27665
rect 271877 27625 271889 27659
rect 271923 27656 271935 27659
rect 272150 27656 272156 27668
rect 271923 27628 272156 27656
rect 271923 27625 271935 27628
rect 271877 27619 271935 27625
rect 272150 27616 272156 27628
rect 272208 27616 272214 27668
rect 157337 27591 157395 27597
rect 157337 27557 157349 27591
rect 157383 27588 157395 27591
rect 157426 27588 157432 27600
rect 157383 27560 157432 27588
rect 157383 27557 157395 27560
rect 157337 27551 157395 27557
rect 157426 27548 157432 27560
rect 157484 27548 157490 27600
rect 276106 27588 276112 27600
rect 276067 27560 276112 27588
rect 276106 27548 276112 27560
rect 276164 27548 276170 27600
rect 325694 27588 325700 27600
rect 325655 27560 325700 27588
rect 325694 27548 325700 27560
rect 325752 27548 325758 27600
rect 420454 27588 420460 27600
rect 420415 27560 420460 27588
rect 420454 27548 420460 27560
rect 420512 27548 420518 27600
rect 357710 26364 357716 26376
rect 357671 26336 357716 26364
rect 357710 26324 357716 26336
rect 357768 26324 357774 26376
rect 175550 26296 175556 26308
rect 175511 26268 175556 26296
rect 175550 26256 175556 26268
rect 175608 26256 175614 26308
rect 179414 26256 179420 26308
rect 179472 26296 179478 26308
rect 179506 26296 179512 26308
rect 179472 26268 179512 26296
rect 179472 26256 179478 26268
rect 179506 26256 179512 26268
rect 179564 26256 179570 26308
rect 243722 26296 243728 26308
rect 243683 26268 243728 26296
rect 243722 26256 243728 26268
rect 243780 26256 243786 26308
rect 301866 26228 301872 26240
rect 301827 26200 301872 26228
rect 301866 26188 301872 26200
rect 301924 26188 301930 26240
rect 357710 26188 357716 26240
rect 357768 26228 357774 26240
rect 357897 26231 357955 26237
rect 357897 26228 357909 26231
rect 357768 26200 357909 26228
rect 357768 26188 357774 26200
rect 357897 26197 357909 26200
rect 357943 26197 357955 26231
rect 415026 26228 415032 26240
rect 414987 26200 415032 26228
rect 357897 26191 357955 26197
rect 415026 26188 415032 26200
rect 415084 26188 415090 26240
rect 431497 26231 431555 26237
rect 431497 26197 431509 26231
rect 431543 26228 431555 26231
rect 431678 26228 431684 26240
rect 431543 26200 431684 26228
rect 431543 26197 431555 26200
rect 431497 26191 431555 26197
rect 431678 26188 431684 26200
rect 431736 26188 431742 26240
rect 383378 25276 383384 25288
rect 383339 25248 383384 25276
rect 383378 25236 383384 25248
rect 383436 25236 383442 25288
rect 178034 25032 178040 25084
rect 178092 25072 178098 25084
rect 178092 25044 178137 25072
rect 178092 25032 178098 25044
rect 73614 24828 73620 24880
rect 73672 24868 73678 24880
rect 73890 24868 73896 24880
rect 73672 24840 73896 24868
rect 73672 24828 73678 24840
rect 73890 24828 73896 24840
rect 73948 24828 73954 24880
rect 175550 24868 175556 24880
rect 175511 24840 175556 24868
rect 175550 24828 175556 24840
rect 175608 24828 175614 24880
rect 179417 24803 179475 24809
rect 179417 24769 179429 24803
rect 179463 24800 179475 24803
rect 179506 24800 179512 24812
rect 179463 24772 179512 24800
rect 179463 24769 179475 24772
rect 179417 24763 179475 24769
rect 179506 24760 179512 24772
rect 179564 24760 179570 24812
rect 178034 24692 178040 24744
rect 178092 24732 178098 24744
rect 178092 24704 178137 24732
rect 178092 24692 178098 24704
rect 147858 24148 147864 24200
rect 147916 24188 147922 24200
rect 148042 24188 148048 24200
rect 147916 24160 148048 24188
rect 147916 24148 147922 24160
rect 148042 24148 148048 24160
rect 148100 24148 148106 24200
rect 220906 24148 220912 24200
rect 220964 24188 220970 24200
rect 221090 24188 221096 24200
rect 220964 24160 221096 24188
rect 220964 24148 220970 24160
rect 221090 24148 221096 24160
rect 221148 24148 221154 24200
rect 234617 22831 234675 22837
rect 234617 22797 234629 22831
rect 234663 22828 234675 22831
rect 234706 22828 234712 22840
rect 234663 22800 234712 22828
rect 234663 22797 234675 22800
rect 234617 22791 234675 22797
rect 234706 22788 234712 22800
rect 234764 22788 234770 22840
rect 394510 22244 394516 22296
rect 394568 22244 394574 22296
rect 205729 22219 205787 22225
rect 205729 22185 205741 22219
rect 205775 22216 205787 22219
rect 205910 22216 205916 22228
rect 205775 22188 205916 22216
rect 205775 22185 205787 22188
rect 205729 22179 205787 22185
rect 205910 22176 205916 22188
rect 205968 22176 205974 22228
rect 394418 22176 394424 22228
rect 394476 22216 394482 22228
rect 394528 22216 394556 22244
rect 394476 22188 394556 22216
rect 394476 22176 394482 22188
rect 181162 22148 181168 22160
rect 181088 22120 181168 22148
rect 181088 22092 181116 22120
rect 181162 22108 181168 22120
rect 181220 22108 181226 22160
rect 212718 22108 212724 22160
rect 212776 22108 212782 22160
rect 233326 22148 233332 22160
rect 233287 22120 233332 22148
rect 233326 22108 233332 22120
rect 233384 22108 233390 22160
rect 243722 22108 243728 22160
rect 243780 22108 243786 22160
rect 404078 22148 404084 22160
rect 404004 22120 404084 22148
rect 3142 22040 3148 22092
rect 3200 22080 3206 22092
rect 132218 22080 132224 22092
rect 3200 22052 132224 22080
rect 3200 22040 3206 22052
rect 132218 22040 132224 22052
rect 132276 22040 132282 22092
rect 181070 22040 181076 22092
rect 181128 22040 181134 22092
rect 200206 22040 200212 22092
rect 200264 22080 200270 22092
rect 200390 22080 200396 22092
rect 200264 22052 200396 22080
rect 200264 22040 200270 22052
rect 200390 22040 200396 22052
rect 200448 22040 200454 22092
rect 212736 22024 212764 22108
rect 214098 22040 214104 22092
rect 214156 22040 214162 22092
rect 212718 21972 212724 22024
rect 212776 21972 212782 22024
rect 214116 22012 214144 22040
rect 243740 22024 243768 22108
rect 404004 22092 404032 22120
rect 404078 22108 404084 22120
rect 404136 22108 404142 22160
rect 244366 22040 244372 22092
rect 244424 22080 244430 22092
rect 244550 22080 244556 22092
rect 244424 22052 244556 22080
rect 244424 22040 244430 22052
rect 244550 22040 244556 22052
rect 244608 22040 244614 22092
rect 245838 22040 245844 22092
rect 245896 22080 245902 22092
rect 246022 22080 246028 22092
rect 245896 22052 246028 22080
rect 245896 22040 245902 22052
rect 246022 22040 246028 22052
rect 246080 22040 246086 22092
rect 403986 22040 403992 22092
rect 404044 22040 404050 22092
rect 214190 22012 214196 22024
rect 214116 21984 214196 22012
rect 214190 21972 214196 21984
rect 214248 21972 214254 22024
rect 243722 21972 243728 22024
rect 243780 21972 243786 22024
rect 357894 22012 357900 22024
rect 357855 21984 357900 22012
rect 357894 21972 357900 21984
rect 357952 21972 357958 22024
rect 73890 20000 73896 20052
rect 73948 20040 73954 20052
rect 74261 20043 74319 20049
rect 74261 20040 74273 20043
rect 73948 20012 74273 20040
rect 73948 20000 73954 20012
rect 74261 20009 74273 20012
rect 74307 20009 74319 20043
rect 74261 20003 74319 20009
rect 173894 20000 173900 20052
rect 173952 20040 173958 20052
rect 173989 20043 174047 20049
rect 173989 20040 174001 20043
rect 173952 20012 174001 20040
rect 173952 20000 173958 20012
rect 173989 20009 174001 20012
rect 174035 20009 174047 20043
rect 173989 20003 174047 20009
rect 190641 19431 190699 19437
rect 190641 19397 190653 19431
rect 190687 19428 190699 19431
rect 190730 19428 190736 19440
rect 190687 19400 190736 19428
rect 190687 19397 190699 19400
rect 190641 19391 190699 19397
rect 190730 19388 190736 19400
rect 190788 19388 190794 19440
rect 159082 19320 159088 19372
rect 159140 19360 159146 19372
rect 159266 19360 159272 19372
rect 159140 19332 159272 19360
rect 159140 19320 159146 19332
rect 159266 19320 159272 19332
rect 159324 19320 159330 19372
rect 162946 19320 162952 19372
rect 163004 19360 163010 19372
rect 163130 19360 163136 19372
rect 163004 19332 163136 19360
rect 163004 19320 163010 19332
rect 163130 19320 163136 19332
rect 163188 19320 163194 19372
rect 184934 19360 184940 19372
rect 184895 19332 184940 19360
rect 184934 19320 184940 19332
rect 184992 19320 184998 19372
rect 205726 19360 205732 19372
rect 205687 19332 205732 19360
rect 205726 19320 205732 19332
rect 205784 19320 205790 19372
rect 211154 19320 211160 19372
rect 211212 19360 211218 19372
rect 211338 19360 211344 19372
rect 211212 19332 211344 19360
rect 211212 19320 211218 19332
rect 211338 19320 211344 19332
rect 211396 19320 211402 19372
rect 216674 19320 216680 19372
rect 216732 19360 216738 19372
rect 216950 19360 216956 19372
rect 216732 19332 216956 19360
rect 216732 19320 216738 19332
rect 216950 19320 216956 19332
rect 217008 19320 217014 19372
rect 229094 19320 229100 19372
rect 229152 19360 229158 19372
rect 229278 19360 229284 19372
rect 229152 19332 229284 19360
rect 229152 19320 229158 19332
rect 229278 19320 229284 19332
rect 229336 19320 229342 19372
rect 279970 19360 279976 19372
rect 279931 19332 279976 19360
rect 279970 19320 279976 19332
rect 280028 19320 280034 19372
rect 383378 19360 383384 19372
rect 383339 19332 383384 19360
rect 383378 19320 383384 19332
rect 383436 19320 383442 19372
rect 143626 19292 143632 19304
rect 143587 19264 143632 19292
rect 143626 19252 143632 19264
rect 143684 19252 143690 19304
rect 200390 19292 200396 19304
rect 200351 19264 200396 19292
rect 200390 19252 200396 19264
rect 200448 19252 200454 19304
rect 233326 19292 233332 19304
rect 233287 19264 233332 19292
rect 233326 19252 233332 19264
rect 233384 19252 233390 19304
rect 244550 19292 244556 19304
rect 244511 19264 244556 19292
rect 244550 19252 244556 19264
rect 244608 19252 244614 19304
rect 394326 19292 394332 19304
rect 394287 19264 394332 19292
rect 394326 19252 394332 19264
rect 394384 19252 394390 19304
rect 425974 19252 425980 19304
rect 426032 19292 426038 19304
rect 426066 19292 426072 19304
rect 426032 19264 426072 19292
rect 426032 19252 426038 19264
rect 426066 19252 426072 19264
rect 426124 19252 426130 19304
rect 274818 18136 274824 18148
rect 274779 18108 274824 18136
rect 274818 18096 274824 18108
rect 274876 18096 274882 18148
rect 190638 18000 190644 18012
rect 190599 17972 190644 18000
rect 190638 17960 190644 17972
rect 190696 17960 190702 18012
rect 234614 18000 234620 18012
rect 234575 17972 234620 18000
rect 234614 17960 234620 17972
rect 234672 17960 234678 18012
rect 276106 18000 276112 18012
rect 276067 17972 276112 18000
rect 276106 17960 276112 17972
rect 276164 17960 276170 18012
rect 420457 18003 420515 18009
rect 420457 17969 420469 18003
rect 420503 18000 420515 18003
rect 420546 18000 420552 18012
rect 420503 17972 420552 18000
rect 420503 17969 420515 17972
rect 420457 17963 420515 17969
rect 420546 17960 420552 17972
rect 420604 17960 420610 18012
rect 436738 17892 436744 17944
rect 436796 17932 436802 17944
rect 579798 17932 579804 17944
rect 436796 17904 579804 17932
rect 436796 17892 436802 17904
rect 579798 17892 579804 17904
rect 579856 17892 579862 17944
rect 415026 16640 415032 16652
rect 414987 16612 415032 16640
rect 415026 16600 415032 16612
rect 415084 16600 415090 16652
rect 431494 16640 431500 16652
rect 431455 16612 431500 16640
rect 431494 16600 431500 16612
rect 431552 16600 431558 16652
rect 383286 12560 383292 12572
rect 383247 12532 383292 12560
rect 383286 12520 383292 12532
rect 383344 12520 383350 12572
rect 168377 12495 168435 12501
rect 168377 12461 168389 12495
rect 168423 12492 168435 12495
rect 168466 12492 168472 12504
rect 168423 12464 168472 12492
rect 168423 12461 168435 12464
rect 168377 12455 168435 12461
rect 168466 12452 168472 12464
rect 168524 12452 168530 12504
rect 183738 12492 183744 12504
rect 183664 12464 183744 12492
rect 183664 12436 183692 12464
rect 183738 12452 183744 12464
rect 183796 12452 183802 12504
rect 211338 12492 211344 12504
rect 211264 12464 211344 12492
rect 211264 12436 211292 12464
rect 211338 12452 211344 12464
rect 211396 12452 211402 12504
rect 276106 12452 276112 12504
rect 276164 12452 276170 12504
rect 415026 12492 415032 12504
rect 414952 12464 415032 12492
rect 183646 12384 183652 12436
rect 183704 12384 183710 12436
rect 211246 12384 211252 12436
rect 211304 12384 211310 12436
rect 74258 12356 74264 12368
rect 74219 12328 74264 12356
rect 74258 12316 74264 12328
rect 74316 12316 74322 12368
rect 178126 12356 178132 12368
rect 178087 12328 178132 12356
rect 178126 12316 178132 12328
rect 178184 12316 178190 12368
rect 276124 12356 276152 12452
rect 414952 12436 414980 12464
rect 415026 12452 415032 12464
rect 415084 12452 415090 12504
rect 420546 12492 420552 12504
rect 420472 12464 420552 12492
rect 420472 12436 420500 12464
rect 420546 12452 420552 12464
rect 420604 12452 420610 12504
rect 280338 12384 280344 12436
rect 280396 12424 280402 12436
rect 281258 12424 281264 12436
rect 280396 12396 281264 12424
rect 280396 12384 280402 12396
rect 281258 12384 281264 12396
rect 281316 12384 281322 12436
rect 321738 12384 321744 12436
rect 321796 12384 321802 12436
rect 414934 12384 414940 12436
rect 414992 12384 414998 12436
rect 420454 12384 420460 12436
rect 420512 12384 420518 12436
rect 463694 12384 463700 12436
rect 463752 12424 463758 12436
rect 464338 12424 464344 12436
rect 463752 12396 464344 12424
rect 463752 12384 463758 12396
rect 464338 12384 464344 12396
rect 464396 12384 464402 12436
rect 276474 12356 276480 12368
rect 276124 12328 276480 12356
rect 276474 12316 276480 12328
rect 276532 12316 276538 12368
rect 321756 12356 321784 12384
rect 322750 12356 322756 12368
rect 321756 12328 322756 12356
rect 322750 12316 322756 12328
rect 322808 12316 322814 12368
rect 200390 12288 200396 12300
rect 200351 12260 200396 12288
rect 200390 12248 200396 12260
rect 200448 12248 200454 12300
rect 205542 12112 205548 12164
rect 205600 12152 205606 12164
rect 205726 12152 205732 12164
rect 205600 12124 205732 12152
rect 205600 12112 205606 12124
rect 205726 12112 205732 12124
rect 205784 12112 205790 12164
rect 246022 11908 246028 11960
rect 246080 11908 246086 11960
rect 244550 11880 244556 11892
rect 244511 11852 244556 11880
rect 244550 11840 244556 11852
rect 244608 11840 244614 11892
rect 246040 11824 246068 11908
rect 246022 11772 246028 11824
rect 246080 11772 246086 11824
rect 371050 10684 371056 10736
rect 371108 10724 371114 10736
rect 459646 10724 459652 10736
rect 371108 10696 459652 10724
rect 371108 10684 371114 10696
rect 459646 10684 459652 10696
rect 459704 10684 459710 10736
rect 372338 10616 372344 10668
rect 372396 10656 372402 10668
rect 463234 10656 463240 10668
rect 372396 10628 463240 10656
rect 372396 10616 372402 10628
rect 463234 10616 463240 10628
rect 463292 10616 463298 10668
rect 375190 10548 375196 10600
rect 375248 10588 375254 10600
rect 466822 10588 466828 10600
rect 375248 10560 466828 10588
rect 375248 10548 375254 10560
rect 466822 10548 466828 10560
rect 466880 10548 466886 10600
rect 376570 10480 376576 10532
rect 376628 10520 376634 10532
rect 470318 10520 470324 10532
rect 376628 10492 470324 10520
rect 376628 10480 376634 10492
rect 470318 10480 470324 10492
rect 470376 10480 470382 10532
rect 377950 10412 377956 10464
rect 378008 10452 378014 10464
rect 473354 10452 473360 10464
rect 378008 10424 473360 10452
rect 378008 10412 378014 10424
rect 473354 10412 473360 10424
rect 473412 10412 473418 10464
rect 380802 10344 380808 10396
rect 380860 10384 380866 10396
rect 477586 10384 477592 10396
rect 380860 10356 477592 10384
rect 380860 10344 380866 10356
rect 477586 10344 477592 10356
rect 477644 10344 477650 10396
rect 382090 10276 382096 10328
rect 382148 10316 382154 10328
rect 481082 10316 481088 10328
rect 382148 10288 481088 10316
rect 382148 10276 382154 10288
rect 481082 10276 481088 10288
rect 481140 10276 481146 10328
rect 143629 9707 143687 9713
rect 143629 9673 143641 9707
rect 143675 9704 143687 9707
rect 143718 9704 143724 9716
rect 143675 9676 143724 9704
rect 143675 9673 143687 9676
rect 143629 9667 143687 9673
rect 143718 9664 143724 9676
rect 143776 9664 143782 9716
rect 157334 9704 157340 9716
rect 157295 9676 157340 9704
rect 157334 9664 157340 9676
rect 157392 9664 157398 9716
rect 168374 9704 168380 9716
rect 168335 9676 168380 9704
rect 168374 9664 168380 9676
rect 168432 9664 168438 9716
rect 190638 9664 190644 9716
rect 190696 9704 190702 9716
rect 190730 9704 190736 9716
rect 190696 9676 190736 9704
rect 190696 9664 190702 9676
rect 190730 9664 190736 9676
rect 190788 9664 190794 9716
rect 228910 9664 228916 9716
rect 228968 9704 228974 9716
rect 229186 9704 229192 9716
rect 228968 9676 229192 9704
rect 228968 9664 228974 9676
rect 229186 9664 229192 9676
rect 229244 9664 229250 9716
rect 234614 9664 234620 9716
rect 234672 9704 234678 9716
rect 234706 9704 234712 9716
rect 234672 9676 234712 9704
rect 234672 9664 234678 9676
rect 234706 9664 234712 9676
rect 234764 9664 234770 9716
rect 274821 9707 274879 9713
rect 274821 9673 274833 9707
rect 274867 9704 274879 9707
rect 275278 9704 275284 9716
rect 274867 9676 275284 9704
rect 274867 9673 274879 9676
rect 274821 9667 274879 9673
rect 275278 9664 275284 9676
rect 275336 9664 275342 9716
rect 325697 9707 325755 9713
rect 325697 9673 325709 9707
rect 325743 9704 325755 9707
rect 326246 9704 326252 9716
rect 325743 9676 326252 9704
rect 325743 9673 325755 9676
rect 325697 9667 325755 9673
rect 326246 9664 326252 9676
rect 326304 9664 326310 9716
rect 383286 9704 383292 9716
rect 383247 9676 383292 9704
rect 383286 9664 383292 9676
rect 383344 9664 383350 9716
rect 394329 9707 394387 9713
rect 394329 9673 394341 9707
rect 394375 9704 394387 9707
rect 394418 9704 394424 9716
rect 394375 9676 394424 9704
rect 394375 9673 394387 9676
rect 394329 9667 394387 9673
rect 394418 9664 394424 9676
rect 394476 9664 394482 9716
rect 87322 9596 87328 9648
rect 87380 9636 87386 9648
rect 168285 9639 168343 9645
rect 168285 9636 168297 9639
rect 87380 9608 168297 9636
rect 87380 9596 87386 9608
rect 168285 9605 168297 9608
rect 168331 9605 168343 9639
rect 168285 9599 168343 9605
rect 168469 9639 168527 9645
rect 168469 9605 168481 9639
rect 168515 9636 168527 9639
rect 178129 9639 178187 9645
rect 178129 9636 178141 9639
rect 168515 9608 178141 9636
rect 168515 9605 168527 9608
rect 168469 9599 168527 9605
rect 178129 9605 178141 9608
rect 178175 9605 178187 9639
rect 183646 9636 183652 9648
rect 183607 9608 183652 9636
rect 178129 9599 178187 9605
rect 183646 9596 183652 9608
rect 183704 9596 183710 9648
rect 368382 9596 368388 9648
rect 368440 9636 368446 9648
rect 454862 9636 454868 9648
rect 368440 9608 454868 9636
rect 368440 9596 368446 9608
rect 454862 9596 454868 9608
rect 454920 9596 454926 9648
rect 75454 9528 75460 9580
rect 75512 9568 75518 9580
rect 168193 9571 168251 9577
rect 168193 9568 168205 9571
rect 75512 9540 168205 9568
rect 75512 9528 75518 9540
rect 168193 9537 168205 9540
rect 168239 9537 168251 9571
rect 168193 9531 168251 9537
rect 371142 9528 371148 9580
rect 371200 9568 371206 9580
rect 458450 9568 458456 9580
rect 371200 9540 458456 9568
rect 371200 9528 371206 9540
rect 458450 9528 458456 9540
rect 458508 9528 458514 9580
rect 68278 9460 68284 9512
rect 68336 9500 68342 9512
rect 168374 9500 168380 9512
rect 68336 9472 168380 9500
rect 68336 9460 68342 9472
rect 168374 9460 168380 9472
rect 168432 9460 168438 9512
rect 183554 9460 183560 9512
rect 183612 9500 183618 9512
rect 183612 9472 183657 9500
rect 183612 9460 183618 9472
rect 372430 9460 372436 9512
rect 372488 9500 372494 9512
rect 462038 9500 462044 9512
rect 372488 9472 462044 9500
rect 372488 9460 372494 9472
rect 462038 9460 462044 9472
rect 462096 9460 462102 9512
rect 61194 9392 61200 9444
rect 61252 9432 61258 9444
rect 164418 9432 164424 9444
rect 61252 9404 164424 9432
rect 61252 9392 61258 9404
rect 164418 9392 164424 9404
rect 164476 9392 164482 9444
rect 168193 9435 168251 9441
rect 168193 9401 168205 9435
rect 168239 9432 168251 9435
rect 172606 9432 172612 9444
rect 168239 9404 172612 9432
rect 168239 9401 168251 9404
rect 168193 9395 168251 9401
rect 172606 9392 172612 9404
rect 172664 9392 172670 9444
rect 419442 9392 419448 9444
rect 419500 9432 419506 9444
rect 552382 9432 552388 9444
rect 419500 9404 552388 9432
rect 419500 9392 419506 9404
rect 552382 9392 552388 9404
rect 552440 9392 552446 9444
rect 55214 9324 55220 9376
rect 55272 9364 55278 9376
rect 161474 9364 161480 9376
rect 55272 9336 161480 9364
rect 55272 9324 55278 9336
rect 161474 9324 161480 9336
rect 161532 9324 161538 9376
rect 420454 9324 420460 9376
rect 420512 9364 420518 9376
rect 555970 9364 555976 9376
rect 420512 9336 555976 9364
rect 420512 9324 420518 9336
rect 555970 9324 555976 9336
rect 556028 9324 556034 9376
rect 58802 9256 58808 9308
rect 58860 9296 58866 9308
rect 164326 9296 164332 9308
rect 58860 9268 164332 9296
rect 58860 9256 58866 9268
rect 164326 9256 164332 9268
rect 164384 9256 164390 9308
rect 422110 9256 422116 9308
rect 422168 9296 422174 9308
rect 559558 9296 559564 9308
rect 422168 9268 559564 9296
rect 422168 9256 422174 9268
rect 559558 9256 559564 9268
rect 559616 9256 559622 9308
rect 54018 9188 54024 9240
rect 54076 9228 54082 9240
rect 161566 9228 161572 9240
rect 54076 9200 161572 9228
rect 54076 9188 54082 9200
rect 161566 9188 161572 9200
rect 161624 9188 161630 9240
rect 409506 9188 409512 9240
rect 409564 9228 409570 9240
rect 409782 9228 409788 9240
rect 409564 9200 409788 9228
rect 409564 9188 409570 9200
rect 409782 9188 409788 9200
rect 409840 9188 409846 9240
rect 424962 9188 424968 9240
rect 425020 9228 425026 9240
rect 563146 9228 563152 9240
rect 425020 9200 563152 9228
rect 425020 9188 425026 9200
rect 563146 9188 563152 9200
rect 563204 9188 563210 9240
rect 46934 9120 46940 9172
rect 46992 9160 46998 9172
rect 157334 9160 157340 9172
rect 46992 9132 157340 9160
rect 46992 9120 46998 9132
rect 157334 9120 157340 9132
rect 157392 9120 157398 9172
rect 350350 9120 350356 9172
rect 350408 9160 350414 9172
rect 420362 9160 420368 9172
rect 350408 9132 420368 9160
rect 350408 9120 350414 9132
rect 420362 9120 420368 9132
rect 420420 9120 420426 9172
rect 425974 9120 425980 9172
rect 426032 9160 426038 9172
rect 566734 9160 566740 9172
rect 426032 9132 566740 9160
rect 426032 9120 426038 9132
rect 566734 9120 566740 9132
rect 566792 9120 566798 9172
rect 40954 9052 40960 9104
rect 41012 9092 41018 9104
rect 154666 9092 154672 9104
rect 41012 9064 154672 9092
rect 41012 9052 41018 9064
rect 154666 9052 154672 9064
rect 154724 9052 154730 9104
rect 353202 9052 353208 9104
rect 353260 9092 353266 9104
rect 423950 9092 423956 9104
rect 353260 9064 423956 9092
rect 353260 9052 353266 9064
rect 423950 9052 423956 9064
rect 424008 9052 424014 9104
rect 427630 9052 427636 9104
rect 427688 9092 427694 9104
rect 570230 9092 570236 9104
rect 427688 9064 570236 9092
rect 427688 9052 427694 9064
rect 570230 9052 570236 9064
rect 570288 9052 570294 9104
rect 26694 8984 26700 9036
rect 26752 9024 26758 9036
rect 147766 9024 147772 9036
rect 26752 8996 147772 9024
rect 26752 8984 26758 8996
rect 147766 8984 147772 8996
rect 147824 8984 147830 9036
rect 354490 8984 354496 9036
rect 354548 9024 354554 9036
rect 427538 9024 427544 9036
rect 354548 8996 427544 9024
rect 354548 8984 354554 8996
rect 427538 8984 427544 8996
rect 427596 8984 427602 9036
rect 431494 8984 431500 9036
rect 431552 9024 431558 9036
rect 577406 9024 577412 9036
rect 431552 8996 577412 9024
rect 431552 8984 431558 8996
rect 577406 8984 577412 8996
rect 577464 8984 577470 9036
rect 6454 8916 6460 8968
rect 6512 8956 6518 8968
rect 136818 8956 136824 8968
rect 6512 8928 136824 8956
rect 6512 8916 6518 8928
rect 136818 8916 136824 8928
rect 136876 8916 136882 8968
rect 355870 8916 355876 8968
rect 355928 8956 355934 8968
rect 431126 8956 431132 8968
rect 355928 8928 431132 8956
rect 355928 8916 355934 8928
rect 431126 8916 431132 8928
rect 431184 8916 431190 8968
rect 433150 8916 433156 8968
rect 433208 8956 433214 8968
rect 580994 8956 581000 8968
rect 433208 8928 581000 8956
rect 433208 8916 433214 8928
rect 580994 8916 581000 8928
rect 581052 8916 581058 8968
rect 106366 8848 106372 8900
rect 106424 8888 106430 8900
rect 187786 8888 187792 8900
rect 106424 8860 187792 8888
rect 106424 8848 106430 8860
rect 187786 8848 187792 8860
rect 187844 8848 187850 8900
rect 369762 8848 369768 8900
rect 369820 8888 369826 8900
rect 456058 8888 456064 8900
rect 369820 8860 456064 8888
rect 369820 8848 369826 8860
rect 456058 8848 456064 8860
rect 456116 8848 456122 8900
rect 119430 8780 119436 8832
rect 119488 8820 119494 8832
rect 194778 8820 194784 8832
rect 119488 8792 194784 8820
rect 119488 8780 119494 8792
rect 194778 8780 194784 8792
rect 194836 8780 194842 8832
rect 366910 8780 366916 8832
rect 366968 8820 366974 8832
rect 452470 8820 452476 8832
rect 366968 8792 452476 8820
rect 366968 8780 366974 8792
rect 452470 8780 452476 8792
rect 452528 8780 452534 8832
rect 120626 8712 120632 8764
rect 120684 8752 120690 8764
rect 190546 8752 190552 8764
rect 120684 8724 190552 8752
rect 120684 8712 120690 8724
rect 190546 8712 190552 8724
rect 190604 8712 190610 8764
rect 365530 8712 365536 8764
rect 365588 8752 365594 8764
rect 448974 8752 448980 8764
rect 365588 8724 448980 8752
rect 365588 8712 365594 8724
rect 448974 8712 448980 8724
rect 449032 8712 449038 8764
rect 361390 8644 361396 8696
rect 361448 8684 361454 8696
rect 441798 8684 441804 8696
rect 361448 8656 441804 8684
rect 361448 8644 361454 8656
rect 441798 8644 441804 8656
rect 441856 8644 441862 8696
rect 364242 8576 364248 8628
rect 364300 8616 364306 8628
rect 445386 8616 445392 8628
rect 364300 8588 445392 8616
rect 364300 8576 364306 8588
rect 445386 8576 445392 8588
rect 445444 8576 445450 8628
rect 360010 8508 360016 8560
rect 360068 8548 360074 8560
rect 438210 8548 438216 8560
rect 360068 8520 438216 8548
rect 360068 8508 360074 8520
rect 438210 8508 438216 8520
rect 438268 8508 438274 8560
rect 358630 8440 358636 8492
rect 358688 8480 358694 8492
rect 434622 8480 434628 8492
rect 358688 8452 434628 8480
rect 358688 8440 358694 8452
rect 434622 8440 434628 8452
rect 434680 8440 434686 8492
rect 247954 8304 247960 8356
rect 248012 8344 248018 8356
rect 248322 8344 248328 8356
rect 248012 8316 248328 8344
rect 248012 8304 248018 8316
rect 248322 8304 248328 8316
rect 248380 8304 248386 8356
rect 301869 8347 301927 8353
rect 301869 8313 301881 8347
rect 301915 8344 301927 8347
rect 302050 8344 302056 8356
rect 301915 8316 302056 8344
rect 301915 8313 301927 8316
rect 301869 8307 301927 8313
rect 302050 8304 302056 8316
rect 302108 8304 302114 8356
rect 357802 8304 357808 8356
rect 357860 8344 357866 8356
rect 357894 8344 357900 8356
rect 357860 8316 357900 8344
rect 357860 8304 357866 8316
rect 357894 8304 357900 8316
rect 357952 8304 357958 8356
rect 3418 8236 3424 8288
rect 3476 8276 3482 8288
rect 131758 8276 131764 8288
rect 3476 8248 131764 8276
rect 3476 8236 3482 8248
rect 131758 8236 131764 8248
rect 131816 8236 131822 8288
rect 133782 8236 133788 8288
rect 133840 8276 133846 8288
rect 203058 8276 203064 8288
rect 133840 8248 203064 8276
rect 133840 8236 133846 8248
rect 203058 8236 203064 8248
rect 203116 8236 203122 8288
rect 384942 8236 384948 8288
rect 385000 8276 385006 8288
rect 414753 8279 414811 8285
rect 414753 8276 414765 8279
rect 385000 8248 414765 8276
rect 385000 8236 385006 8248
rect 414753 8245 414765 8248
rect 414799 8245 414811 8279
rect 414753 8239 414811 8245
rect 415029 8279 415087 8285
rect 415029 8245 415041 8279
rect 415075 8276 415087 8279
rect 486970 8276 486976 8288
rect 415075 8248 486976 8276
rect 415075 8245 415087 8248
rect 415029 8239 415087 8245
rect 486970 8236 486976 8248
rect 487028 8236 487034 8288
rect 34974 8168 34980 8220
rect 35032 8208 35038 8220
rect 127618 8208 127624 8220
rect 35032 8180 127624 8208
rect 35032 8168 35038 8180
rect 127618 8168 127624 8180
rect 127676 8168 127682 8220
rect 127802 8168 127808 8220
rect 127860 8208 127866 8220
rect 198734 8208 198740 8220
rect 127860 8180 198740 8208
rect 127860 8168 127866 8180
rect 198734 8168 198740 8180
rect 198792 8168 198798 8220
rect 387610 8168 387616 8220
rect 387668 8208 387674 8220
rect 490558 8208 490564 8220
rect 387668 8180 490564 8208
rect 387668 8168 387674 8180
rect 490558 8168 490564 8180
rect 490616 8168 490622 8220
rect 51626 8100 51632 8152
rect 51684 8140 51690 8152
rect 160186 8140 160192 8152
rect 51684 8112 160192 8140
rect 51684 8100 51690 8112
rect 160186 8100 160192 8112
rect 160244 8100 160250 8152
rect 388898 8100 388904 8152
rect 388956 8140 388962 8152
rect 494146 8140 494152 8152
rect 388956 8112 494152 8140
rect 388956 8100 388962 8112
rect 494146 8100 494152 8112
rect 494204 8100 494210 8152
rect 48130 8032 48136 8084
rect 48188 8072 48194 8084
rect 158806 8072 158812 8084
rect 48188 8044 158812 8072
rect 48188 8032 48194 8044
rect 158806 8032 158812 8044
rect 158864 8032 158870 8084
rect 390462 8032 390468 8084
rect 390520 8072 390526 8084
rect 497734 8072 497740 8084
rect 390520 8044 497740 8072
rect 390520 8032 390526 8044
rect 497734 8032 497740 8044
rect 497792 8032 497798 8084
rect 20714 7964 20720 8016
rect 20772 8004 20778 8016
rect 143718 8004 143724 8016
rect 20772 7976 143724 8004
rect 20772 7964 20778 7976
rect 143718 7964 143724 7976
rect 143776 7964 143782 8016
rect 144454 7964 144460 8016
rect 144512 8004 144518 8016
rect 208486 8004 208492 8016
rect 144512 7976 208492 8004
rect 144512 7964 144518 7976
rect 208486 7964 208492 7976
rect 208544 7964 208550 8016
rect 393130 7964 393136 8016
rect 393188 8004 393194 8016
rect 501230 8004 501236 8016
rect 393188 7976 501236 8004
rect 393188 7964 393194 7976
rect 501230 7964 501236 7976
rect 501288 7964 501294 8016
rect 13630 7896 13636 7948
rect 13688 7936 13694 7948
rect 140866 7936 140872 7948
rect 13688 7908 140872 7936
rect 13688 7896 13694 7908
rect 140866 7896 140872 7908
rect 140924 7896 140930 7948
rect 143258 7896 143264 7948
rect 143316 7936 143322 7948
rect 207198 7936 207204 7948
rect 143316 7908 207204 7936
rect 143316 7896 143322 7908
rect 207198 7896 207204 7908
rect 207256 7896 207262 7948
rect 394326 7896 394332 7948
rect 394384 7936 394390 7948
rect 504818 7936 504824 7948
rect 394384 7908 504824 7936
rect 394384 7896 394390 7908
rect 504818 7896 504824 7908
rect 504876 7896 504882 7948
rect 7650 7828 7656 7880
rect 7708 7868 7714 7880
rect 136726 7868 136732 7880
rect 7708 7840 136732 7868
rect 7708 7828 7714 7840
rect 136726 7828 136732 7840
rect 136784 7828 136790 7880
rect 140958 7828 140964 7880
rect 141016 7868 141022 7880
rect 205542 7868 205548 7880
rect 141016 7840 205548 7868
rect 141016 7828 141022 7840
rect 205542 7828 205548 7840
rect 205600 7828 205606 7880
rect 395890 7828 395896 7880
rect 395948 7868 395954 7880
rect 508406 7868 508412 7880
rect 395948 7840 508412 7868
rect 395948 7828 395954 7840
rect 508406 7828 508412 7840
rect 508464 7828 508470 7880
rect 1670 7760 1676 7812
rect 1728 7800 1734 7812
rect 133874 7800 133880 7812
rect 1728 7772 133880 7800
rect 1728 7760 1734 7772
rect 133874 7760 133880 7772
rect 133932 7760 133938 7812
rect 136082 7760 136088 7812
rect 136140 7800 136146 7812
rect 202874 7800 202880 7812
rect 136140 7772 202880 7800
rect 136140 7760 136146 7772
rect 202874 7760 202880 7772
rect 202932 7760 202938 7812
rect 413922 7760 413928 7812
rect 413980 7800 413986 7812
rect 541710 7800 541716 7812
rect 413980 7772 541716 7800
rect 413980 7760 413986 7772
rect 541710 7760 541716 7772
rect 541768 7760 541774 7812
rect 5258 7692 5264 7744
rect 5316 7732 5322 7744
rect 136634 7732 136640 7744
rect 5316 7704 136640 7732
rect 5316 7692 5322 7704
rect 136634 7692 136640 7704
rect 136692 7692 136698 7744
rect 139670 7692 139676 7744
rect 139728 7732 139734 7744
rect 205634 7732 205640 7744
rect 139728 7704 205640 7732
rect 139728 7692 139734 7704
rect 205634 7692 205640 7704
rect 205692 7692 205698 7744
rect 344738 7692 344744 7744
rect 344796 7732 344802 7744
rect 409690 7732 409696 7744
rect 344796 7704 409696 7732
rect 344796 7692 344802 7704
rect 409690 7692 409696 7704
rect 409748 7692 409754 7744
rect 414934 7692 414940 7744
rect 414992 7732 414998 7744
rect 545298 7732 545304 7744
rect 414992 7704 545304 7732
rect 414992 7692 414998 7704
rect 545298 7692 545304 7704
rect 545356 7692 545362 7744
rect 2866 7624 2872 7676
rect 2924 7664 2930 7676
rect 135346 7664 135352 7676
rect 2924 7636 135352 7664
rect 2924 7624 2930 7636
rect 135346 7624 135352 7636
rect 135404 7624 135410 7676
rect 137278 7624 137284 7676
rect 137336 7664 137342 7676
rect 204346 7664 204352 7676
rect 137336 7636 204352 7664
rect 137336 7624 137342 7636
rect 204346 7624 204352 7636
rect 204404 7624 204410 7676
rect 347682 7624 347688 7676
rect 347740 7664 347746 7676
rect 413278 7664 413284 7676
rect 347740 7636 413284 7664
rect 347740 7624 347746 7636
rect 413278 7624 413284 7636
rect 413336 7624 413342 7676
rect 416590 7624 416596 7676
rect 416648 7664 416654 7676
rect 548886 7664 548892 7676
rect 416648 7636 548892 7664
rect 416648 7624 416654 7636
rect 548886 7624 548892 7636
rect 548944 7624 548950 7676
rect 566 7556 572 7608
rect 624 7596 630 7608
rect 134150 7596 134156 7608
rect 624 7568 134156 7596
rect 624 7556 630 7568
rect 134150 7556 134156 7568
rect 134208 7556 134214 7608
rect 134886 7556 134892 7608
rect 134944 7596 134950 7608
rect 202966 7596 202972 7608
rect 134944 7568 202972 7596
rect 134944 7556 134950 7568
rect 202966 7556 202972 7568
rect 203024 7556 203030 7608
rect 348970 7556 348976 7608
rect 349028 7596 349034 7608
rect 412637 7599 412695 7605
rect 412637 7596 412649 7599
rect 349028 7568 412649 7596
rect 349028 7556 349034 7568
rect 412637 7565 412649 7568
rect 412683 7565 412695 7599
rect 412637 7559 412695 7565
rect 416774 7556 416780 7608
rect 416832 7596 416838 7608
rect 417970 7596 417976 7608
rect 416832 7568 417976 7596
rect 416832 7556 416838 7568
rect 417970 7556 417976 7568
rect 418028 7556 418034 7608
rect 430482 7556 430488 7608
rect 430540 7596 430546 7608
rect 573818 7596 573824 7608
rect 430540 7568 573824 7596
rect 430540 7556 430546 7568
rect 573818 7556 573824 7568
rect 573876 7556 573882 7608
rect 115934 7488 115940 7540
rect 115992 7528 115998 7540
rect 117130 7528 117136 7540
rect 115992 7500 117136 7528
rect 115992 7488 115998 7500
rect 117130 7488 117136 7500
rect 117188 7488 117194 7540
rect 118234 7488 118240 7540
rect 118292 7528 118298 7540
rect 194594 7528 194600 7540
rect 118292 7500 194600 7528
rect 118292 7488 118298 7500
rect 194594 7488 194600 7500
rect 194652 7488 194658 7540
rect 383286 7488 383292 7540
rect 383344 7528 383350 7540
rect 383344 7500 477448 7528
rect 383344 7488 383350 7500
rect 121822 7420 121828 7472
rect 121880 7460 121886 7472
rect 196066 7460 196072 7472
rect 121880 7432 196072 7460
rect 121880 7420 121886 7432
rect 196066 7420 196072 7432
rect 196124 7420 196130 7472
rect 367002 7420 367008 7472
rect 367060 7460 367066 7472
rect 451274 7460 451280 7472
rect 367060 7432 451280 7460
rect 367060 7420 367066 7432
rect 451274 7420 451280 7432
rect 451332 7420 451338 7472
rect 477420 7460 477448 7500
rect 477494 7488 477500 7540
rect 477552 7528 477558 7540
rect 478690 7528 478696 7540
rect 477552 7500 478696 7528
rect 477552 7488 477558 7500
rect 478690 7488 478696 7500
rect 478748 7488 478754 7540
rect 483474 7460 483480 7472
rect 477420 7432 483480 7460
rect 483474 7420 483480 7432
rect 483532 7420 483538 7472
rect 126606 7352 126612 7404
rect 126664 7392 126670 7404
rect 198826 7392 198832 7404
rect 126664 7364 198832 7392
rect 126664 7352 126670 7364
rect 198826 7352 198832 7364
rect 198884 7352 198890 7404
rect 365622 7352 365628 7404
rect 365680 7392 365686 7404
rect 447778 7392 447784 7404
rect 365680 7364 447784 7392
rect 365680 7352 365686 7364
rect 447778 7352 447784 7364
rect 447836 7352 447842 7404
rect 77846 7284 77852 7336
rect 77904 7324 77910 7336
rect 77904 7296 126008 7324
rect 77904 7284 77910 7296
rect 84930 7216 84936 7268
rect 84988 7256 84994 7268
rect 125980 7256 126008 7296
rect 128998 7284 129004 7336
rect 129056 7324 129062 7336
rect 200114 7324 200120 7336
rect 129056 7296 200120 7324
rect 129056 7284 129062 7296
rect 200114 7284 200120 7296
rect 200172 7284 200178 7336
rect 362862 7284 362868 7336
rect 362920 7324 362926 7336
rect 444190 7324 444196 7336
rect 362920 7296 444196 7324
rect 362920 7284 362926 7296
rect 444190 7284 444196 7296
rect 444248 7284 444254 7336
rect 129090 7256 129096 7268
rect 84988 7228 125916 7256
rect 125980 7228 129096 7256
rect 84988 7216 84994 7228
rect 95694 7148 95700 7200
rect 95752 7188 95758 7200
rect 125781 7191 125839 7197
rect 125781 7188 125793 7191
rect 95752 7160 125793 7188
rect 95752 7148 95758 7160
rect 125781 7157 125793 7160
rect 125827 7157 125839 7191
rect 125888 7188 125916 7228
rect 129090 7216 129096 7228
rect 129148 7216 129154 7268
rect 130194 7216 130200 7268
rect 130252 7256 130258 7268
rect 200390 7256 200396 7268
rect 130252 7228 200396 7256
rect 130252 7216 130258 7228
rect 200390 7216 200396 7228
rect 200448 7216 200454 7268
rect 361482 7216 361488 7268
rect 361540 7256 361546 7268
rect 440602 7256 440608 7268
rect 361540 7228 440608 7256
rect 361540 7216 361546 7228
rect 440602 7216 440608 7228
rect 440660 7216 440666 7268
rect 129182 7188 129188 7200
rect 125888 7160 129188 7188
rect 125781 7151 125839 7157
rect 129182 7148 129188 7160
rect 129240 7148 129246 7200
rect 131390 7148 131396 7200
rect 131448 7188 131454 7200
rect 201586 7188 201592 7200
rect 131448 7160 201592 7188
rect 131448 7148 131454 7160
rect 201586 7148 201592 7160
rect 201644 7148 201650 7200
rect 358722 7148 358728 7200
rect 358780 7188 358786 7200
rect 435818 7188 435824 7200
rect 358780 7160 435824 7188
rect 358780 7148 358786 7160
rect 435818 7148 435824 7160
rect 435876 7148 435882 7200
rect 109954 7080 109960 7132
rect 110012 7120 110018 7132
rect 133046 7120 133052 7132
rect 110012 7092 133052 7120
rect 110012 7080 110018 7092
rect 133046 7080 133052 7092
rect 133104 7080 133110 7132
rect 133138 7080 133144 7132
rect 133196 7120 133202 7132
rect 201494 7120 201500 7132
rect 133196 7092 201500 7120
rect 133196 7080 133202 7092
rect 201494 7080 201500 7092
rect 201552 7080 201558 7132
rect 360102 7080 360108 7132
rect 360160 7120 360166 7132
rect 437014 7120 437020 7132
rect 360160 7092 437020 7120
rect 360160 7080 360166 7092
rect 437014 7080 437020 7092
rect 437072 7080 437078 7132
rect 125781 7055 125839 7061
rect 125781 7021 125793 7055
rect 125827 7052 125839 7055
rect 129274 7052 129280 7064
rect 125827 7024 129280 7052
rect 125827 7021 125839 7024
rect 125781 7015 125839 7021
rect 129274 7012 129280 7024
rect 129332 7012 129338 7064
rect 412637 7055 412695 7061
rect 412637 7021 412649 7055
rect 412683 7052 412695 7055
rect 416866 7052 416872 7064
rect 412683 7024 416872 7052
rect 412683 7021 412695 7024
rect 412637 7015 412695 7021
rect 416866 7012 416872 7024
rect 416924 7012 416930 7064
rect 173986 6916 173992 6928
rect 173947 6888 173992 6916
rect 173986 6876 173992 6888
rect 174044 6876 174050 6928
rect 179414 6916 179420 6928
rect 179375 6888 179420 6916
rect 179414 6876 179420 6888
rect 179472 6876 179478 6928
rect 96890 6808 96896 6860
rect 96948 6848 96954 6860
rect 183557 6851 183615 6857
rect 183557 6848 183569 6851
rect 96948 6820 183569 6848
rect 96948 6808 96954 6820
rect 183557 6817 183569 6820
rect 183603 6817 183615 6851
rect 183557 6811 183615 6817
rect 317138 6808 317144 6860
rect 317196 6848 317202 6860
rect 356146 6848 356152 6860
rect 317196 6820 356152 6848
rect 317196 6808 317202 6820
rect 356146 6808 356152 6820
rect 356204 6808 356210 6860
rect 391750 6808 391756 6860
rect 391808 6848 391814 6860
rect 498930 6848 498936 6860
rect 391808 6820 498936 6848
rect 391808 6808 391814 6820
rect 498930 6808 498936 6820
rect 498988 6808 498994 6860
rect 94498 6740 94504 6792
rect 94556 6780 94562 6792
rect 182266 6780 182272 6792
rect 94556 6752 182272 6780
rect 94556 6740 94562 6752
rect 182266 6740 182272 6752
rect 182324 6740 182330 6792
rect 326890 6740 326896 6792
rect 326948 6780 326954 6792
rect 373994 6780 374000 6792
rect 326948 6752 374000 6780
rect 326948 6740 326954 6752
rect 373994 6740 374000 6752
rect 374052 6740 374058 6792
rect 393222 6740 393228 6792
rect 393280 6780 393286 6792
rect 502426 6780 502432 6792
rect 393280 6752 502432 6780
rect 393280 6740 393286 6752
rect 502426 6740 502432 6752
rect 502484 6740 502490 6792
rect 89714 6672 89720 6724
rect 89772 6712 89778 6724
rect 179414 6712 179420 6724
rect 89772 6684 179420 6712
rect 89772 6672 89778 6684
rect 179414 6672 179420 6684
rect 179472 6672 179478 6724
rect 328178 6672 328184 6724
rect 328236 6712 328242 6724
rect 377582 6712 377588 6724
rect 328236 6684 377588 6712
rect 328236 6672 328242 6684
rect 377582 6672 377588 6684
rect 377640 6672 377646 6724
rect 394602 6672 394608 6724
rect 394660 6712 394666 6724
rect 506014 6712 506020 6724
rect 394660 6684 506020 6712
rect 394660 6672 394666 6684
rect 506014 6672 506020 6684
rect 506072 6672 506078 6724
rect 90910 6604 90916 6656
rect 90968 6644 90974 6656
rect 180886 6644 180892 6656
rect 90968 6616 180892 6644
rect 90968 6604 90974 6616
rect 180886 6604 180892 6616
rect 180944 6604 180950 6656
rect 331030 6604 331036 6656
rect 331088 6644 331094 6656
rect 381170 6644 381176 6656
rect 331088 6616 381176 6644
rect 331088 6604 331094 6616
rect 381170 6604 381176 6616
rect 381228 6604 381234 6656
rect 397362 6604 397368 6656
rect 397420 6644 397426 6656
rect 509602 6644 509608 6656
rect 397420 6616 509608 6644
rect 397420 6604 397426 6616
rect 509602 6604 509608 6616
rect 509660 6604 509666 6656
rect 86126 6536 86132 6588
rect 86184 6576 86190 6588
rect 178034 6576 178040 6588
rect 86184 6548 178040 6576
rect 86184 6536 86190 6548
rect 178034 6536 178040 6548
rect 178092 6536 178098 6588
rect 332410 6536 332416 6588
rect 332468 6576 332474 6588
rect 384666 6576 384672 6588
rect 332468 6548 384672 6576
rect 332468 6536 332474 6548
rect 384666 6536 384672 6548
rect 384724 6536 384730 6588
rect 398650 6536 398656 6588
rect 398708 6576 398714 6588
rect 513190 6576 513196 6588
rect 398708 6548 513196 6576
rect 398708 6536 398714 6548
rect 513190 6536 513196 6548
rect 513248 6536 513254 6588
rect 79042 6468 79048 6520
rect 79100 6508 79106 6520
rect 173986 6508 173992 6520
rect 79100 6480 173992 6508
rect 79100 6468 79106 6480
rect 173986 6468 173992 6480
rect 174044 6468 174050 6520
rect 336642 6468 336648 6520
rect 336700 6508 336706 6520
rect 391842 6508 391848 6520
rect 336700 6480 391848 6508
rect 336700 6468 336706 6480
rect 391842 6468 391848 6480
rect 391900 6468 391906 6520
rect 399938 6468 399944 6520
rect 399996 6508 400002 6520
rect 516778 6508 516784 6520
rect 399996 6480 516784 6508
rect 399996 6468 400002 6480
rect 516778 6468 516784 6480
rect 516836 6468 516842 6520
rect 71866 6400 71872 6452
rect 71924 6440 71930 6452
rect 169846 6440 169852 6452
rect 71924 6412 169852 6440
rect 71924 6400 71930 6412
rect 169846 6400 169852 6412
rect 169904 6400 169910 6452
rect 333698 6400 333704 6452
rect 333756 6440 333762 6452
rect 388254 6440 388260 6452
rect 333756 6412 388260 6440
rect 333756 6400 333762 6412
rect 388254 6400 388260 6412
rect 388312 6400 388318 6452
rect 402790 6400 402796 6452
rect 402848 6440 402854 6452
rect 520274 6440 520280 6452
rect 402848 6412 520280 6440
rect 402848 6400 402854 6412
rect 520274 6400 520280 6412
rect 520332 6400 520338 6452
rect 64782 6332 64788 6384
rect 64840 6372 64846 6384
rect 167086 6372 167092 6384
rect 64840 6344 167092 6372
rect 64840 6332 64846 6344
rect 167086 6332 167092 6344
rect 167144 6332 167150 6384
rect 337930 6332 337936 6384
rect 337988 6372 337994 6384
rect 395430 6372 395436 6384
rect 337988 6344 395436 6372
rect 337988 6332 337994 6344
rect 395430 6332 395436 6344
rect 395488 6332 395494 6384
rect 404170 6332 404176 6384
rect 404228 6372 404234 6384
rect 523862 6372 523868 6384
rect 404228 6344 523868 6372
rect 404228 6332 404234 6344
rect 523862 6332 523868 6344
rect 523920 6332 523926 6384
rect 57606 6264 57612 6316
rect 57664 6304 57670 6316
rect 162854 6304 162860 6316
rect 57664 6276 162860 6304
rect 57664 6264 57670 6276
rect 162854 6264 162860 6276
rect 162912 6264 162918 6316
rect 177482 6264 177488 6316
rect 177540 6304 177546 6316
rect 214190 6304 214196 6316
rect 177540 6276 214196 6304
rect 177540 6264 177546 6276
rect 214190 6264 214196 6276
rect 214248 6264 214254 6316
rect 342162 6264 342168 6316
rect 342220 6304 342226 6316
rect 402514 6304 402520 6316
rect 342220 6276 402520 6304
rect 342220 6264 342226 6276
rect 402514 6264 402520 6276
rect 402572 6264 402578 6316
rect 408402 6264 408408 6316
rect 408460 6304 408466 6316
rect 531038 6304 531044 6316
rect 408460 6276 531044 6304
rect 408460 6264 408466 6276
rect 531038 6264 531044 6276
rect 531096 6264 531102 6316
rect 36170 6196 36176 6248
rect 36228 6236 36234 6248
rect 151814 6236 151820 6248
rect 36228 6208 151820 6236
rect 36228 6196 36234 6208
rect 151814 6196 151820 6208
rect 151872 6196 151878 6248
rect 183554 6196 183560 6248
rect 183612 6236 183618 6248
rect 222286 6236 222292 6248
rect 183612 6208 222292 6236
rect 183612 6196 183618 6208
rect 222286 6196 222292 6208
rect 222344 6196 222350 6248
rect 339310 6196 339316 6248
rect 339368 6236 339374 6248
rect 399018 6236 399024 6248
rect 339368 6208 399024 6236
rect 339368 6196 339374 6208
rect 399018 6196 399024 6208
rect 399076 6196 399082 6248
rect 405550 6196 405556 6248
rect 405608 6236 405614 6248
rect 527450 6236 527456 6248
rect 405608 6208 527456 6236
rect 405608 6196 405614 6208
rect 527450 6196 527456 6208
rect 527508 6196 527514 6248
rect 29086 6128 29092 6180
rect 29144 6168 29150 6180
rect 148042 6168 148048 6180
rect 29144 6140 148048 6168
rect 29144 6128 29150 6140
rect 148042 6128 148048 6140
rect 148100 6128 148106 6180
rect 153930 6128 153936 6180
rect 153988 6168 153994 6180
rect 212718 6168 212724 6180
rect 153988 6140 212724 6168
rect 153988 6128 153994 6140
rect 212718 6128 212724 6140
rect 212776 6128 212782 6180
rect 343450 6128 343456 6180
rect 343508 6168 343514 6180
rect 406102 6168 406108 6180
rect 343508 6140 406108 6168
rect 343508 6128 343514 6140
rect 406102 6128 406108 6140
rect 406160 6128 406166 6180
rect 409598 6128 409604 6180
rect 409656 6168 409662 6180
rect 534534 6168 534540 6180
rect 409656 6140 534540 6168
rect 409656 6128 409662 6140
rect 534534 6128 534540 6140
rect 534592 6128 534598 6180
rect 98086 6060 98092 6112
rect 98144 6100 98150 6112
rect 183649 6103 183707 6109
rect 183649 6100 183661 6103
rect 98144 6072 183661 6100
rect 98144 6060 98150 6072
rect 183649 6069 183661 6072
rect 183695 6069 183707 6103
rect 183649 6063 183707 6069
rect 318702 6060 318708 6112
rect 318760 6100 318766 6112
rect 358538 6100 358544 6112
rect 318760 6072 358544 6100
rect 318760 6060 318766 6072
rect 358538 6060 358544 6072
rect 358596 6060 358602 6112
rect 388990 6060 388996 6112
rect 389048 6100 389054 6112
rect 495342 6100 495348 6112
rect 389048 6072 495348 6100
rect 389048 6060 389054 6072
rect 495342 6060 495348 6072
rect 495400 6060 495406 6112
rect 101582 5992 101588 6044
rect 101640 6032 101646 6044
rect 186314 6032 186320 6044
rect 101640 6004 186320 6032
rect 101640 5992 101646 6004
rect 186314 5992 186320 6004
rect 186372 5992 186378 6044
rect 317230 5992 317236 6044
rect 317288 6032 317294 6044
rect 354950 6032 354956 6044
rect 317288 6004 354956 6032
rect 317288 5992 317294 6004
rect 354950 5992 354956 6004
rect 355008 5992 355014 6044
rect 387702 5992 387708 6044
rect 387760 6032 387766 6044
rect 491754 6032 491760 6044
rect 387760 6004 491760 6032
rect 387760 5992 387766 6004
rect 491754 5992 491760 6004
rect 491812 5992 491818 6044
rect 103974 5924 103980 5976
rect 104032 5964 104038 5976
rect 186498 5964 186504 5976
rect 104032 5936 186504 5964
rect 104032 5924 104038 5936
rect 186498 5924 186504 5936
rect 186556 5924 186562 5976
rect 315942 5924 315948 5976
rect 316000 5964 316006 5976
rect 352558 5964 352564 5976
rect 316000 5936 352564 5964
rect 316000 5924 316006 5936
rect 352558 5924 352564 5936
rect 352616 5924 352622 5976
rect 383470 5924 383476 5976
rect 383528 5964 383534 5976
rect 484578 5964 484584 5976
rect 383528 5936 484584 5964
rect 383528 5924 383534 5936
rect 484578 5924 484584 5936
rect 484636 5924 484642 5976
rect 105170 5856 105176 5908
rect 105228 5896 105234 5908
rect 187694 5896 187700 5908
rect 105228 5868 187700 5896
rect 105228 5856 105234 5868
rect 187694 5856 187700 5868
rect 187752 5856 187758 5908
rect 315850 5856 315856 5908
rect 315908 5896 315914 5908
rect 351362 5896 351368 5908
rect 315908 5868 351368 5896
rect 315908 5856 315914 5868
rect 351362 5856 351368 5868
rect 351420 5856 351426 5908
rect 386322 5856 386328 5908
rect 386380 5896 386386 5908
rect 488166 5896 488172 5908
rect 386380 5868 488172 5896
rect 386380 5856 386386 5868
rect 488166 5856 488172 5868
rect 488224 5856 488230 5908
rect 56410 5788 56416 5840
rect 56468 5828 56474 5840
rect 108298 5828 108304 5840
rect 56468 5800 108304 5828
rect 56468 5788 56474 5800
rect 108298 5788 108304 5800
rect 108356 5788 108362 5840
rect 108758 5788 108764 5840
rect 108816 5828 108822 5840
rect 189166 5828 189172 5840
rect 108816 5800 189172 5828
rect 108816 5788 108822 5800
rect 189166 5788 189172 5800
rect 189224 5788 189230 5840
rect 379330 5788 379336 5840
rect 379388 5828 379394 5840
rect 476298 5828 476304 5840
rect 379388 5800 476304 5828
rect 379388 5788 379394 5800
rect 476298 5788 476304 5800
rect 476356 5788 476362 5840
rect 112346 5720 112352 5772
rect 112404 5760 112410 5772
rect 191926 5760 191932 5772
rect 112404 5732 191932 5760
rect 112404 5720 112410 5732
rect 191926 5720 191932 5732
rect 191984 5720 191990 5772
rect 382182 5720 382188 5772
rect 382240 5760 382246 5772
rect 479886 5760 479892 5772
rect 382240 5732 479892 5760
rect 382240 5720 382246 5732
rect 479886 5720 479892 5732
rect 479944 5720 479950 5772
rect 111150 5652 111156 5704
rect 111208 5692 111214 5704
rect 190546 5692 190552 5704
rect 111208 5664 190552 5692
rect 111208 5652 111214 5664
rect 190546 5652 190552 5664
rect 190604 5652 190610 5704
rect 378042 5652 378048 5704
rect 378100 5692 378106 5704
rect 472710 5692 472716 5704
rect 378100 5664 472716 5692
rect 378100 5652 378106 5664
rect 472710 5652 472716 5664
rect 472768 5652 472774 5704
rect 115934 5584 115940 5636
rect 115992 5624 115998 5636
rect 193214 5624 193220 5636
rect 115992 5596 193220 5624
rect 115992 5584 115998 5596
rect 193214 5584 193220 5596
rect 193272 5584 193278 5636
rect 373902 5584 373908 5636
rect 373960 5624 373966 5636
rect 465626 5624 465632 5636
rect 373960 5596 465632 5624
rect 373960 5584 373966 5596
rect 465626 5584 465632 5596
rect 465684 5584 465690 5636
rect 123018 5516 123024 5568
rect 123076 5556 123082 5568
rect 197446 5556 197452 5568
rect 123076 5528 197452 5556
rect 123076 5516 123082 5528
rect 197446 5516 197452 5528
rect 197504 5516 197510 5568
rect 376662 5516 376668 5568
rect 376720 5556 376726 5568
rect 469122 5556 469128 5568
rect 376720 5528 469128 5556
rect 376720 5516 376726 5528
rect 469122 5516 469128 5528
rect 469180 5516 469186 5568
rect 69474 5448 69480 5500
rect 69532 5488 69538 5500
rect 169938 5488 169944 5500
rect 69532 5460 169944 5488
rect 69532 5448 69538 5460
rect 169938 5448 169944 5460
rect 169996 5448 170002 5500
rect 174170 5448 174176 5500
rect 174228 5488 174234 5500
rect 223666 5488 223672 5500
rect 174228 5460 223672 5488
rect 174228 5448 174234 5460
rect 223666 5448 223672 5460
rect 223724 5448 223730 5500
rect 335170 5448 335176 5500
rect 335228 5488 335234 5500
rect 390646 5488 390652 5500
rect 335228 5460 390652 5488
rect 335228 5448 335234 5460
rect 390646 5448 390652 5460
rect 390704 5448 390710 5500
rect 415302 5448 415308 5500
rect 415360 5488 415366 5500
rect 544102 5488 544108 5500
rect 415360 5460 544108 5488
rect 415360 5448 415366 5460
rect 544102 5448 544108 5460
rect 544160 5448 544166 5500
rect 65978 5380 65984 5432
rect 66036 5420 66042 5432
rect 166994 5420 167000 5432
rect 66036 5392 167000 5420
rect 66036 5380 66042 5392
rect 166994 5380 167000 5392
rect 167052 5380 167058 5432
rect 170582 5380 170588 5432
rect 170640 5420 170646 5432
rect 221090 5420 221096 5432
rect 170640 5392 221096 5420
rect 170640 5380 170646 5392
rect 221090 5380 221096 5392
rect 221148 5380 221154 5432
rect 339402 5380 339408 5432
rect 339460 5420 339466 5432
rect 397822 5420 397828 5432
rect 339460 5392 397828 5420
rect 339460 5380 339466 5392
rect 397822 5380 397828 5392
rect 397880 5380 397886 5432
rect 416682 5380 416688 5432
rect 416740 5420 416746 5432
rect 547690 5420 547696 5432
rect 416740 5392 547696 5420
rect 416740 5380 416746 5392
rect 547690 5380 547696 5392
rect 547748 5380 547754 5432
rect 62390 5312 62396 5364
rect 62448 5352 62454 5364
rect 165706 5352 165712 5364
rect 62448 5324 165712 5352
rect 62448 5312 62454 5324
rect 165706 5312 165712 5324
rect 165764 5312 165770 5364
rect 167086 5312 167092 5364
rect 167144 5352 167150 5364
rect 219526 5352 219532 5364
rect 167144 5324 219532 5352
rect 167144 5312 167150 5324
rect 219526 5312 219532 5324
rect 219584 5312 219590 5364
rect 340690 5312 340696 5364
rect 340748 5352 340754 5364
rect 401318 5352 401324 5364
rect 340748 5324 401324 5352
rect 340748 5312 340754 5324
rect 401318 5312 401324 5324
rect 401376 5312 401382 5364
rect 418062 5312 418068 5364
rect 418120 5352 418126 5364
rect 551186 5352 551192 5364
rect 418120 5324 551192 5352
rect 418120 5312 418126 5324
rect 551186 5312 551192 5324
rect 551244 5312 551250 5364
rect 44542 5244 44548 5296
rect 44600 5284 44606 5296
rect 156230 5284 156236 5296
rect 44600 5256 156236 5284
rect 44600 5244 44606 5256
rect 156230 5244 156236 5256
rect 156288 5244 156294 5296
rect 158714 5244 158720 5296
rect 158772 5284 158778 5296
rect 215386 5284 215392 5296
rect 158772 5256 215392 5284
rect 158772 5244 158778 5256
rect 215386 5244 215392 5256
rect 215444 5244 215450 5296
rect 343542 5244 343548 5296
rect 343600 5284 343606 5296
rect 404906 5284 404912 5296
rect 343600 5256 404912 5284
rect 343600 5244 343606 5256
rect 404906 5244 404912 5256
rect 404964 5244 404970 5296
rect 420822 5244 420828 5296
rect 420880 5284 420886 5296
rect 554774 5284 554780 5296
rect 420880 5256 554780 5284
rect 420880 5244 420886 5256
rect 554774 5244 554780 5256
rect 554832 5244 554838 5296
rect 37366 5176 37372 5228
rect 37424 5216 37430 5228
rect 153286 5216 153292 5228
rect 37424 5188 153292 5216
rect 37424 5176 37430 5188
rect 153286 5176 153292 5188
rect 153344 5176 153350 5228
rect 156322 5176 156328 5228
rect 156380 5216 156386 5228
rect 213914 5216 213920 5228
rect 156380 5188 213920 5216
rect 156380 5176 156386 5188
rect 213914 5176 213920 5188
rect 213972 5176 213978 5228
rect 344830 5176 344836 5228
rect 344888 5216 344894 5228
rect 408678 5216 408684 5228
rect 344888 5188 408684 5216
rect 344888 5176 344894 5188
rect 408678 5176 408684 5188
rect 408736 5176 408742 5228
rect 422202 5176 422208 5228
rect 422260 5216 422266 5228
rect 558362 5216 558368 5228
rect 422260 5188 558368 5216
rect 422260 5176 422266 5188
rect 558362 5176 558368 5188
rect 558420 5176 558426 5228
rect 33870 5108 33876 5160
rect 33928 5148 33934 5160
rect 150710 5148 150716 5160
rect 33928 5120 150716 5148
rect 33928 5108 33934 5120
rect 150710 5108 150716 5120
rect 150768 5108 150774 5160
rect 155126 5108 155132 5160
rect 155184 5148 155190 5160
rect 214006 5148 214012 5160
rect 155184 5120 214012 5148
rect 155184 5108 155190 5120
rect 214006 5108 214012 5120
rect 214064 5108 214070 5160
rect 346302 5108 346308 5160
rect 346360 5148 346366 5160
rect 412082 5148 412088 5160
rect 346360 5120 412088 5148
rect 346360 5108 346366 5120
rect 412082 5108 412088 5120
rect 412140 5108 412146 5160
rect 423582 5108 423588 5160
rect 423640 5148 423646 5160
rect 561950 5148 561956 5160
rect 423640 5120 561956 5148
rect 423640 5108 423646 5120
rect 561950 5108 561956 5120
rect 562008 5108 562014 5160
rect 18322 5040 18328 5092
rect 18380 5080 18386 5092
rect 135438 5080 135444 5092
rect 18380 5052 135444 5080
rect 18380 5040 18386 5052
rect 135438 5040 135444 5052
rect 135496 5040 135502 5092
rect 138474 5040 138480 5092
rect 138532 5080 138538 5092
rect 204254 5080 204260 5092
rect 138532 5052 204260 5080
rect 138532 5040 138538 5052
rect 204254 5040 204260 5052
rect 204312 5040 204318 5092
rect 204346 5040 204352 5092
rect 204404 5080 204410 5092
rect 237466 5080 237472 5092
rect 204404 5052 237472 5080
rect 204404 5040 204410 5052
rect 237466 5040 237472 5052
rect 237524 5040 237530 5092
rect 349062 5040 349068 5092
rect 349120 5080 349126 5092
rect 415670 5080 415676 5092
rect 349120 5052 415676 5080
rect 349120 5040 349126 5052
rect 415670 5040 415676 5052
rect 415728 5040 415734 5092
rect 426342 5040 426348 5092
rect 426400 5080 426406 5092
rect 565538 5080 565544 5092
rect 426400 5052 565544 5080
rect 426400 5040 426406 5052
rect 565538 5040 565544 5052
rect 565596 5040 565602 5092
rect 21910 4972 21916 5024
rect 21968 5012 21974 5024
rect 145098 5012 145104 5024
rect 21968 4984 145104 5012
rect 21968 4972 21974 4984
rect 145098 4972 145104 4984
rect 145156 4972 145162 5024
rect 152734 4972 152740 5024
rect 152792 5012 152798 5024
rect 212534 5012 212540 5024
rect 152792 4984 212540 5012
rect 152792 4972 152798 4984
rect 212534 4972 212540 4984
rect 212592 4972 212598 5024
rect 350442 4972 350448 5024
rect 350500 5012 350506 5024
rect 419166 5012 419172 5024
rect 350500 4984 419172 5012
rect 350500 4972 350506 4984
rect 419166 4972 419172 4984
rect 419224 4972 419230 5024
rect 427722 4972 427728 5024
rect 427780 5012 427786 5024
rect 569034 5012 569040 5024
rect 427780 4984 569040 5012
rect 427780 4972 427786 4984
rect 569034 4972 569040 4984
rect 569092 4972 569098 5024
rect 17218 4904 17224 4956
rect 17276 4944 17282 4956
rect 142246 4944 142252 4956
rect 17276 4916 142252 4944
rect 17276 4904 17282 4916
rect 142246 4904 142252 4916
rect 142304 4904 142310 4956
rect 149238 4904 149244 4956
rect 149296 4944 149302 4956
rect 209866 4944 209872 4956
rect 149296 4916 209872 4944
rect 149296 4904 149302 4916
rect 209866 4904 209872 4916
rect 209924 4904 209930 4956
rect 215846 4904 215852 4956
rect 215904 4944 215910 4956
rect 244550 4944 244556 4956
rect 215904 4916 244556 4944
rect 215904 4904 215910 4916
rect 244550 4904 244556 4916
rect 244608 4904 244614 4956
rect 310422 4904 310428 4956
rect 310480 4944 310486 4956
rect 341886 4944 341892 4956
rect 310480 4916 341892 4944
rect 310480 4904 310486 4916
rect 341886 4904 341892 4916
rect 341944 4904 341950 4956
rect 354582 4904 354588 4956
rect 354640 4944 354646 4956
rect 426342 4944 426348 4956
rect 354640 4916 426348 4944
rect 354640 4904 354646 4916
rect 426342 4904 426348 4916
rect 426400 4904 426406 4956
rect 429102 4904 429108 4956
rect 429160 4944 429166 4956
rect 572622 4944 572628 4956
rect 429160 4916 572628 4944
rect 429160 4904 429166 4916
rect 572622 4904 572628 4916
rect 572680 4904 572686 4956
rect 12434 4836 12440 4888
rect 12492 4876 12498 4888
rect 139486 4876 139492 4888
rect 12492 4848 139492 4876
rect 12492 4836 12498 4848
rect 139486 4836 139492 4848
rect 139544 4836 139550 4888
rect 145650 4836 145656 4888
rect 145708 4876 145714 4888
rect 208578 4876 208584 4888
rect 145708 4848 208584 4876
rect 145708 4836 145714 4848
rect 208578 4836 208584 4848
rect 208636 4836 208642 4888
rect 212258 4836 212264 4888
rect 212316 4876 212322 4888
rect 242986 4876 242992 4888
rect 212316 4848 242992 4876
rect 212316 4836 212322 4848
rect 242986 4836 242992 4848
rect 243044 4836 243050 4888
rect 314562 4836 314568 4888
rect 314620 4876 314626 4888
rect 349062 4876 349068 4888
rect 314620 4848 349068 4876
rect 314620 4836 314626 4848
rect 349062 4836 349068 4848
rect 349120 4836 349126 4888
rect 351730 4836 351736 4888
rect 351788 4876 351794 4888
rect 422754 4876 422760 4888
rect 351788 4848 422760 4876
rect 351788 4836 351794 4848
rect 422754 4836 422760 4848
rect 422812 4836 422818 4888
rect 431862 4836 431868 4888
rect 431920 4876 431926 4888
rect 576210 4876 576216 4888
rect 431920 4848 576216 4876
rect 431920 4836 431926 4848
rect 576210 4836 576216 4848
rect 576268 4836 576274 4888
rect 4062 4768 4068 4820
rect 4120 4808 4126 4820
rect 135254 4808 135260 4820
rect 4120 4780 135260 4808
rect 4120 4768 4126 4780
rect 135254 4768 135260 4780
rect 135312 4768 135318 4820
rect 142062 4768 142068 4820
rect 142120 4808 142126 4820
rect 207014 4808 207020 4820
rect 142120 4780 207020 4808
rect 142120 4768 142126 4780
rect 207014 4768 207020 4780
rect 207072 4768 207078 4820
rect 208210 4768 208216 4820
rect 208268 4808 208274 4820
rect 238938 4808 238944 4820
rect 208268 4780 238944 4808
rect 208268 4768 208274 4780
rect 238938 4768 238944 4780
rect 238996 4768 239002 4820
rect 313090 4768 313096 4820
rect 313148 4808 313154 4820
rect 347866 4808 347872 4820
rect 313148 4780 347872 4808
rect 313148 4768 313154 4780
rect 347866 4768 347872 4780
rect 347924 4768 347930 4820
rect 355962 4768 355968 4820
rect 356020 4808 356026 4820
rect 429930 4808 429936 4820
rect 356020 4780 429936 4808
rect 356020 4768 356026 4780
rect 429930 4768 429936 4780
rect 429988 4768 429994 4820
rect 433242 4768 433248 4820
rect 433300 4808 433306 4820
rect 579798 4808 579804 4820
rect 433300 4780 579804 4808
rect 433300 4768 433306 4780
rect 579798 4768 579804 4780
rect 579856 4768 579862 4820
rect 73062 4700 73068 4752
rect 73120 4740 73126 4752
rect 171226 4740 171232 4752
rect 73120 4712 171232 4740
rect 73120 4700 73126 4712
rect 171226 4700 171232 4712
rect 171284 4700 171290 4752
rect 173894 4700 173900 4752
rect 173952 4740 173958 4752
rect 211246 4740 211252 4752
rect 173952 4712 211252 4740
rect 173952 4700 173958 4712
rect 211246 4700 211252 4712
rect 211304 4700 211310 4752
rect 338022 4700 338028 4752
rect 338080 4740 338086 4752
rect 394234 4740 394240 4752
rect 338080 4712 394240 4740
rect 338080 4700 338086 4712
rect 394234 4700 394240 4712
rect 394292 4700 394298 4752
rect 412542 4700 412548 4752
rect 412600 4740 412606 4752
rect 540514 4740 540520 4752
rect 412600 4712 540520 4740
rect 412600 4700 412606 4712
rect 540514 4700 540520 4712
rect 540572 4700 540578 4752
rect 76650 4632 76656 4684
rect 76708 4672 76714 4684
rect 172514 4672 172520 4684
rect 76708 4644 172520 4672
rect 76708 4632 76714 4644
rect 172514 4632 172520 4644
rect 172572 4632 172578 4684
rect 208670 4632 208676 4684
rect 208728 4672 208734 4684
rect 240134 4672 240140 4684
rect 208728 4644 240140 4672
rect 208728 4632 208734 4644
rect 240134 4632 240140 4644
rect 240192 4632 240198 4684
rect 333790 4632 333796 4684
rect 333848 4672 333854 4684
rect 387058 4672 387064 4684
rect 333848 4644 387064 4672
rect 333848 4632 333854 4644
rect 387058 4632 387064 4644
rect 387116 4632 387122 4684
rect 411162 4632 411168 4684
rect 411220 4672 411226 4684
rect 536926 4672 536932 4684
rect 411220 4644 536932 4672
rect 411220 4632 411226 4644
rect 536926 4632 536932 4644
rect 536984 4632 536990 4684
rect 80238 4564 80244 4616
rect 80296 4604 80302 4616
rect 175366 4604 175372 4616
rect 80296 4576 175372 4604
rect 80296 4564 80302 4576
rect 175366 4564 175372 4576
rect 175424 4564 175430 4616
rect 202874 4564 202880 4616
rect 202932 4604 202938 4616
rect 233326 4604 233332 4616
rect 202932 4576 233332 4604
rect 202932 4564 202938 4576
rect 233326 4564 233332 4576
rect 233384 4564 233390 4616
rect 329742 4564 329748 4616
rect 329800 4604 329806 4616
rect 379974 4604 379980 4616
rect 329800 4576 379980 4604
rect 329800 4564 329806 4576
rect 379974 4564 379980 4576
rect 380032 4564 380038 4616
rect 409782 4564 409788 4616
rect 409840 4604 409846 4616
rect 533430 4604 533436 4616
rect 409840 4576 533436 4604
rect 409840 4564 409846 4576
rect 533430 4564 533436 4576
rect 533488 4564 533494 4616
rect 83826 4496 83832 4548
rect 83884 4536 83890 4548
rect 176746 4536 176752 4548
rect 83884 4508 176752 4536
rect 83884 4496 83890 4508
rect 176746 4496 176752 4508
rect 176804 4496 176810 4548
rect 204254 4496 204260 4548
rect 204312 4536 204318 4548
rect 234706 4536 234712 4548
rect 204312 4508 234712 4536
rect 204312 4496 204318 4508
rect 234706 4496 234712 4508
rect 234764 4496 234770 4548
rect 332502 4496 332508 4548
rect 332560 4536 332566 4548
rect 383562 4536 383568 4548
rect 332560 4508 383568 4536
rect 332560 4496 332566 4508
rect 383562 4496 383568 4508
rect 383620 4496 383626 4548
rect 406930 4496 406936 4548
rect 406988 4536 406994 4548
rect 529842 4536 529848 4548
rect 406988 4508 529848 4536
rect 406988 4496 406994 4508
rect 529842 4496 529848 4508
rect 529900 4496 529906 4548
rect 49326 4428 49332 4480
rect 49384 4468 49390 4480
rect 130378 4468 130384 4480
rect 49384 4440 130384 4468
rect 49384 4428 49390 4440
rect 130378 4428 130384 4440
rect 130436 4428 130442 4480
rect 163498 4428 163504 4480
rect 163556 4468 163562 4480
rect 218146 4468 218152 4480
rect 163556 4440 218152 4468
rect 163556 4428 163562 4440
rect 218146 4428 218152 4440
rect 218204 4428 218210 4480
rect 328270 4428 328276 4480
rect 328328 4468 328334 4480
rect 376386 4468 376392 4480
rect 328328 4440 376392 4468
rect 328328 4428 328334 4440
rect 376386 4428 376392 4440
rect 376444 4428 376450 4480
rect 405642 4428 405648 4480
rect 405700 4468 405706 4480
rect 526254 4468 526260 4480
rect 405700 4440 526260 4468
rect 405700 4428 405706 4440
rect 526254 4428 526260 4440
rect 526312 4428 526318 4480
rect 45738 4360 45744 4412
rect 45796 4400 45802 4412
rect 126238 4400 126244 4412
rect 45796 4372 126244 4400
rect 45796 4360 45802 4372
rect 126238 4360 126244 4372
rect 126296 4360 126302 4412
rect 169665 4403 169723 4409
rect 169665 4369 169677 4403
rect 169711 4400 169723 4403
rect 205637 4403 205695 4409
rect 205637 4400 205649 4403
rect 169711 4372 205649 4400
rect 169711 4369 169723 4372
rect 169665 4363 169723 4369
rect 205637 4369 205649 4372
rect 205683 4369 205695 4403
rect 205637 4363 205695 4369
rect 326982 4360 326988 4412
rect 327040 4400 327046 4412
rect 372798 4400 372804 4412
rect 327040 4372 372804 4400
rect 327040 4360 327046 4372
rect 372798 4360 372804 4372
rect 372856 4360 372862 4412
rect 401502 4360 401508 4412
rect 401560 4400 401566 4412
rect 519078 4400 519084 4412
rect 401560 4372 519084 4400
rect 401560 4360 401566 4372
rect 519078 4360 519084 4372
rect 519136 4360 519142 4412
rect 52822 4292 52828 4344
rect 52880 4332 52886 4344
rect 122098 4332 122104 4344
rect 52880 4304 122104 4332
rect 52880 4292 52886 4304
rect 122098 4292 122104 4304
rect 122156 4292 122162 4344
rect 164694 4292 164700 4344
rect 164752 4332 164758 4344
rect 218054 4332 218060 4344
rect 164752 4304 218060 4332
rect 164752 4292 164758 4304
rect 218054 4292 218060 4304
rect 218112 4292 218118 4344
rect 324130 4292 324136 4344
rect 324188 4332 324194 4344
rect 369118 4332 369124 4344
rect 324188 4304 369124 4332
rect 324188 4292 324194 4304
rect 369118 4292 369124 4304
rect 369176 4292 369182 4344
rect 404262 4292 404268 4344
rect 404320 4332 404326 4344
rect 522666 4332 522672 4344
rect 404320 4304 522672 4332
rect 404320 4292 404326 4304
rect 522666 4292 522672 4304
rect 522724 4292 522730 4344
rect 63586 4224 63592 4276
rect 63644 4264 63650 4276
rect 128814 4264 128820 4276
rect 63644 4236 128820 4264
rect 63644 4224 63650 4236
rect 128814 4224 128820 4236
rect 128872 4224 128878 4276
rect 205637 4267 205695 4273
rect 205637 4233 205649 4267
rect 205683 4264 205695 4267
rect 215294 4264 215300 4276
rect 205683 4236 215300 4264
rect 205683 4233 205695 4236
rect 205637 4227 205695 4233
rect 215294 4224 215300 4236
rect 215352 4224 215358 4276
rect 322566 4224 322572 4276
rect 322624 4264 322630 4276
rect 365714 4264 365720 4276
rect 322624 4236 365720 4264
rect 322624 4224 322630 4236
rect 365714 4224 365720 4236
rect 365772 4224 365778 4276
rect 400030 4224 400036 4276
rect 400088 4264 400094 4276
rect 515582 4264 515588 4276
rect 400088 4236 515588 4264
rect 400088 4224 400094 4236
rect 515582 4224 515588 4236
rect 515640 4224 515646 4276
rect 67177 4199 67235 4205
rect 67177 4165 67189 4199
rect 67223 4196 67235 4199
rect 67542 4196 67548 4208
rect 67223 4168 67548 4196
rect 67223 4165 67235 4168
rect 67177 4159 67235 4165
rect 67542 4156 67548 4168
rect 67600 4156 67606 4208
rect 70670 4156 70676 4208
rect 70728 4196 70734 4208
rect 120718 4196 120724 4208
rect 70728 4168 120724 4196
rect 70728 4156 70734 4168
rect 120718 4156 120724 4168
rect 120776 4156 120782 4208
rect 169665 4199 169723 4205
rect 169665 4196 169677 4199
rect 161492 4168 169677 4196
rect 42150 4088 42156 4140
rect 42208 4128 42214 4140
rect 151906 4128 151912 4140
rect 42208 4100 151912 4128
rect 42208 4088 42214 4100
rect 151906 4088 151912 4100
rect 151964 4088 151970 4140
rect 159910 4088 159916 4140
rect 159968 4128 159974 4140
rect 161492 4128 161520 4168
rect 169665 4165 169677 4168
rect 169711 4165 169723 4199
rect 169665 4159 169723 4165
rect 321370 4156 321376 4208
rect 321428 4196 321434 4208
rect 362126 4196 362132 4208
rect 321428 4168 362132 4196
rect 321428 4156 321434 4168
rect 362126 4156 362132 4168
rect 362184 4156 362190 4208
rect 398742 4156 398748 4208
rect 398800 4196 398806 4208
rect 511994 4196 512000 4208
rect 398800 4168 512000 4196
rect 398800 4156 398806 4168
rect 511994 4156 512000 4168
rect 512052 4156 512058 4208
rect 159968 4100 161520 4128
rect 159968 4088 159974 4100
rect 168190 4088 168196 4140
rect 168248 4128 168254 4140
rect 174538 4128 174544 4140
rect 168248 4100 174544 4128
rect 168248 4088 168254 4100
rect 174538 4088 174544 4100
rect 174596 4088 174602 4140
rect 175366 4088 175372 4140
rect 175424 4128 175430 4140
rect 176562 4128 176568 4140
rect 175424 4100 176568 4128
rect 175424 4088 175430 4100
rect 176562 4088 176568 4100
rect 176620 4088 176626 4140
rect 177758 4088 177764 4140
rect 177816 4128 177822 4140
rect 180058 4128 180064 4140
rect 177816 4100 180064 4128
rect 177816 4088 177822 4100
rect 180058 4088 180064 4100
rect 180116 4088 180122 4140
rect 182542 4088 182548 4140
rect 182600 4128 182606 4140
rect 183462 4128 183468 4140
rect 182600 4100 183468 4128
rect 182600 4088 182606 4100
rect 183462 4088 183468 4100
rect 183520 4088 183526 4140
rect 190822 4088 190828 4140
rect 190880 4128 190886 4140
rect 190880 4100 225184 4128
rect 190880 4088 190886 4100
rect 43346 4020 43352 4072
rect 43404 4060 43410 4072
rect 155954 4060 155960 4072
rect 43404 4032 155960 4060
rect 43404 4020 43410 4032
rect 155954 4020 155960 4032
rect 156012 4020 156018 4072
rect 187234 4020 187240 4072
rect 187292 4060 187298 4072
rect 225049 4063 225107 4069
rect 225049 4060 225061 4063
rect 187292 4032 225061 4060
rect 187292 4020 187298 4032
rect 225049 4029 225061 4032
rect 225095 4029 225107 4063
rect 225049 4023 225107 4029
rect 39758 3952 39764 4004
rect 39816 3992 39822 4004
rect 153194 3992 153200 4004
rect 39816 3964 153200 3992
rect 39816 3952 39822 3964
rect 153194 3952 153200 3964
rect 153252 3952 153258 4004
rect 171778 3952 171784 4004
rect 171836 3992 171842 4004
rect 183554 3992 183560 4004
rect 171836 3964 183560 3992
rect 171836 3952 171842 3964
rect 183554 3952 183560 3964
rect 183612 3952 183618 4004
rect 188430 3952 188436 4004
rect 188488 3992 188494 4004
rect 220081 3995 220139 4001
rect 220081 3992 220093 3995
rect 188488 3964 220093 3992
rect 188488 3952 188494 3964
rect 220081 3961 220093 3964
rect 220127 3961 220139 3995
rect 225156 3992 225184 4100
rect 225322 4088 225328 4140
rect 225380 4128 225386 4140
rect 226242 4128 226248 4140
rect 225380 4100 226248 4128
rect 225380 4088 225386 4100
rect 226242 4088 226248 4100
rect 226300 4088 226306 4140
rect 226518 4088 226524 4140
rect 226576 4128 226582 4140
rect 227622 4128 227628 4140
rect 226576 4100 227628 4128
rect 226576 4088 226582 4100
rect 227622 4088 227628 4100
rect 227680 4088 227686 4140
rect 227714 4088 227720 4140
rect 227772 4128 227778 4140
rect 229002 4128 229008 4140
rect 227772 4100 229008 4128
rect 227772 4088 227778 4100
rect 229002 4088 229008 4100
rect 229060 4088 229066 4140
rect 231302 4088 231308 4140
rect 231360 4128 231366 4140
rect 231762 4128 231768 4140
rect 231360 4100 231768 4128
rect 231360 4088 231366 4100
rect 231762 4088 231768 4100
rect 231820 4088 231826 4140
rect 233694 4088 233700 4140
rect 233752 4128 233758 4140
rect 234522 4128 234528 4140
rect 233752 4100 234528 4128
rect 233752 4088 233758 4100
rect 234522 4088 234528 4100
rect 234580 4088 234586 4140
rect 239582 4088 239588 4140
rect 239640 4128 239646 4140
rect 240042 4128 240048 4140
rect 239640 4100 240048 4128
rect 239640 4088 239646 4100
rect 240042 4088 240048 4100
rect 240100 4088 240106 4140
rect 243170 4088 243176 4140
rect 243228 4128 243234 4140
rect 244182 4128 244188 4140
rect 243228 4100 244188 4128
rect 243228 4088 243234 4100
rect 244182 4088 244188 4100
rect 244240 4088 244246 4140
rect 244366 4088 244372 4140
rect 244424 4128 244430 4140
rect 245562 4128 245568 4140
rect 244424 4100 245568 4128
rect 244424 4088 244430 4100
rect 245562 4088 245568 4100
rect 245620 4088 245626 4140
rect 246758 4088 246764 4140
rect 246816 4128 246822 4140
rect 247678 4128 247684 4140
rect 246816 4100 247684 4128
rect 246816 4088 246822 4100
rect 247678 4088 247684 4100
rect 247736 4088 247742 4140
rect 249150 4088 249156 4140
rect 249208 4128 249214 4140
rect 249702 4128 249708 4140
rect 249208 4100 249708 4128
rect 249208 4088 249214 4100
rect 249702 4088 249708 4100
rect 249760 4088 249766 4140
rect 251450 4088 251456 4140
rect 251508 4128 251514 4140
rect 252462 4128 252468 4140
rect 251508 4100 252468 4128
rect 251508 4088 251514 4100
rect 252462 4088 252468 4100
rect 252520 4088 252526 4140
rect 265802 4088 265808 4140
rect 265860 4128 265866 4140
rect 266262 4128 266268 4140
rect 265860 4100 266268 4128
rect 265860 4088 265866 4100
rect 266262 4088 266268 4100
rect 266320 4088 266326 4140
rect 268102 4088 268108 4140
rect 268160 4128 268166 4140
rect 269758 4128 269764 4140
rect 268160 4100 269764 4128
rect 268160 4088 268166 4100
rect 269758 4088 269764 4100
rect 269816 4088 269822 4140
rect 271690 4088 271696 4140
rect 271748 4128 271754 4140
rect 272518 4128 272524 4140
rect 271748 4100 272524 4128
rect 271748 4088 271754 4100
rect 272518 4088 272524 4100
rect 272576 4088 272582 4140
rect 274082 4088 274088 4140
rect 274140 4128 274146 4140
rect 274542 4128 274548 4140
rect 274140 4100 274548 4128
rect 274140 4088 274146 4100
rect 274542 4088 274548 4100
rect 274600 4088 274606 4140
rect 277302 4088 277308 4140
rect 277360 4128 277366 4140
rect 277670 4128 277676 4140
rect 277360 4100 277676 4128
rect 277360 4088 277366 4100
rect 277670 4088 277676 4100
rect 277728 4088 277734 4140
rect 280062 4088 280068 4140
rect 280120 4128 280126 4140
rect 282454 4128 282460 4140
rect 280120 4100 282460 4128
rect 280120 4088 280126 4100
rect 282454 4088 282460 4100
rect 282512 4088 282518 4140
rect 292390 4088 292396 4140
rect 292448 4128 292454 4140
rect 307386 4128 307392 4140
rect 292448 4100 307392 4128
rect 292448 4088 292454 4100
rect 307386 4088 307392 4100
rect 307444 4088 307450 4140
rect 315298 4088 315304 4140
rect 315356 4128 315362 4140
rect 315850 4128 315856 4140
rect 315356 4100 315856 4128
rect 315356 4088 315362 4100
rect 315850 4088 315856 4100
rect 315908 4088 315914 4140
rect 321462 4088 321468 4140
rect 321520 4128 321526 4140
rect 363322 4128 363328 4140
rect 321520 4100 363328 4128
rect 321520 4088 321526 4100
rect 363322 4088 363328 4100
rect 363380 4088 363386 4140
rect 363598 4088 363604 4140
rect 363656 4128 363662 4140
rect 364518 4128 364524 4140
rect 363656 4100 364524 4128
rect 363656 4088 363662 4100
rect 364518 4088 364524 4100
rect 364576 4088 364582 4140
rect 391750 4088 391756 4140
rect 391808 4128 391814 4140
rect 500126 4128 500132 4140
rect 391808 4100 500132 4128
rect 391808 4088 391814 4100
rect 500126 4088 500132 4100
rect 500184 4088 500190 4140
rect 502978 4088 502984 4140
rect 503036 4128 503042 4140
rect 507029 4131 507087 4137
rect 507029 4128 507041 4131
rect 503036 4100 507041 4128
rect 503036 4088 503042 4100
rect 507029 4097 507041 4100
rect 507075 4097 507087 4131
rect 507029 4091 507087 4097
rect 507118 4088 507124 4140
rect 507176 4128 507182 4140
rect 571426 4128 571432 4140
rect 507176 4100 571432 4128
rect 507176 4088 507182 4100
rect 571426 4088 571432 4100
rect 571484 4088 571490 4140
rect 241974 4020 241980 4072
rect 242032 4060 242038 4072
rect 243722 4060 243728 4072
rect 242032 4032 243728 4060
rect 242032 4020 242038 4032
rect 243722 4020 243728 4032
rect 243780 4020 243786 4072
rect 284202 4020 284208 4072
rect 284260 4060 284266 4072
rect 289538 4060 289544 4072
rect 284260 4032 289544 4060
rect 284260 4020 284266 4032
rect 289538 4020 289544 4032
rect 289596 4020 289602 4072
rect 297910 4020 297916 4072
rect 297968 4020 297974 4072
rect 298002 4020 298008 4072
rect 298060 4060 298066 4072
rect 316954 4060 316960 4072
rect 298060 4032 316960 4060
rect 298060 4020 298066 4032
rect 316954 4020 316960 4032
rect 317012 4020 317018 4072
rect 322842 4020 322848 4072
rect 322900 4060 322906 4072
rect 361025 4063 361083 4069
rect 361025 4060 361037 4063
rect 322900 4032 361037 4060
rect 322900 4020 322906 4032
rect 361025 4029 361037 4032
rect 361071 4029 361083 4063
rect 361025 4023 361083 4029
rect 395982 4020 395988 4072
rect 396040 4060 396046 4072
rect 507210 4060 507216 4072
rect 396040 4032 507216 4060
rect 396040 4020 396046 4032
rect 507210 4020 507216 4032
rect 507268 4020 507274 4072
rect 507305 4063 507363 4069
rect 507305 4029 507317 4063
rect 507351 4060 507363 4063
rect 514021 4063 514079 4069
rect 514021 4060 514033 4063
rect 507351 4032 514033 4060
rect 507351 4029 507363 4032
rect 507305 4023 507363 4029
rect 514021 4029 514033 4032
rect 514067 4029 514079 4063
rect 514021 4023 514079 4029
rect 514113 4063 514171 4069
rect 514113 4029 514125 4063
rect 514159 4060 514171 4063
rect 578602 4060 578608 4072
rect 514159 4032 578608 4060
rect 514159 4029 514171 4032
rect 514113 4023 514171 4029
rect 578602 4020 578608 4032
rect 578660 4020 578666 4072
rect 231946 3992 231952 4004
rect 225156 3964 231952 3992
rect 220081 3955 220139 3961
rect 231946 3952 231952 3964
rect 232004 3952 232010 4004
rect 269298 3952 269304 4004
rect 269356 3992 269362 4004
rect 272150 3992 272156 4004
rect 269356 3964 272156 3992
rect 269356 3952 269362 3964
rect 272150 3952 272156 3964
rect 272208 3952 272214 4004
rect 285582 3952 285588 4004
rect 285640 3992 285646 4004
rect 293126 3992 293132 4004
rect 285640 3964 293132 3992
rect 285640 3952 285646 3964
rect 293126 3952 293132 3964
rect 293184 3952 293190 4004
rect 297928 3992 297956 4020
rect 318058 3992 318064 4004
rect 297928 3964 318064 3992
rect 318058 3952 318064 3964
rect 318116 3952 318122 4004
rect 324222 3952 324228 4004
rect 324280 3992 324286 4004
rect 368014 3992 368020 4004
rect 324280 3964 368020 3992
rect 324280 3952 324286 3964
rect 368014 3952 368020 3964
rect 368072 3952 368078 4004
rect 400122 3952 400128 4004
rect 400180 3992 400186 4004
rect 514386 3992 514392 4004
rect 400180 3964 514392 3992
rect 400180 3952 400186 3964
rect 514386 3952 514392 3964
rect 514444 3952 514450 4004
rect 32674 3884 32680 3936
rect 32732 3924 32738 3936
rect 150434 3924 150440 3936
rect 32732 3896 150440 3924
rect 32732 3884 32738 3896
rect 150434 3884 150440 3896
rect 150492 3884 150498 3936
rect 161106 3884 161112 3936
rect 161164 3924 161170 3936
rect 178678 3924 178684 3936
rect 161164 3896 178684 3924
rect 161164 3884 161170 3896
rect 178678 3884 178684 3896
rect 178736 3884 178742 3936
rect 183738 3884 183744 3936
rect 183796 3924 183802 3936
rect 227898 3924 227904 3936
rect 183796 3896 227904 3924
rect 183796 3884 183802 3896
rect 227898 3884 227904 3896
rect 227956 3884 227962 3936
rect 235994 3884 236000 3936
rect 236052 3924 236058 3936
rect 237282 3924 237288 3936
rect 236052 3896 237288 3924
rect 236052 3884 236058 3896
rect 237282 3884 237288 3896
rect 237340 3884 237346 3936
rect 283558 3884 283564 3936
rect 283616 3924 283622 3936
rect 287146 3924 287152 3936
rect 283616 3896 287152 3924
rect 283616 3884 283622 3896
rect 287146 3884 287152 3896
rect 287204 3884 287210 3936
rect 288342 3884 288348 3936
rect 288400 3924 288406 3936
rect 297910 3924 297916 3936
rect 288400 3896 297916 3924
rect 288400 3884 288406 3896
rect 297910 3884 297916 3896
rect 297968 3884 297974 3936
rect 302142 3884 302148 3936
rect 302200 3924 302206 3936
rect 324038 3924 324044 3936
rect 302200 3896 324044 3924
rect 302200 3884 302206 3896
rect 324038 3884 324044 3896
rect 324096 3884 324102 3936
rect 326338 3884 326344 3936
rect 326396 3924 326402 3936
rect 370406 3924 370412 3936
rect 326396 3896 370412 3924
rect 326396 3884 326402 3896
rect 370406 3884 370412 3896
rect 370464 3884 370470 3936
rect 374638 3884 374644 3936
rect 374696 3924 374702 3936
rect 374696 3896 375420 3924
rect 374696 3884 374702 3896
rect 25498 3816 25504 3868
rect 25556 3856 25562 3868
rect 146294 3856 146300 3868
rect 25556 3828 146300 3856
rect 25556 3816 25562 3828
rect 146294 3816 146300 3828
rect 146352 3816 146358 3868
rect 157518 3816 157524 3868
rect 157576 3856 157582 3868
rect 177482 3856 177488 3868
rect 157576 3828 177488 3856
rect 157576 3816 157582 3828
rect 177482 3816 177488 3828
rect 177540 3816 177546 3868
rect 180150 3816 180156 3868
rect 180208 3856 180214 3868
rect 226426 3856 226432 3868
rect 180208 3828 226432 3856
rect 180208 3816 180214 3828
rect 226426 3816 226432 3828
rect 226484 3816 226490 3868
rect 228910 3816 228916 3868
rect 228968 3856 228974 3868
rect 235258 3856 235264 3868
rect 228968 3828 235264 3856
rect 228968 3816 228974 3828
rect 235258 3816 235264 3828
rect 235316 3816 235322 3868
rect 286870 3816 286876 3868
rect 286928 3856 286934 3868
rect 295518 3856 295524 3868
rect 286928 3828 295524 3856
rect 286928 3816 286934 3828
rect 295518 3816 295524 3828
rect 295576 3816 295582 3868
rect 299382 3816 299388 3868
rect 299440 3856 299446 3868
rect 320450 3856 320456 3868
rect 299440 3828 320456 3856
rect 299440 3816 299446 3828
rect 320450 3816 320456 3828
rect 320508 3816 320514 3868
rect 328362 3816 328368 3868
rect 328420 3856 328426 3868
rect 375190 3856 375196 3868
rect 328420 3828 375196 3856
rect 328420 3816 328426 3828
rect 375190 3816 375196 3828
rect 375248 3816 375254 3868
rect 375392 3856 375420 3896
rect 384298 3884 384304 3936
rect 384356 3924 384362 3936
rect 396626 3924 396632 3936
rect 384356 3896 396632 3924
rect 384356 3884 384362 3896
rect 396626 3884 396632 3896
rect 396684 3884 396690 3936
rect 402882 3884 402888 3936
rect 402940 3924 402946 3936
rect 521470 3924 521476 3936
rect 402940 3896 521476 3924
rect 402940 3884 402946 3896
rect 521470 3884 521476 3896
rect 521528 3884 521534 3936
rect 393038 3856 393044 3868
rect 375392 3828 393044 3856
rect 393038 3816 393044 3828
rect 393096 3816 393102 3868
rect 398837 3859 398895 3865
rect 398837 3825 398849 3859
rect 398883 3856 398895 3859
rect 398883 3828 403848 3856
rect 398883 3825 398895 3828
rect 398837 3819 398895 3825
rect 24302 3748 24308 3800
rect 24360 3788 24366 3800
rect 146386 3788 146392 3800
rect 24360 3760 146392 3788
rect 24360 3748 24366 3760
rect 146386 3748 146392 3760
rect 146444 3748 146450 3800
rect 151538 3748 151544 3800
rect 151596 3788 151602 3800
rect 173894 3788 173900 3800
rect 151596 3760 173900 3788
rect 151596 3748 151602 3760
rect 173894 3748 173900 3760
rect 173952 3748 173958 3800
rect 176470 3748 176476 3800
rect 176528 3788 176534 3800
rect 217965 3791 218023 3797
rect 217965 3788 217977 3791
rect 176528 3760 217977 3788
rect 176528 3748 176534 3760
rect 217965 3757 217977 3760
rect 218011 3757 218023 3791
rect 219713 3791 219771 3797
rect 219713 3788 219725 3791
rect 217965 3751 218023 3757
rect 218072 3760 219725 3788
rect 19518 3680 19524 3732
rect 19576 3720 19582 3732
rect 143534 3720 143540 3732
rect 19576 3692 143540 3720
rect 19576 3680 19582 3692
rect 143534 3680 143540 3692
rect 143592 3680 143598 3732
rect 172974 3680 172980 3732
rect 173032 3720 173038 3732
rect 218072 3720 218100 3760
rect 219713 3757 219725 3760
rect 219759 3757 219771 3791
rect 219713 3751 219771 3757
rect 220081 3791 220139 3797
rect 220081 3757 220093 3791
rect 220127 3788 220139 3791
rect 230566 3788 230572 3800
rect 220127 3760 230572 3788
rect 220127 3757 220139 3760
rect 220081 3751 220139 3757
rect 230566 3748 230572 3760
rect 230624 3748 230630 3800
rect 286962 3748 286968 3800
rect 287020 3788 287026 3800
rect 296714 3788 296720 3800
rect 287020 3760 296720 3788
rect 287020 3748 287026 3760
rect 296714 3748 296720 3760
rect 296772 3748 296778 3800
rect 302050 3748 302056 3800
rect 302108 3788 302114 3800
rect 325234 3788 325240 3800
rect 302108 3760 325240 3788
rect 302108 3748 302114 3760
rect 325234 3748 325240 3760
rect 325292 3748 325298 3800
rect 326154 3748 326160 3800
rect 326212 3788 326218 3800
rect 326433 3791 326491 3797
rect 326433 3788 326445 3791
rect 326212 3760 326445 3788
rect 326212 3748 326218 3760
rect 326433 3757 326445 3760
rect 326479 3757 326491 3791
rect 326433 3751 326491 3757
rect 334618 3748 334624 3800
rect 334676 3788 334682 3800
rect 335906 3788 335912 3800
rect 334676 3760 335912 3788
rect 334676 3748 334682 3760
rect 335906 3748 335912 3760
rect 335964 3748 335970 3800
rect 340141 3791 340199 3797
rect 340141 3757 340153 3791
rect 340187 3788 340199 3791
rect 382366 3788 382372 3800
rect 340187 3760 382372 3788
rect 340187 3757 340199 3760
rect 340141 3751 340199 3757
rect 382366 3748 382372 3760
rect 382424 3748 382430 3800
rect 389818 3748 389824 3800
rect 389876 3788 389882 3800
rect 403710 3788 403716 3800
rect 389876 3760 403716 3788
rect 389876 3748 389882 3760
rect 403710 3748 403716 3760
rect 403768 3748 403774 3800
rect 403820 3788 403848 3828
rect 407022 3816 407028 3868
rect 407080 3856 407086 3868
rect 528646 3856 528652 3868
rect 407080 3828 528652 3856
rect 407080 3816 407086 3828
rect 528646 3816 528652 3828
rect 528704 3816 528710 3868
rect 407393 3791 407451 3797
rect 407393 3788 407405 3791
rect 403820 3760 407405 3788
rect 407393 3757 407405 3760
rect 407439 3757 407451 3791
rect 407393 3751 407451 3757
rect 409506 3748 409512 3800
rect 409564 3788 409570 3800
rect 535730 3788 535736 3800
rect 409564 3760 535736 3788
rect 409564 3748 409570 3760
rect 535730 3748 535736 3760
rect 535788 3748 535794 3800
rect 173032 3692 218100 3720
rect 173032 3680 173038 3692
rect 218146 3680 218152 3732
rect 218204 3720 218210 3732
rect 224218 3720 224224 3732
rect 218204 3692 224224 3720
rect 218204 3680 218210 3692
rect 224218 3680 224224 3692
rect 224276 3680 224282 3732
rect 225049 3723 225107 3729
rect 225049 3689 225061 3723
rect 225095 3720 225107 3723
rect 229186 3720 229192 3732
rect 225095 3692 229192 3720
rect 225095 3689 225107 3692
rect 225049 3683 225107 3689
rect 229186 3680 229192 3692
rect 229244 3680 229250 3732
rect 288250 3680 288256 3732
rect 288308 3720 288314 3732
rect 299106 3720 299112 3732
rect 288308 3692 299112 3720
rect 288308 3680 288314 3692
rect 299106 3680 299112 3692
rect 299164 3680 299170 3732
rect 303522 3680 303528 3732
rect 303580 3720 303586 3732
rect 327626 3720 327632 3732
rect 303580 3692 327632 3720
rect 303580 3680 303586 3692
rect 327626 3680 327632 3692
rect 327684 3680 327690 3732
rect 333882 3680 333888 3732
rect 333940 3720 333946 3732
rect 385862 3720 385868 3732
rect 333940 3692 385868 3720
rect 333940 3680 333946 3692
rect 385862 3680 385868 3692
rect 385920 3680 385926 3732
rect 396718 3680 396724 3732
rect 396776 3720 396782 3732
rect 410886 3720 410892 3732
rect 396776 3692 410892 3720
rect 396776 3680 396782 3692
rect 410886 3680 410892 3692
rect 410944 3680 410950 3732
rect 418154 3680 418160 3732
rect 418212 3720 418218 3732
rect 542906 3720 542912 3732
rect 418212 3692 542912 3720
rect 418212 3680 418218 3692
rect 542906 3680 542912 3692
rect 542964 3680 542970 3732
rect 14826 3612 14832 3664
rect 14884 3652 14890 3664
rect 140774 3652 140780 3664
rect 14884 3624 140780 3652
rect 14884 3612 14890 3624
rect 140774 3612 140780 3624
rect 140832 3612 140838 3664
rect 148042 3612 148048 3664
rect 148100 3652 148106 3664
rect 196713 3655 196771 3661
rect 196713 3652 196725 3655
rect 148100 3624 196725 3652
rect 148100 3612 148106 3624
rect 196713 3621 196725 3624
rect 196759 3621 196771 3655
rect 196713 3615 196771 3621
rect 196802 3612 196808 3664
rect 196860 3652 196866 3664
rect 197262 3652 197268 3664
rect 196860 3624 197268 3652
rect 196860 3612 196866 3624
rect 197262 3612 197268 3624
rect 197320 3612 197326 3664
rect 200390 3612 200396 3664
rect 200448 3652 200454 3664
rect 201402 3652 201408 3664
rect 200448 3624 201408 3652
rect 200448 3612 200454 3624
rect 201402 3612 201408 3624
rect 201460 3612 201466 3664
rect 201494 3612 201500 3664
rect 201552 3652 201558 3664
rect 204346 3652 204352 3664
rect 201552 3624 204352 3652
rect 201552 3612 201558 3624
rect 204346 3612 204352 3624
rect 204404 3612 204410 3664
rect 207474 3612 207480 3664
rect 207532 3652 207538 3664
rect 208302 3652 208308 3664
rect 207532 3624 208308 3652
rect 207532 3612 207538 3624
rect 208302 3612 208308 3624
rect 208360 3612 208366 3664
rect 209866 3612 209872 3664
rect 209924 3652 209930 3664
rect 211062 3652 211068 3664
rect 209924 3624 211068 3652
rect 209924 3612 209930 3624
rect 211062 3612 211068 3624
rect 211120 3612 211126 3664
rect 211157 3655 211215 3661
rect 211157 3621 211169 3655
rect 211203 3652 211215 3655
rect 233878 3652 233884 3664
rect 211203 3624 233884 3652
rect 211203 3621 211215 3624
rect 211157 3615 211215 3621
rect 233878 3612 233884 3624
rect 233936 3612 233942 3664
rect 234798 3612 234804 3664
rect 234856 3652 234862 3664
rect 250438 3652 250444 3664
rect 234856 3624 250444 3652
rect 234856 3612 234862 3624
rect 250438 3612 250444 3624
rect 250496 3612 250502 3664
rect 284938 3612 284944 3664
rect 284996 3652 285002 3664
rect 288342 3652 288348 3664
rect 284996 3624 288348 3652
rect 284996 3612 285002 3624
rect 288342 3612 288348 3624
rect 288400 3612 288406 3664
rect 291010 3612 291016 3664
rect 291068 3652 291074 3664
rect 303798 3652 303804 3664
rect 291068 3624 303804 3652
rect 291068 3612 291074 3624
rect 303798 3612 303804 3624
rect 303856 3612 303862 3664
rect 306282 3612 306288 3664
rect 306340 3652 306346 3664
rect 332410 3652 332416 3664
rect 306340 3624 332416 3652
rect 306340 3612 306346 3624
rect 332410 3612 332416 3624
rect 332468 3612 332474 3664
rect 335262 3612 335268 3664
rect 335320 3652 335326 3664
rect 389450 3652 389456 3664
rect 335320 3624 389456 3652
rect 335320 3612 335326 3624
rect 389450 3612 389456 3624
rect 389508 3612 389514 3664
rect 393958 3612 393964 3664
rect 394016 3652 394022 3664
rect 398837 3655 398895 3661
rect 398837 3652 398849 3655
rect 394016 3624 398849 3652
rect 394016 3612 394022 3624
rect 398837 3621 398849 3624
rect 398883 3621 398895 3655
rect 398837 3615 398895 3621
rect 413186 3612 413192 3664
rect 413244 3652 413250 3664
rect 417973 3655 418031 3661
rect 417973 3652 417985 3655
rect 413244 3624 417985 3652
rect 413244 3612 413250 3624
rect 417973 3621 417985 3624
rect 418019 3621 418031 3655
rect 417973 3615 418031 3621
rect 420178 3612 420184 3664
rect 420236 3652 420242 3664
rect 553578 3652 553584 3664
rect 420236 3624 553584 3652
rect 420236 3612 420242 3624
rect 553578 3612 553584 3624
rect 553636 3612 553642 3664
rect 16022 3544 16028 3596
rect 16080 3584 16086 3596
rect 142338 3584 142344 3596
rect 16080 3556 142344 3584
rect 16080 3544 16086 3556
rect 142338 3544 142344 3556
rect 142396 3544 142402 3596
rect 169386 3544 169392 3596
rect 169444 3584 169450 3596
rect 210421 3587 210479 3593
rect 210421 3584 210433 3587
rect 169444 3556 210433 3584
rect 169444 3544 169450 3556
rect 210421 3553 210433 3556
rect 210467 3553 210479 3587
rect 210421 3547 210479 3553
rect 214650 3544 214656 3596
rect 214708 3584 214714 3596
rect 220078 3584 220084 3596
rect 214708 3556 220084 3584
rect 214708 3544 214714 3556
rect 220078 3544 220084 3556
rect 220136 3544 220142 3596
rect 224126 3544 224132 3596
rect 224184 3584 224190 3596
rect 248506 3584 248512 3596
rect 224184 3556 248512 3584
rect 224184 3544 224190 3556
rect 248506 3544 248512 3556
rect 248564 3544 248570 3596
rect 291102 3544 291108 3596
rect 291160 3584 291166 3596
rect 302602 3584 302608 3596
rect 291160 3556 302608 3584
rect 291160 3544 291166 3556
rect 302602 3544 302608 3556
rect 302660 3544 302666 3596
rect 303430 3544 303436 3596
rect 303488 3584 303494 3596
rect 328822 3584 328828 3596
rect 303488 3556 328828 3584
rect 303488 3544 303494 3556
rect 328822 3544 328828 3556
rect 328880 3544 328886 3596
rect 331122 3544 331128 3596
rect 331180 3584 331186 3596
rect 340141 3587 340199 3593
rect 340141 3584 340153 3587
rect 331180 3556 340153 3584
rect 331180 3544 331186 3556
rect 340141 3553 340153 3556
rect 340187 3553 340199 3587
rect 340141 3547 340199 3553
rect 341610 3544 341616 3596
rect 341668 3584 341674 3596
rect 343082 3584 343088 3596
rect 341668 3556 343088 3584
rect 341668 3544 341674 3556
rect 343082 3544 343088 3556
rect 343140 3544 343146 3596
rect 358170 3544 358176 3596
rect 358228 3584 358234 3596
rect 360930 3584 360936 3596
rect 358228 3556 360936 3584
rect 358228 3544 358234 3556
rect 360930 3544 360936 3556
rect 360988 3544 360994 3596
rect 361025 3587 361083 3593
rect 361025 3553 361037 3587
rect 361071 3584 361083 3587
rect 366910 3584 366916 3596
rect 361071 3556 366916 3584
rect 361071 3553 361083 3556
rect 361025 3547 361083 3553
rect 366910 3544 366916 3556
rect 366968 3544 366974 3596
rect 369210 3544 369216 3596
rect 369268 3584 369274 3596
rect 371602 3584 371608 3596
rect 369268 3556 371608 3584
rect 369268 3544 369274 3556
rect 371602 3544 371608 3556
rect 371660 3544 371666 3596
rect 398098 3544 398104 3596
rect 398156 3584 398162 3596
rect 408310 3584 408316 3596
rect 398156 3556 408316 3584
rect 398156 3544 398162 3556
rect 408310 3544 408316 3556
rect 408368 3544 408374 3596
rect 408494 3544 408500 3596
rect 408552 3584 408558 3596
rect 408552 3556 422984 3584
rect 408552 3544 408558 3556
rect 8846 3476 8852 3528
rect 8904 3516 8910 3528
rect 9582 3516 9588 3528
rect 8904 3488 9588 3516
rect 8904 3476 8910 3488
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 10042 3476 10048 3528
rect 10100 3516 10106 3528
rect 138014 3516 138020 3528
rect 10100 3488 138020 3516
rect 10100 3476 10106 3488
rect 138014 3476 138020 3488
rect 138072 3476 138078 3528
rect 154577 3519 154635 3525
rect 154577 3485 154589 3519
rect 154623 3516 154635 3519
rect 164145 3519 164203 3525
rect 164145 3516 164157 3519
rect 154623 3488 164157 3516
rect 154623 3485 154635 3488
rect 154577 3479 154635 3485
rect 164145 3485 164157 3488
rect 164191 3485 164203 3519
rect 164145 3479 164203 3485
rect 165890 3476 165896 3528
rect 165948 3516 165954 3528
rect 219618 3516 219624 3528
rect 165948 3488 219624 3516
rect 165948 3476 165954 3488
rect 219618 3476 219624 3488
rect 219676 3476 219682 3528
rect 219713 3519 219771 3525
rect 219713 3485 219725 3519
rect 219759 3516 219771 3519
rect 222194 3516 222200 3528
rect 219759 3488 222200 3516
rect 219759 3485 219771 3488
rect 219713 3479 219771 3485
rect 222194 3476 222200 3488
rect 222252 3476 222258 3528
rect 222930 3476 222936 3528
rect 222988 3516 222994 3528
rect 248598 3516 248604 3528
rect 222988 3488 248604 3516
rect 222988 3476 222994 3488
rect 248598 3476 248604 3488
rect 248656 3476 248662 3528
rect 257430 3476 257436 3528
rect 257488 3516 257494 3528
rect 257982 3516 257988 3528
rect 257488 3488 257988 3516
rect 257488 3476 257494 3488
rect 257982 3476 257988 3488
rect 258040 3476 258046 3528
rect 259822 3476 259828 3528
rect 259880 3516 259886 3528
rect 261478 3516 261484 3528
rect 259880 3488 261484 3516
rect 259880 3476 259886 3488
rect 261478 3476 261484 3488
rect 261536 3476 261542 3528
rect 262214 3476 262220 3528
rect 262272 3516 262278 3528
rect 263502 3516 263508 3528
rect 262272 3488 263508 3516
rect 262272 3476 262278 3488
rect 263502 3476 263508 3488
rect 263560 3476 263566 3528
rect 290918 3476 290924 3528
rect 290976 3516 290982 3528
rect 304994 3516 305000 3528
rect 290976 3488 305000 3516
rect 290976 3476 290982 3488
rect 304994 3476 305000 3488
rect 305052 3476 305058 3528
rect 305638 3476 305644 3528
rect 305696 3516 305702 3528
rect 306282 3516 306288 3528
rect 305696 3488 306288 3516
rect 305696 3476 305702 3488
rect 306282 3476 306288 3488
rect 306340 3476 306346 3528
rect 309042 3476 309048 3528
rect 309100 3516 309106 3528
rect 339494 3516 339500 3528
rect 309100 3488 339500 3516
rect 309100 3476 309106 3488
rect 339494 3476 339500 3488
rect 339552 3476 339558 3528
rect 344922 3476 344928 3528
rect 344980 3516 344986 3528
rect 407298 3516 407304 3528
rect 344980 3488 407304 3516
rect 344980 3476 344986 3488
rect 407298 3476 407304 3488
rect 407356 3476 407362 3528
rect 407393 3519 407451 3525
rect 407393 3485 407405 3519
rect 407439 3516 407451 3519
rect 417878 3516 417884 3528
rect 407439 3488 417884 3516
rect 407439 3485 407451 3488
rect 407393 3479 407451 3485
rect 417878 3476 417884 3488
rect 417936 3476 417942 3528
rect 417973 3519 418031 3525
rect 417973 3485 417985 3519
rect 418019 3516 418031 3519
rect 418157 3519 418215 3525
rect 418157 3516 418169 3519
rect 418019 3488 418169 3516
rect 418019 3485 418031 3488
rect 417973 3479 418031 3485
rect 418157 3485 418169 3488
rect 418203 3485 418215 3519
rect 421558 3516 421564 3528
rect 418157 3479 418215 3485
rect 418264 3488 421564 3516
rect 11238 3408 11244 3460
rect 11296 3448 11302 3460
rect 139578 3448 139584 3460
rect 11296 3420 139584 3448
rect 11296 3408 11302 3420
rect 139578 3408 139584 3420
rect 139636 3408 139642 3460
rect 147677 3451 147735 3457
rect 147677 3417 147689 3451
rect 147723 3448 147735 3451
rect 147723 3420 159404 3448
rect 147723 3417 147735 3420
rect 147677 3411 147735 3417
rect 27890 3340 27896 3392
rect 27948 3380 27954 3392
rect 28902 3380 28908 3392
rect 27948 3352 28908 3380
rect 27948 3340 27954 3352
rect 28902 3340 28908 3352
rect 28960 3340 28966 3392
rect 50522 3340 50528 3392
rect 50580 3380 50586 3392
rect 159082 3380 159088 3392
rect 50580 3352 159088 3380
rect 50580 3340 50586 3352
rect 159082 3340 159088 3352
rect 159140 3340 159146 3392
rect 59998 3272 60004 3324
rect 60056 3312 60062 3324
rect 60642 3312 60648 3324
rect 60056 3284 60648 3312
rect 60056 3272 60062 3284
rect 60642 3272 60648 3284
rect 60700 3272 60706 3324
rect 62761 3315 62819 3321
rect 62761 3281 62773 3315
rect 62807 3312 62819 3315
rect 62807 3284 73200 3312
rect 62807 3281 62819 3284
rect 62761 3275 62819 3281
rect 38562 3204 38568 3256
rect 38620 3244 38626 3256
rect 38620 3216 41460 3244
rect 38620 3204 38626 3216
rect 41432 3176 41460 3216
rect 57977 3179 58035 3185
rect 57977 3176 57989 3179
rect 41432 3148 57989 3176
rect 57977 3145 57989 3148
rect 58023 3145 58035 3179
rect 73172 3176 73200 3284
rect 81434 3272 81440 3324
rect 81492 3312 81498 3324
rect 82538 3312 82544 3324
rect 81492 3284 82544 3312
rect 81492 3272 81498 3284
rect 82538 3272 82544 3284
rect 82596 3272 82602 3324
rect 82630 3272 82636 3324
rect 82688 3312 82694 3324
rect 103517 3315 103575 3321
rect 103517 3312 103529 3315
rect 82688 3284 103529 3312
rect 82688 3272 82694 3284
rect 103517 3281 103529 3284
rect 103563 3281 103575 3315
rect 103517 3275 103575 3281
rect 110601 3315 110659 3321
rect 110601 3281 110613 3315
rect 110647 3312 110659 3315
rect 122837 3315 122895 3321
rect 122837 3312 122849 3315
rect 110647 3284 122849 3312
rect 110647 3281 110659 3284
rect 110601 3275 110659 3281
rect 122837 3281 122849 3284
rect 122883 3281 122895 3315
rect 122837 3275 122895 3281
rect 132586 3272 132592 3324
rect 132644 3312 132650 3324
rect 133138 3312 133144 3324
rect 132644 3284 133144 3312
rect 132644 3272 132650 3284
rect 133138 3272 133144 3284
rect 133196 3272 133202 3324
rect 137925 3315 137983 3321
rect 137925 3281 137937 3315
rect 137971 3312 137983 3315
rect 147677 3315 147735 3321
rect 147677 3312 147689 3315
rect 137971 3284 147689 3312
rect 137971 3281 137983 3284
rect 137925 3275 137983 3281
rect 147677 3281 147689 3284
rect 147723 3281 147735 3315
rect 159376 3312 159404 3420
rect 162302 3408 162308 3460
rect 162360 3448 162366 3460
rect 208857 3451 208915 3457
rect 208857 3448 208869 3451
rect 162360 3420 208869 3448
rect 162360 3408 162366 3420
rect 208857 3417 208869 3420
rect 208903 3417 208915 3451
rect 208857 3411 208915 3417
rect 210329 3451 210387 3457
rect 210329 3417 210341 3451
rect 210375 3448 210387 3451
rect 211157 3451 211215 3457
rect 211157 3448 211169 3451
rect 210375 3420 211169 3448
rect 210375 3417 210387 3420
rect 210329 3411 210387 3417
rect 211157 3417 211169 3420
rect 211203 3417 211215 3451
rect 211157 3411 211215 3417
rect 219342 3408 219348 3460
rect 219400 3448 219406 3460
rect 246022 3448 246028 3460
rect 219400 3420 246028 3448
rect 219400 3408 219406 3420
rect 246022 3408 246028 3420
rect 246080 3408 246086 3460
rect 270494 3408 270500 3460
rect 270552 3448 270558 3460
rect 273346 3448 273352 3460
rect 270552 3420 273352 3448
rect 270552 3408 270558 3420
rect 273346 3408 273352 3420
rect 273404 3408 273410 3460
rect 285490 3408 285496 3460
rect 285548 3448 285554 3460
rect 294322 3448 294328 3460
rect 285548 3420 294328 3448
rect 285548 3408 285554 3420
rect 294322 3408 294328 3420
rect 294380 3408 294386 3460
rect 295242 3408 295248 3460
rect 295300 3448 295306 3460
rect 310974 3448 310980 3460
rect 295300 3420 310980 3448
rect 295300 3408 295306 3420
rect 310974 3408 310980 3420
rect 311032 3408 311038 3460
rect 313182 3408 313188 3460
rect 313240 3448 313246 3460
rect 346670 3448 346676 3460
rect 313240 3420 346676 3448
rect 313240 3408 313246 3420
rect 346670 3408 346676 3420
rect 346728 3408 346734 3460
rect 351822 3408 351828 3460
rect 351880 3448 351886 3460
rect 418264 3448 418292 3488
rect 421558 3476 421564 3488
rect 421616 3476 421622 3528
rect 422956 3516 422984 3556
rect 424318 3544 424324 3596
rect 424376 3584 424382 3596
rect 560754 3584 560760 3596
rect 424376 3556 560760 3584
rect 424376 3544 424382 3556
rect 560754 3544 560760 3556
rect 560812 3544 560818 3596
rect 439406 3516 439412 3528
rect 422956 3488 439412 3516
rect 439406 3476 439412 3488
rect 439464 3476 439470 3528
rect 442261 3519 442319 3525
rect 442261 3485 442273 3519
rect 442307 3516 442319 3519
rect 567838 3516 567844 3528
rect 442307 3488 567844 3516
rect 442307 3485 442319 3488
rect 442261 3479 442319 3485
rect 567838 3476 567844 3488
rect 567896 3476 567902 3528
rect 351880 3420 418292 3448
rect 351880 3408 351886 3420
rect 418338 3408 418344 3460
rect 418396 3448 418402 3460
rect 432322 3448 432328 3460
rect 418396 3420 432328 3448
rect 418396 3408 418402 3420
rect 432322 3408 432328 3420
rect 432380 3408 432386 3460
rect 432509 3451 432567 3457
rect 432509 3417 432521 3451
rect 432555 3448 432567 3451
rect 437385 3451 437443 3457
rect 437385 3448 437397 3451
rect 432555 3420 437397 3448
rect 432555 3417 432567 3420
rect 432509 3411 432567 3417
rect 437385 3417 437397 3420
rect 437431 3417 437443 3451
rect 437385 3411 437443 3417
rect 442166 3408 442172 3460
rect 442224 3448 442230 3460
rect 582190 3448 582196 3460
rect 442224 3420 582196 3448
rect 442224 3408 442230 3420
rect 582190 3408 582196 3420
rect 582248 3408 582254 3460
rect 189626 3340 189632 3392
rect 189684 3380 189690 3392
rect 190362 3380 190368 3392
rect 189684 3352 190368 3380
rect 189684 3340 189690 3352
rect 190362 3340 190368 3352
rect 190420 3340 190426 3392
rect 196713 3383 196771 3389
rect 196713 3349 196725 3383
rect 196759 3380 196771 3383
rect 197906 3380 197912 3392
rect 196759 3352 197912 3380
rect 196759 3349 196771 3352
rect 196713 3343 196771 3349
rect 197906 3340 197912 3352
rect 197964 3340 197970 3392
rect 207661 3383 207719 3389
rect 207661 3349 207673 3383
rect 207707 3380 207719 3383
rect 231854 3380 231860 3392
rect 207707 3352 231860 3380
rect 207707 3349 207719 3352
rect 207661 3343 207719 3349
rect 231854 3340 231860 3352
rect 231912 3340 231918 3392
rect 250346 3340 250352 3392
rect 250404 3380 250410 3392
rect 251082 3380 251088 3392
rect 250404 3352 251088 3380
rect 250404 3340 250410 3352
rect 251082 3340 251088 3352
rect 251140 3340 251146 3392
rect 293862 3340 293868 3392
rect 293920 3380 293926 3392
rect 308582 3380 308588 3392
rect 293920 3352 308588 3380
rect 293920 3340 293926 3352
rect 308582 3340 308588 3352
rect 308640 3340 308646 3392
rect 320082 3340 320088 3392
rect 320140 3380 320146 3392
rect 359734 3380 359740 3392
rect 320140 3352 359740 3380
rect 320140 3340 320146 3352
rect 359734 3340 359740 3352
rect 359792 3340 359798 3392
rect 389082 3340 389088 3392
rect 389140 3380 389146 3392
rect 492950 3380 492956 3392
rect 389140 3352 492956 3380
rect 389140 3340 389146 3352
rect 492950 3340 492956 3352
rect 493008 3340 493014 3392
rect 493318 3340 493324 3392
rect 493376 3380 493382 3392
rect 495989 3383 496047 3389
rect 495989 3380 496001 3383
rect 493376 3352 496001 3380
rect 493376 3340 493382 3352
rect 495989 3349 496001 3352
rect 496035 3349 496047 3383
rect 495989 3343 496047 3349
rect 496078 3340 496084 3392
rect 496136 3380 496142 3392
rect 504361 3383 504419 3389
rect 504361 3380 504373 3383
rect 496136 3352 504373 3380
rect 496136 3340 496142 3352
rect 504361 3349 504373 3352
rect 504407 3349 504419 3383
rect 504361 3343 504419 3349
rect 504453 3383 504511 3389
rect 504453 3349 504465 3383
rect 504499 3380 504511 3383
rect 510798 3380 510804 3392
rect 504499 3352 510804 3380
rect 504499 3349 504511 3352
rect 504453 3343 504511 3349
rect 510798 3340 510804 3352
rect 510856 3340 510862 3392
rect 511258 3340 511264 3392
rect 511316 3380 511322 3392
rect 513929 3383 513987 3389
rect 513929 3380 513941 3383
rect 511316 3352 513941 3380
rect 511316 3340 511322 3352
rect 513929 3349 513941 3352
rect 513975 3349 513987 3383
rect 513929 3343 513987 3349
rect 514021 3383 514079 3389
rect 514021 3349 514033 3383
rect 514067 3380 514079 3383
rect 564342 3380 564348 3392
rect 514067 3352 564348 3380
rect 514067 3349 514079 3352
rect 514021 3343 514079 3349
rect 564342 3340 564348 3352
rect 564400 3340 564406 3392
rect 175642 3312 175648 3324
rect 159376 3284 175648 3312
rect 147677 3275 147735 3281
rect 175642 3272 175648 3284
rect 175700 3272 175706 3324
rect 181070 3312 181076 3324
rect 177500 3284 181076 3312
rect 93302 3204 93308 3256
rect 93360 3244 93366 3256
rect 154577 3247 154635 3253
rect 154577 3244 154589 3247
rect 93360 3216 154589 3244
rect 93360 3204 93366 3216
rect 154577 3213 154589 3216
rect 154623 3213 154635 3247
rect 154577 3207 154635 3213
rect 164145 3247 164203 3253
rect 164145 3213 164157 3247
rect 164191 3244 164203 3247
rect 177500 3244 177528 3284
rect 181070 3272 181076 3284
rect 181128 3272 181134 3324
rect 197998 3272 198004 3324
rect 198056 3312 198062 3324
rect 204254 3312 204260 3324
rect 198056 3284 204260 3312
rect 198056 3272 198062 3284
rect 204254 3272 204260 3284
rect 204312 3272 204318 3324
rect 217042 3272 217048 3324
rect 217100 3312 217106 3324
rect 217100 3284 238064 3312
rect 217100 3272 217106 3284
rect 184934 3244 184940 3256
rect 164191 3216 177528 3244
rect 180812 3216 184940 3244
rect 164191 3213 164203 3216
rect 164145 3207 164203 3213
rect 76006 3176 76012 3188
rect 73172 3148 76012 3176
rect 57977 3139 58035 3145
rect 76006 3136 76012 3148
rect 76064 3136 76070 3188
rect 99282 3136 99288 3188
rect 99340 3176 99346 3188
rect 100018 3176 100024 3188
rect 99340 3148 100024 3176
rect 99340 3136 99346 3148
rect 100018 3136 100024 3148
rect 100076 3136 100082 3188
rect 100478 3136 100484 3188
rect 100536 3176 100542 3188
rect 180812 3176 180840 3216
rect 184934 3204 184940 3216
rect 184992 3204 184998 3256
rect 192018 3204 192024 3256
rect 192076 3244 192082 3256
rect 196621 3247 196679 3253
rect 196621 3244 196633 3247
rect 192076 3216 196633 3244
rect 192076 3204 192082 3216
rect 196621 3213 196633 3216
rect 196667 3213 196679 3247
rect 196621 3207 196679 3213
rect 199194 3204 199200 3256
rect 199252 3244 199258 3256
rect 199252 3216 200896 3244
rect 199252 3204 199258 3216
rect 100536 3148 180840 3176
rect 100536 3136 100542 3148
rect 181346 3136 181352 3188
rect 181404 3176 181410 3188
rect 195609 3179 195667 3185
rect 195609 3176 195621 3179
rect 181404 3148 195621 3176
rect 181404 3136 181410 3148
rect 195609 3145 195621 3148
rect 195655 3145 195667 3179
rect 200868 3176 200896 3216
rect 202690 3204 202696 3256
rect 202748 3244 202754 3256
rect 229738 3244 229744 3256
rect 202748 3216 229744 3244
rect 202748 3204 202754 3216
rect 229738 3204 229744 3216
rect 229796 3204 229802 3256
rect 238036 3244 238064 3284
rect 240778 3272 240784 3324
rect 240836 3312 240842 3324
rect 241422 3312 241428 3324
rect 240836 3284 241428 3312
rect 240836 3272 240842 3284
rect 241422 3272 241428 3284
rect 241480 3272 241486 3324
rect 253842 3272 253848 3324
rect 253900 3312 253906 3324
rect 257338 3312 257344 3324
rect 253900 3284 257344 3312
rect 253900 3272 253906 3284
rect 257338 3272 257344 3284
rect 257396 3272 257402 3324
rect 266998 3272 267004 3324
rect 267056 3312 267062 3324
rect 267642 3312 267648 3324
rect 267056 3284 267648 3312
rect 267056 3272 267062 3284
rect 267642 3272 267648 3284
rect 267700 3272 267706 3324
rect 292482 3272 292488 3324
rect 292540 3312 292546 3324
rect 306190 3312 306196 3324
rect 292540 3284 306196 3312
rect 292540 3272 292546 3284
rect 306190 3272 306196 3284
rect 306248 3272 306254 3324
rect 306282 3272 306288 3324
rect 306340 3312 306346 3324
rect 314562 3312 314568 3324
rect 306340 3284 314568 3312
rect 306340 3272 306346 3284
rect 314562 3272 314568 3284
rect 314620 3272 314626 3324
rect 317322 3272 317328 3324
rect 317380 3312 317386 3324
rect 353754 3312 353760 3324
rect 317380 3284 353760 3312
rect 317380 3272 317386 3284
rect 353754 3272 353760 3284
rect 353812 3272 353818 3324
rect 357802 3272 357808 3324
rect 357860 3312 357866 3324
rect 378778 3312 378784 3324
rect 357860 3284 378784 3312
rect 357860 3272 357866 3284
rect 378778 3272 378784 3284
rect 378836 3272 378842 3324
rect 383470 3272 383476 3324
rect 383528 3312 383534 3324
rect 482278 3312 482284 3324
rect 383528 3284 482284 3312
rect 383528 3272 383534 3284
rect 482278 3272 482284 3284
rect 482336 3272 482342 3324
rect 482373 3315 482431 3321
rect 482373 3281 482385 3315
rect 482419 3312 482431 3315
rect 485685 3315 485743 3321
rect 485685 3312 485697 3315
rect 482419 3284 485697 3312
rect 482419 3281 482431 3284
rect 482373 3275 482431 3281
rect 485685 3281 485697 3284
rect 485731 3281 485743 3315
rect 485685 3275 485743 3281
rect 486418 3272 486424 3324
rect 486476 3312 486482 3324
rect 489549 3315 489607 3321
rect 489549 3312 489561 3315
rect 486476 3284 489561 3312
rect 486476 3272 486482 3284
rect 489549 3281 489561 3284
rect 489595 3281 489607 3315
rect 489549 3275 489607 3281
rect 500218 3272 500224 3324
rect 500276 3312 500282 3324
rect 557166 3312 557172 3324
rect 500276 3284 557172 3312
rect 500276 3272 500282 3284
rect 557166 3272 557172 3284
rect 557224 3272 557230 3324
rect 243538 3244 243544 3256
rect 238036 3216 243544 3244
rect 243538 3204 243544 3216
rect 243596 3204 243602 3256
rect 261018 3204 261024 3256
rect 261076 3244 261082 3256
rect 262122 3244 262128 3256
rect 261076 3216 262128 3244
rect 261076 3204 261082 3216
rect 262122 3204 262128 3216
rect 262180 3204 262186 3256
rect 281442 3204 281448 3256
rect 281500 3244 281506 3256
rect 285950 3244 285956 3256
rect 281500 3216 285956 3244
rect 281500 3204 281506 3216
rect 285950 3204 285956 3216
rect 286008 3204 286014 3256
rect 294598 3204 294604 3256
rect 294656 3244 294662 3256
rect 301406 3244 301412 3256
rect 294656 3216 301412 3244
rect 294656 3204 294662 3216
rect 301406 3204 301412 3216
rect 301464 3204 301470 3256
rect 315850 3204 315856 3256
rect 315908 3244 315914 3256
rect 321646 3244 321652 3256
rect 315908 3216 321652 3244
rect 315908 3204 315914 3216
rect 321646 3204 321652 3216
rect 321704 3204 321710 3256
rect 322198 3204 322204 3256
rect 322256 3244 322262 3256
rect 357342 3244 357348 3256
rect 322256 3216 357348 3244
rect 322256 3204 322262 3216
rect 357342 3204 357348 3216
rect 357400 3204 357406 3256
rect 379422 3204 379428 3256
rect 379480 3244 379486 3256
rect 475102 3244 475108 3256
rect 379480 3216 475108 3244
rect 379480 3204 379486 3216
rect 475102 3204 475108 3216
rect 475160 3204 475166 3256
rect 496538 3244 496544 3256
rect 475212 3216 496544 3244
rect 225598 3176 225604 3188
rect 200868 3148 225604 3176
rect 195609 3139 195667 3145
rect 225598 3136 225604 3148
rect 225656 3136 225662 3188
rect 281350 3136 281356 3188
rect 281408 3176 281414 3188
rect 284754 3176 284760 3188
rect 281408 3148 284760 3176
rect 281408 3136 281414 3148
rect 284754 3136 284760 3148
rect 284812 3136 284818 3188
rect 297358 3136 297364 3188
rect 297416 3176 297422 3188
rect 300302 3176 300308 3188
rect 297416 3148 300308 3176
rect 297416 3136 297422 3148
rect 300302 3136 300308 3148
rect 300360 3136 300366 3188
rect 302878 3136 302884 3188
rect 302936 3176 302942 3188
rect 309778 3176 309784 3188
rect 302936 3148 309784 3176
rect 302936 3136 302942 3148
rect 309778 3136 309784 3148
rect 309836 3136 309842 3188
rect 320818 3136 320824 3188
rect 320876 3176 320882 3188
rect 350258 3176 350264 3188
rect 320876 3148 350264 3176
rect 320876 3136 320882 3148
rect 350258 3136 350264 3148
rect 350316 3136 350322 3188
rect 375282 3136 375288 3188
rect 375340 3176 375346 3188
rect 467926 3176 467932 3188
rect 375340 3148 467932 3176
rect 375340 3136 375346 3148
rect 467926 3136 467932 3148
rect 467984 3136 467990 3188
rect 473998 3136 474004 3188
rect 474056 3176 474062 3188
rect 475212 3176 475240 3216
rect 496538 3204 496544 3216
rect 496596 3204 496602 3256
rect 496633 3247 496691 3253
rect 496633 3213 496645 3247
rect 496679 3244 496691 3247
rect 546494 3244 546500 3256
rect 496679 3216 546500 3244
rect 496679 3213 496691 3216
rect 496633 3207 496691 3213
rect 546494 3204 546500 3216
rect 546552 3204 546558 3256
rect 474056 3148 475240 3176
rect 474056 3136 474062 3148
rect 478138 3136 478144 3188
rect 478196 3176 478202 3188
rect 485133 3179 485191 3185
rect 485133 3176 485145 3179
rect 478196 3148 485145 3176
rect 478196 3136 478202 3148
rect 485133 3145 485145 3148
rect 485179 3145 485191 3179
rect 485133 3139 485191 3145
rect 489825 3179 489883 3185
rect 489825 3145 489837 3179
rect 489871 3176 489883 3179
rect 503622 3176 503628 3188
rect 489871 3148 503628 3176
rect 489871 3145 489883 3148
rect 489825 3139 489883 3145
rect 503622 3136 503628 3148
rect 503680 3136 503686 3188
rect 504361 3179 504419 3185
rect 504361 3145 504373 3179
rect 504407 3176 504419 3179
rect 550082 3176 550088 3188
rect 504407 3148 550088 3176
rect 504407 3145 504419 3148
rect 504361 3139 504419 3145
rect 550082 3136 550088 3148
rect 550140 3136 550146 3188
rect 107562 3068 107568 3120
rect 107620 3108 107626 3120
rect 189258 3108 189264 3120
rect 107620 3080 189264 3108
rect 107620 3068 107626 3080
rect 189258 3068 189264 3080
rect 189316 3068 189322 3120
rect 206278 3068 206284 3120
rect 206336 3108 206342 3120
rect 231118 3108 231124 3120
rect 206336 3080 231124 3108
rect 206336 3068 206342 3080
rect 231118 3068 231124 3080
rect 231176 3068 231182 3120
rect 232498 3068 232504 3120
rect 232556 3108 232562 3120
rect 235350 3108 235356 3120
rect 232556 3080 235356 3108
rect 232556 3068 232562 3080
rect 235350 3068 235356 3080
rect 235408 3068 235414 3120
rect 258626 3068 258632 3120
rect 258684 3108 258690 3120
rect 259362 3108 259368 3120
rect 258684 3080 259368 3108
rect 258684 3068 258690 3080
rect 259362 3068 259368 3080
rect 259420 3068 259426 3120
rect 264606 3068 264612 3120
rect 264664 3108 264670 3120
rect 268378 3108 268384 3120
rect 264664 3080 268384 3108
rect 264664 3068 264670 3080
rect 268378 3068 268384 3080
rect 268436 3068 268442 3120
rect 372522 3068 372528 3120
rect 372580 3108 372586 3120
rect 460842 3108 460848 3120
rect 372580 3080 460848 3108
rect 372580 3068 372586 3080
rect 460842 3068 460848 3080
rect 460900 3068 460906 3120
rect 469858 3068 469864 3120
rect 469916 3108 469922 3120
rect 477865 3111 477923 3117
rect 477865 3108 477877 3111
rect 469916 3080 477877 3108
rect 469916 3068 469922 3080
rect 477865 3077 477877 3080
rect 477911 3077 477923 3111
rect 477865 3071 477923 3077
rect 478049 3111 478107 3117
rect 478049 3077 478061 3111
rect 478095 3108 478107 3111
rect 489362 3108 489368 3120
rect 478095 3080 489368 3108
rect 478095 3077 478107 3080
rect 478049 3071 478107 3077
rect 489362 3068 489368 3080
rect 489420 3068 489426 3120
rect 539318 3108 539324 3120
rect 489472 3080 539324 3108
rect 57977 3043 58035 3049
rect 57977 3009 57989 3043
rect 58023 3040 58035 3043
rect 62761 3043 62819 3049
rect 62761 3040 62773 3043
rect 58023 3012 62773 3040
rect 58023 3009 58035 3012
rect 57977 3003 58035 3009
rect 62761 3009 62773 3012
rect 62807 3009 62819 3043
rect 62761 3003 62819 3009
rect 103517 3043 103575 3049
rect 103517 3009 103529 3043
rect 103563 3040 103575 3043
rect 110601 3043 110659 3049
rect 110601 3040 110613 3043
rect 103563 3012 110613 3040
rect 103563 3009 103575 3012
rect 103517 3003 103575 3009
rect 110601 3009 110613 3012
rect 110647 3009 110659 3043
rect 110601 3003 110659 3009
rect 114738 3000 114744 3052
rect 114796 3040 114802 3052
rect 191834 3040 191840 3052
rect 114796 3012 191840 3040
rect 114796 3000 114802 3012
rect 191834 3000 191840 3012
rect 191892 3000 191898 3052
rect 193214 3000 193220 3052
rect 193272 3040 193278 3052
rect 194502 3040 194508 3052
rect 193272 3012 194508 3040
rect 193272 3000 193278 3012
rect 194502 3000 194508 3012
rect 194560 3000 194566 3052
rect 202785 3043 202843 3049
rect 202785 3009 202797 3043
rect 202831 3040 202843 3043
rect 202874 3040 202880 3052
rect 202831 3012 202880 3040
rect 202831 3009 202843 3012
rect 202785 3003 202843 3009
rect 202874 3000 202880 3012
rect 202932 3000 202938 3052
rect 204441 3043 204499 3049
rect 204441 3009 204453 3043
rect 204487 3040 204499 3043
rect 207661 3043 207719 3049
rect 207661 3040 207673 3043
rect 204487 3012 207673 3040
rect 204487 3009 204499 3012
rect 204441 3003 204499 3009
rect 207661 3009 207673 3012
rect 207707 3009 207719 3043
rect 207661 3003 207719 3009
rect 211062 3000 211068 3052
rect 211120 3040 211126 3052
rect 217318 3040 217324 3052
rect 211120 3012 217324 3040
rect 211120 3000 211126 3012
rect 217318 3000 217324 3012
rect 217376 3000 217382 3052
rect 220538 3000 220544 3052
rect 220596 3040 220602 3052
rect 232406 3040 232412 3052
rect 220596 3012 232412 3040
rect 220596 3000 220602 3012
rect 232406 3000 232412 3012
rect 232464 3000 232470 3052
rect 252646 3000 252652 3052
rect 252704 3040 252710 3052
rect 254578 3040 254584 3052
rect 252704 3012 254584 3040
rect 252704 3000 252710 3012
rect 254578 3000 254584 3012
rect 254636 3000 254642 3052
rect 377398 3000 377404 3052
rect 377456 3040 377462 3052
rect 453666 3040 453672 3052
rect 377456 3012 453672 3040
rect 377456 3000 377462 3012
rect 453666 3000 453672 3012
rect 453724 3000 453730 3052
rect 475378 3000 475384 3052
rect 475436 3040 475442 3052
rect 489089 3043 489147 3049
rect 489089 3040 489101 3043
rect 475436 3012 489101 3040
rect 475436 3000 475442 3012
rect 489089 3009 489101 3012
rect 489135 3009 489147 3043
rect 489089 3003 489147 3009
rect 489178 3000 489184 3052
rect 489236 3040 489242 3052
rect 489472 3040 489500 3080
rect 539318 3068 539324 3080
rect 539376 3068 539382 3120
rect 489236 3012 489500 3040
rect 489549 3043 489607 3049
rect 489236 3000 489242 3012
rect 489549 3009 489561 3043
rect 489595 3040 489607 3043
rect 532234 3040 532240 3052
rect 489595 3012 532240 3040
rect 489595 3009 489607 3012
rect 489549 3003 489607 3009
rect 532234 3000 532240 3012
rect 532292 3000 532298 3052
rect 124214 2932 124220 2984
rect 124272 2972 124278 2984
rect 125502 2972 125508 2984
rect 124272 2944 125508 2972
rect 124272 2932 124278 2944
rect 125502 2932 125508 2944
rect 125560 2932 125566 2984
rect 197354 2972 197360 2984
rect 125612 2944 197360 2972
rect 125410 2864 125416 2916
rect 125468 2904 125474 2916
rect 125612 2904 125640 2944
rect 197354 2932 197360 2944
rect 197412 2932 197418 2984
rect 203886 2932 203892 2984
rect 203944 2972 203950 2984
rect 210329 2975 210387 2981
rect 210329 2972 210341 2975
rect 203944 2944 210341 2972
rect 203944 2932 203950 2944
rect 210329 2941 210341 2944
rect 210375 2941 210387 2975
rect 210329 2935 210387 2941
rect 210421 2975 210479 2981
rect 210421 2941 210433 2975
rect 210467 2972 210479 2975
rect 220814 2972 220820 2984
rect 210467 2944 220820 2972
rect 210467 2941 210479 2944
rect 210421 2935 210479 2941
rect 220814 2932 220820 2944
rect 220872 2932 220878 2984
rect 221734 2932 221740 2984
rect 221792 2972 221798 2984
rect 228358 2972 228364 2984
rect 221792 2944 228364 2972
rect 221792 2932 221798 2944
rect 228358 2932 228364 2944
rect 228416 2932 228422 2984
rect 308398 2932 308404 2984
rect 308456 2972 308462 2984
rect 313366 2972 313372 2984
rect 308456 2944 313372 2972
rect 308456 2932 308462 2944
rect 313366 2932 313372 2944
rect 313424 2932 313430 2984
rect 376018 2932 376024 2984
rect 376076 2972 376082 2984
rect 414474 2972 414480 2984
rect 376076 2944 414480 2972
rect 376076 2932 376082 2944
rect 414474 2932 414480 2944
rect 414532 2932 414538 2984
rect 416038 2932 416044 2984
rect 416096 2972 416102 2984
rect 418154 2972 418160 2984
rect 416096 2944 418160 2972
rect 416096 2932 416102 2944
rect 418154 2932 418160 2944
rect 418212 2932 418218 2984
rect 418249 2975 418307 2981
rect 418249 2941 418261 2975
rect 418295 2972 418307 2975
rect 422297 2975 422355 2981
rect 422297 2972 422309 2975
rect 418295 2944 422309 2972
rect 418295 2941 418307 2944
rect 418249 2935 418307 2941
rect 422297 2941 422309 2944
rect 422343 2941 422355 2975
rect 422297 2935 422355 2941
rect 437385 2975 437443 2981
rect 437385 2941 437397 2975
rect 437431 2972 437443 2975
rect 482281 2975 482339 2981
rect 482281 2972 482293 2975
rect 437431 2944 456840 2972
rect 437431 2941 437443 2944
rect 437385 2935 437443 2941
rect 125468 2876 125640 2904
rect 125468 2864 125474 2876
rect 150434 2864 150440 2916
rect 150492 2904 150498 2916
rect 192478 2904 192484 2916
rect 150492 2876 192484 2904
rect 150492 2864 150498 2876
rect 192478 2864 192484 2876
rect 192536 2864 192542 2916
rect 195609 2907 195667 2913
rect 195609 2873 195621 2907
rect 195655 2904 195667 2907
rect 208857 2907 208915 2913
rect 195655 2876 208808 2904
rect 195655 2873 195667 2876
rect 195609 2867 195667 2873
rect 92106 2796 92112 2848
rect 92164 2836 92170 2848
rect 92382 2836 92388 2848
rect 92164 2808 92388 2836
rect 92164 2796 92170 2808
rect 92382 2796 92388 2808
rect 92440 2796 92446 2848
rect 122837 2839 122895 2845
rect 122837 2805 122849 2839
rect 122883 2836 122895 2839
rect 137925 2839 137983 2845
rect 137925 2836 137937 2839
rect 122883 2808 137937 2836
rect 122883 2805 122895 2808
rect 122837 2799 122895 2805
rect 137925 2805 137937 2808
rect 137971 2805 137983 2839
rect 137925 2799 137983 2805
rect 146846 2796 146852 2848
rect 146904 2836 146910 2848
rect 185578 2836 185584 2848
rect 146904 2808 185584 2836
rect 146904 2796 146910 2808
rect 185578 2796 185584 2808
rect 185636 2796 185642 2848
rect 196621 2839 196679 2845
rect 196621 2805 196633 2839
rect 196667 2836 196679 2839
rect 204441 2839 204499 2845
rect 204441 2836 204453 2839
rect 196667 2808 204453 2836
rect 196667 2805 196679 2808
rect 196621 2799 196679 2805
rect 204441 2805 204453 2808
rect 204487 2805 204499 2839
rect 204441 2799 204499 2805
rect 205082 2796 205088 2848
rect 205140 2836 205146 2848
rect 208210 2836 208216 2848
rect 205140 2808 208216 2836
rect 205140 2796 205146 2808
rect 208210 2796 208216 2808
rect 208268 2796 208274 2848
rect 208780 2836 208808 2876
rect 208857 2873 208869 2907
rect 208903 2904 208915 2907
rect 216950 2904 216956 2916
rect 208903 2876 216956 2904
rect 208903 2873 208915 2876
rect 208857 2867 208915 2873
rect 216950 2864 216956 2876
rect 217008 2864 217014 2916
rect 217965 2907 218023 2913
rect 217965 2873 217977 2907
rect 218011 2904 218023 2907
rect 223758 2904 223764 2916
rect 218011 2876 223764 2904
rect 218011 2873 218023 2876
rect 217965 2867 218023 2873
rect 223758 2864 223764 2876
rect 223816 2864 223822 2916
rect 368934 2864 368940 2916
rect 368992 2904 368998 2916
rect 428734 2904 428740 2916
rect 368992 2876 428740 2904
rect 368992 2864 368998 2876
rect 428734 2864 428740 2876
rect 428792 2864 428798 2916
rect 429838 2864 429844 2916
rect 429896 2904 429902 2916
rect 442261 2907 442319 2913
rect 442261 2904 442273 2907
rect 429896 2876 442273 2904
rect 429896 2864 429902 2876
rect 442261 2873 442273 2876
rect 442307 2873 442319 2907
rect 456812 2904 456840 2944
rect 466472 2944 482293 2972
rect 466472 2904 466500 2944
rect 482281 2941 482293 2944
rect 482327 2941 482339 2975
rect 482281 2935 482339 2941
rect 482370 2932 482376 2984
rect 482428 2972 482434 2984
rect 485041 2975 485099 2981
rect 485041 2972 485053 2975
rect 482428 2944 485053 2972
rect 482428 2932 482434 2944
rect 485041 2941 485053 2944
rect 485087 2941 485099 2975
rect 485041 2935 485099 2941
rect 485133 2975 485191 2981
rect 485133 2941 485145 2975
rect 485179 2972 485191 2975
rect 504453 2975 504511 2981
rect 504453 2972 504465 2975
rect 485179 2944 504465 2972
rect 485179 2941 485191 2944
rect 485133 2935 485191 2941
rect 504453 2941 504465 2944
rect 504499 2941 504511 2975
rect 504453 2935 504511 2941
rect 456812 2876 466500 2904
rect 442261 2867 442319 2873
rect 480898 2864 480904 2916
rect 480956 2904 480962 2916
rect 484949 2907 485007 2913
rect 484949 2904 484961 2907
rect 480956 2876 484961 2904
rect 480956 2864 480962 2876
rect 484949 2873 484961 2876
rect 484995 2873 485007 2907
rect 484949 2867 485007 2873
rect 485685 2907 485743 2913
rect 485685 2873 485697 2907
rect 485731 2904 485743 2907
rect 485774 2904 485780 2916
rect 485731 2876 485780 2904
rect 485731 2873 485743 2876
rect 485685 2867 485743 2873
rect 485774 2864 485780 2876
rect 485832 2864 485838 2916
rect 525058 2904 525064 2916
rect 485884 2876 525064 2904
rect 213178 2836 213184 2848
rect 208780 2808 213184 2836
rect 213178 2796 213184 2808
rect 213236 2796 213242 2848
rect 340782 2796 340788 2848
rect 340840 2836 340846 2848
rect 400214 2836 400220 2848
rect 340840 2808 400220 2836
rect 340840 2796 340846 2808
rect 400214 2796 400220 2808
rect 400272 2796 400278 2848
rect 402238 2796 402244 2848
rect 402296 2836 402302 2848
rect 446582 2836 446588 2848
rect 402296 2808 446588 2836
rect 402296 2796 402302 2808
rect 446582 2796 446588 2808
rect 446640 2796 446646 2848
rect 485041 2839 485099 2845
rect 485041 2805 485053 2839
rect 485087 2836 485099 2839
rect 485884 2836 485912 2876
rect 525058 2864 525064 2876
rect 525116 2864 525122 2916
rect 517882 2836 517888 2848
rect 485087 2808 485912 2836
rect 485976 2808 517888 2836
rect 485087 2805 485099 2808
rect 485041 2799 485099 2805
rect 422297 2771 422355 2777
rect 422297 2737 422309 2771
rect 422343 2768 422355 2771
rect 432509 2771 432567 2777
rect 432509 2768 432521 2771
rect 422343 2740 432521 2768
rect 422343 2737 422355 2740
rect 422297 2731 422355 2737
rect 432509 2737 432521 2740
rect 432555 2737 432567 2771
rect 432509 2731 432567 2737
rect 484949 2771 485007 2777
rect 484949 2737 484961 2771
rect 484995 2768 485007 2771
rect 485976 2768 486004 2808
rect 517882 2796 517888 2808
rect 517940 2796 517946 2848
rect 484995 2740 486004 2768
rect 484995 2737 485007 2740
rect 484949 2731 485007 2737
rect 194410 1300 194416 1352
rect 194468 1340 194474 1352
rect 202785 1343 202843 1349
rect 202785 1340 202797 1343
rect 194468 1312 202797 1340
rect 194468 1300 194474 1312
rect 202785 1309 202797 1312
rect 202831 1309 202843 1343
rect 202785 1303 202843 1309
rect 23106 552 23112 604
rect 23164 592 23170 604
rect 23382 592 23388 604
rect 23164 564 23388 592
rect 23164 552 23170 564
rect 23382 552 23388 564
rect 23440 552 23446 604
rect 67174 592 67180 604
rect 67135 564 67180 592
rect 67174 552 67180 564
rect 67232 552 67238 604
rect 178954 552 178960 604
rect 179012 592 179018 604
rect 179322 592 179328 604
rect 179012 564 179328 592
rect 179012 552 179018 564
rect 179322 552 179328 564
rect 179380 552 179386 604
rect 230106 552 230112 604
rect 230164 592 230170 604
rect 230382 592 230388 604
rect 230164 564 230388 592
rect 230164 552 230170 564
rect 230382 552 230388 564
rect 230440 552 230446 604
rect 238386 552 238392 604
rect 238444 592 238450 604
rect 238662 592 238668 604
rect 238444 564 238668 592
rect 238444 552 238450 564
rect 238662 552 238668 564
rect 238720 552 238726 604
rect 272886 552 272892 604
rect 272944 592 272950 604
rect 273162 592 273168 604
rect 272944 564 273168 592
rect 272944 552 272950 564
rect 273162 552 273168 564
rect 273220 552 273226 604
rect 290090 552 290096 604
rect 290148 592 290154 604
rect 290734 592 290740 604
rect 290148 564 290740 592
rect 290148 552 290154 564
rect 290734 552 290740 564
rect 290792 552 290798 604
rect 291378 552 291384 604
rect 291436 592 291442 604
rect 291930 592 291936 604
rect 291436 564 291936 592
rect 291436 552 291442 564
rect 291930 552 291936 564
rect 291988 552 291994 604
rect 318978 552 318984 604
rect 319036 592 319042 604
rect 319254 592 319260 604
rect 319036 564 319260 592
rect 319036 552 319042 564
rect 319254 552 319260 564
rect 319312 552 319318 604
rect 326430 592 326436 604
rect 326391 564 326436 592
rect 326430 552 326436 564
rect 326488 552 326494 604
rect 332870 552 332876 604
rect 332928 592 332934 604
rect 333606 592 333612 604
rect 332928 564 333612 592
rect 332928 552 332934 564
rect 333606 552 333612 564
rect 333664 552 333670 604
rect 336918 552 336924 604
rect 336976 592 336982 604
rect 337102 592 337108 604
rect 336976 564 337108 592
rect 336976 552 336982 564
rect 337102 552 337108 564
rect 337160 552 337166 604
rect 343910 552 343916 604
rect 343968 592 343974 604
rect 344278 592 344284 604
rect 343968 564 344284 592
rect 343968 552 343974 564
rect 344278 552 344284 564
rect 344336 552 344342 604
rect 456794 552 456800 604
rect 456852 592 456858 604
rect 457254 592 457260 604
rect 456852 564 457260 592
rect 456852 552 456858 564
rect 457254 552 457260 564
rect 457312 552 457318 604
rect 470594 552 470600 604
rect 470652 592 470658 604
rect 471514 592 471520 604
rect 470652 564 471520 592
rect 470652 552 470658 564
rect 471514 552 471520 564
rect 471572 552 471578 604
rect 473354 552 473360 604
rect 473412 592 473418 604
rect 473906 592 473912 604
rect 473412 564 473912 592
rect 473412 552 473418 564
rect 473906 552 473912 564
rect 473964 552 473970 604
<< via1 >>
rect 133880 700952 133932 701004
rect 267648 700952 267700 701004
rect 133788 700884 133840 700936
rect 283840 700884 283892 700936
rect 300124 700884 300176 700936
rect 434076 700884 434128 700936
rect 132500 700816 132552 700868
rect 332508 700816 332560 700868
rect 133696 700748 133748 700800
rect 218980 700748 219032 700800
rect 235172 700748 235224 700800
rect 434168 700748 434220 700800
rect 131120 700680 131172 700732
rect 348792 700680 348844 700732
rect 364984 700680 365036 700732
rect 433984 700680 434036 700732
rect 170312 700612 170364 700664
rect 434352 700612 434404 700664
rect 131212 700544 131264 700596
rect 397460 700544 397512 700596
rect 132316 700476 132368 700528
rect 413652 700476 413704 700528
rect 105452 700408 105504 700460
rect 434444 700408 434496 700460
rect 438124 700408 438176 700460
rect 494796 700408 494848 700460
rect 8116 700340 8168 700392
rect 13084 700340 13136 700392
rect 89168 700340 89220 700392
rect 126244 700340 126296 700392
rect 132592 700340 132644 700392
rect 462320 700340 462372 700392
rect 40500 700272 40552 700324
rect 434260 700272 434312 700324
rect 447784 700272 447836 700324
rect 559656 700272 559708 700324
rect 133420 700204 133472 700256
rect 202788 700204 202840 700256
rect 24308 699660 24360 699712
rect 24768 699660 24820 699712
rect 72424 699660 72476 699712
rect 72976 699660 73028 699712
rect 133328 699660 133380 699712
rect 137836 699660 137888 699712
rect 429844 699660 429896 699712
rect 433892 699660 433944 699712
rect 153568 698232 153620 698284
rect 154212 698232 154264 698284
rect 147588 697076 147640 697128
rect 154488 697076 154540 697128
rect 166908 697076 166960 697128
rect 173808 697076 173860 697128
rect 186228 697076 186280 697128
rect 193128 697076 193180 697128
rect 205548 697076 205600 697128
rect 212448 697076 212500 697128
rect 224868 697076 224920 697128
rect 231768 697076 231820 697128
rect 244188 697076 244240 697128
rect 251088 697076 251140 697128
rect 263508 697076 263560 697128
rect 270408 697076 270460 697128
rect 282828 697076 282880 697128
rect 289728 697076 289780 697128
rect 302148 697076 302200 697128
rect 309048 697076 309100 697128
rect 321468 697076 321520 697128
rect 328368 697076 328420 697128
rect 154580 686264 154632 686316
rect 159456 686264 159508 686316
rect 135260 686128 135312 686180
rect 142896 686128 142948 686180
rect 153292 685924 153344 685976
rect 153660 685924 153712 685976
rect 153292 684428 153344 684480
rect 3516 681708 3568 681760
rect 434720 681708 434772 681760
rect 446404 673480 446456 673532
rect 580172 673480 580224 673532
rect 3424 667904 3476 667956
rect 19984 667904 20036 667956
rect 153660 666544 153712 666596
rect 153476 656863 153528 656872
rect 153476 656829 153485 656863
rect 153485 656829 153519 656863
rect 153519 656829 153528 656863
rect 153476 656820 153528 656829
rect 154580 650360 154632 650412
rect 159456 650360 159508 650412
rect 135260 650224 135312 650276
rect 142896 650224 142948 650276
rect 153568 647232 153620 647284
rect 153568 645804 153620 645856
rect 153292 636259 153344 636268
rect 153292 636225 153301 636259
rect 153301 636225 153335 636259
rect 153335 636225 153344 636259
rect 153292 636216 153344 636225
rect 153292 630504 153344 630556
rect 153568 630504 153620 630556
rect 445024 626560 445076 626612
rect 580172 626560 580224 626612
rect 3424 623772 3476 623824
rect 434812 623772 434864 623824
rect 153568 621052 153620 621104
rect 153476 620916 153528 620968
rect 3424 609968 3476 610020
rect 21364 609968 21416 610020
rect 153292 598927 153344 598936
rect 153292 598893 153301 598927
rect 153301 598893 153335 598927
rect 153335 598893 153344 598927
rect 153292 598884 153344 598893
rect 4068 594804 4120 594856
rect 4896 594804 4948 594856
rect 154580 592424 154632 592476
rect 159456 592424 159508 592476
rect 135260 592288 135312 592340
rect 142896 592288 142948 592340
rect 153476 589296 153528 589348
rect 270408 583652 270460 583704
rect 307024 583652 307076 583704
rect 287704 583584 287756 583636
rect 319720 583584 319772 583636
rect 130384 583516 130436 583568
rect 311256 583516 311308 583568
rect 129004 583448 129056 583500
rect 330392 583448 330444 583500
rect 129280 583380 129332 583432
rect 347504 583380 347556 583432
rect 119344 583312 119396 583364
rect 336832 583312 336884 583364
rect 85396 583244 85448 583296
rect 334624 583244 334676 583296
rect 298468 583176 298520 583228
rect 332600 583176 332652 583228
rect 298376 583108 298428 583160
rect 341064 583108 341116 583160
rect 293868 583040 293920 583092
rect 338856 583040 338908 583092
rect 281448 582972 281500 583024
rect 326160 582972 326212 583024
rect 298284 582904 298336 582956
rect 353760 582904 353812 582956
rect 298560 582836 298612 582888
rect 355968 582836 356020 582888
rect 291108 582768 291160 582820
rect 351736 582768 351788 582820
rect 300492 582700 300544 582752
rect 362408 582700 362460 582752
rect 298192 582632 298244 582684
rect 345296 582632 345348 582684
rect 366640 582632 366692 582684
rect 378232 582632 378284 582684
rect 294604 582564 294656 582616
rect 313464 582564 313516 582616
rect 357992 582564 358044 582616
rect 378416 582564 378468 582616
rect 298652 582496 298704 582548
rect 321928 582496 321980 582548
rect 370872 582496 370924 582548
rect 378600 582496 378652 582548
rect 298744 582428 298796 582480
rect 328368 582428 328420 582480
rect 300400 582360 300452 582412
rect 309232 582360 309284 582412
rect 372896 582360 372948 582412
rect 378508 582360 378560 582412
rect 153384 579640 153436 579692
rect 153476 579640 153528 579692
rect 299388 579640 299440 579692
rect 304816 579640 304868 579692
rect 442264 579640 442316 579692
rect 580172 579640 580224 579692
rect 299480 579300 299532 579352
rect 300676 579300 300728 579352
rect 315212 579343 315264 579352
rect 315212 579309 315221 579343
rect 315221 579309 315255 579343
rect 315255 579309 315264 579343
rect 315212 579300 315264 579309
rect 317420 579343 317472 579352
rect 317420 579309 317429 579343
rect 317429 579309 317463 579343
rect 317463 579309 317472 579343
rect 317420 579300 317472 579309
rect 342996 579343 343048 579352
rect 342996 579309 343005 579343
rect 343005 579309 343039 579343
rect 343039 579309 343048 579343
rect 342996 579300 343048 579309
rect 364248 579343 364300 579352
rect 364248 579309 364257 579343
rect 364257 579309 364291 579343
rect 364291 579309 364300 579343
rect 364248 579300 364300 579309
rect 375380 579300 375432 579352
rect 378324 579300 378376 579352
rect 122748 578416 122800 578468
rect 115388 578348 115440 578400
rect 115204 578280 115256 578332
rect 129188 578212 129240 578264
rect 110328 575492 110380 575544
rect 298008 575492 298060 575544
rect 272524 569916 272576 569968
rect 298008 569916 298060 569968
rect 129648 563048 129700 563100
rect 296904 563048 296956 563100
rect 195888 561960 195940 562012
rect 197084 561892 197136 561944
rect 208676 561892 208728 561944
rect 217876 561892 217928 561944
rect 197268 561824 197320 561876
rect 214748 561824 214800 561876
rect 196992 561756 197044 561808
rect 202420 561756 202472 561808
rect 197176 561688 197228 561740
rect 205548 561688 205600 561740
rect 153292 560260 153344 560312
rect 153384 560260 153436 560312
rect 391204 556248 391256 556300
rect 484400 556248 484452 556300
rect 273168 556180 273220 556232
rect 297272 556180 297324 556232
rect 395344 556180 395396 556232
rect 511264 556180 511316 556232
rect 109408 554752 109460 554804
rect 110328 554752 110380 554804
rect 115940 554752 115992 554804
rect 92112 553936 92164 553988
rect 115296 553936 115348 553988
rect 89168 553868 89220 553920
rect 160744 553868 160796 553920
rect 115112 553800 115164 553852
rect 128360 553800 128412 553852
rect 129280 553800 129332 553852
rect 95056 553732 95108 553784
rect 120724 553732 120776 553784
rect 100760 553664 100812 553716
rect 129096 553664 129148 553716
rect 106464 553596 106516 553648
rect 140044 553596 140096 553648
rect 103704 553528 103756 553580
rect 146944 553528 146996 553580
rect 97816 553460 97868 553512
rect 153844 553460 153896 553512
rect 112352 553392 112404 553444
rect 116032 553392 116084 553444
rect 3148 552032 3200 552084
rect 28264 552032 28316 552084
rect 85488 549856 85540 549908
rect 86408 549856 86460 549908
rect 115388 549856 115440 549908
rect 118608 542376 118660 542428
rect 152464 542376 152516 542428
rect 286968 538228 287020 538280
rect 297640 538228 297692 538280
rect 117780 536800 117832 536852
rect 144184 536800 144236 536852
rect 296076 534012 296128 534064
rect 297456 534012 297508 534064
rect 117780 532720 117832 532772
rect 159364 532720 159416 532772
rect 514024 532720 514076 532772
rect 580172 532720 580224 532772
rect 153384 531292 153436 531344
rect 153476 531292 153528 531344
rect 117964 529864 118016 529916
rect 119344 529864 119396 529916
rect 118608 525036 118660 525088
rect 128728 525036 128780 525088
rect 128728 524764 128780 524816
rect 129188 524764 129240 524816
rect 70124 524424 70176 524476
rect 82820 524424 82872 524476
rect 153384 524424 153436 524476
rect 153476 524356 153528 524408
rect 280068 521636 280120 521688
rect 297180 521636 297232 521688
rect 128452 521568 128504 521620
rect 129004 521568 129056 521620
rect 295340 521568 295392 521620
rect 296076 521568 296128 521620
rect 85212 521228 85264 521280
rect 295340 521228 295392 521280
rect 199384 521160 199436 521212
rect 222384 521160 222436 521212
rect 199476 521092 199528 521144
rect 222568 521092 222620 521144
rect 198188 521024 198240 521076
rect 222660 521024 222712 521076
rect 117320 520956 117372 521008
rect 128452 520956 128504 521008
rect 198280 520956 198332 521008
rect 222476 520956 222528 521008
rect 85304 520888 85356 520940
rect 295984 520888 296036 520940
rect 298192 520888 298244 520940
rect 279424 518916 279476 518968
rect 297272 518916 297324 518968
rect 89352 518848 89404 518900
rect 130384 518848 130436 518900
rect 109592 518780 109644 518832
rect 113180 518780 113232 518832
rect 115204 518780 115256 518832
rect 86592 518712 86644 518764
rect 122748 518712 122800 518764
rect 127716 518780 127768 518832
rect 98000 518372 98052 518424
rect 126336 518372 126388 518424
rect 106648 518304 106700 518356
rect 151084 518304 151136 518356
rect 100944 518236 100996 518288
rect 157984 518236 158036 518288
rect 198096 518236 198148 518288
rect 218980 518236 219032 518288
rect 391296 518236 391348 518288
rect 479984 518236 480036 518288
rect 92296 518168 92348 518220
rect 126980 518168 127032 518220
rect 297456 518168 297508 518220
rect 398104 518168 398156 518220
rect 506848 518168 506900 518220
rect 205640 517488 205692 517540
rect 206652 517488 206704 517540
rect 284944 516128 284996 516180
rect 297824 516128 297876 516180
rect 153292 511980 153344 512032
rect 153568 511980 153620 512032
rect 294696 509260 294748 509312
rect 297732 509260 297784 509312
rect 192484 506472 192536 506524
rect 297732 506472 297784 506524
rect 153568 505180 153620 505232
rect 128636 505044 128688 505096
rect 128820 505044 128872 505096
rect 153384 505044 153436 505096
rect 96528 500896 96580 500948
rect 379520 500896 379572 500948
rect 103520 500828 103572 500880
rect 104808 500828 104860 500880
rect 379428 500828 379480 500880
rect 69848 500216 69900 500268
rect 95240 500216 95292 500268
rect 96528 500216 96580 500268
rect 118056 499468 118108 499520
rect 302884 499468 302936 499520
rect 300492 499128 300544 499180
rect 311900 499128 311952 499180
rect 298376 499060 298428 499112
rect 310612 499060 310664 499112
rect 324228 499060 324280 499112
rect 378416 499060 378468 499112
rect 298284 498992 298336 499044
rect 314752 498992 314804 499044
rect 321468 498992 321520 499044
rect 378324 498992 378376 499044
rect 298560 498924 298612 498976
rect 316040 498924 316092 498976
rect 317328 498924 317380 498976
rect 378232 498924 378284 498976
rect 298468 498856 298520 498908
rect 309140 498856 309192 498908
rect 310428 498856 310480 498908
rect 378600 498856 378652 498908
rect 298652 498788 298704 498840
rect 306472 498788 306524 498840
rect 309048 498788 309100 498840
rect 378508 498788 378560 498840
rect 300400 498584 300452 498636
rect 302240 498584 302292 498636
rect 132132 498176 132184 498228
rect 580172 498176 580224 498228
rect 129096 498108 129148 498160
rect 364248 498108 364300 498160
rect 116032 498040 116084 498092
rect 347320 498040 347372 498092
rect 120724 497972 120776 498024
rect 121368 497972 121420 498024
rect 338856 497972 338908 498024
rect 126336 497904 126388 497956
rect 334440 497904 334492 497956
rect 337476 497904 337528 497956
rect 370688 497904 370740 497956
rect 152464 497836 152516 497888
rect 153108 497836 153160 497888
rect 319720 497836 319772 497888
rect 320088 497836 320140 497888
rect 357992 497836 358044 497888
rect 289728 497768 289780 497820
rect 366456 497768 366508 497820
rect 284300 497700 284352 497752
rect 368480 497700 368532 497752
rect 111708 497632 111760 497684
rect 115296 497632 115348 497684
rect 291016 497632 291068 497684
rect 377128 497632 377180 497684
rect 108948 497564 109000 497616
rect 116032 497564 116084 497616
rect 284208 497564 284260 497616
rect 374920 497564 374972 497616
rect 83924 497496 83976 497548
rect 127072 497496 127124 497548
rect 360016 497496 360068 497548
rect 111800 497428 111852 497480
rect 125968 497428 126020 497480
rect 372712 497428 372764 497480
rect 285588 497360 285640 497412
rect 345112 497360 345164 497412
rect 292488 497292 292540 497344
rect 351552 497292 351604 497344
rect 301504 497224 301556 497276
rect 353576 497224 353628 497276
rect 295248 497156 295300 497208
rect 340880 497156 340932 497208
rect 277308 497088 277360 497140
rect 317512 497088 317564 497140
rect 319444 497088 319496 497140
rect 349344 497088 349396 497140
rect 288348 497020 288400 497072
rect 321744 497020 321796 497072
rect 334624 497020 334676 497072
rect 362224 497020 362276 497072
rect 279516 496952 279568 497004
rect 311072 496952 311124 497004
rect 333244 496952 333296 497004
rect 355784 496952 355836 497004
rect 304264 496884 304316 496936
rect 332416 496884 332468 496936
rect 126336 496816 126388 496868
rect 126888 496816 126940 496868
rect 285036 496816 285088 496868
rect 306840 496816 306892 496868
rect 308956 496816 309008 496868
rect 316684 496816 316736 496868
rect 322204 496816 322256 496868
rect 323952 496816 324004 496868
rect 330484 496816 330536 496868
rect 336648 496816 336700 496868
rect 337384 496816 337436 496868
rect 343088 496816 343140 496868
rect 3332 495456 3384 495508
rect 31024 495456 31076 495508
rect 153384 495388 153436 495440
rect 153568 495388 153620 495440
rect 153292 492600 153344 492652
rect 153568 492600 153620 492652
rect 128636 491240 128688 491292
rect 128728 491240 128780 491292
rect 284024 491283 284076 491292
rect 284024 491249 284033 491283
rect 284033 491249 284067 491283
rect 284067 491249 284076 491283
rect 284024 491240 284076 491249
rect 299756 485800 299808 485852
rect 300584 485800 300636 485852
rect 438216 485800 438268 485852
rect 580172 485800 580224 485852
rect 284116 485732 284168 485784
rect 125968 481584 126020 481636
rect 126060 481584 126112 481636
rect 284116 481584 284168 481636
rect 4068 480632 4120 480684
rect 4988 480632 5040 480684
rect 153292 476076 153344 476128
rect 153476 476076 153528 476128
rect 299572 476076 299624 476128
rect 299756 476076 299808 476128
rect 153384 473331 153436 473340
rect 153384 473297 153393 473331
rect 153393 473297 153427 473331
rect 153427 473297 153436 473331
rect 153384 473288 153436 473297
rect 299664 473331 299716 473340
rect 299664 473297 299673 473331
rect 299673 473297 299707 473331
rect 299707 473297 299716 473331
rect 299664 473288 299716 473297
rect 153384 466395 153436 466404
rect 153384 466361 153393 466395
rect 153393 466361 153427 466395
rect 153427 466361 153436 466395
rect 153384 466352 153436 466361
rect 299664 466395 299716 466404
rect 299664 466361 299673 466395
rect 299673 466361 299707 466395
rect 299707 466361 299716 466395
rect 299664 466352 299716 466361
rect 284116 463768 284168 463820
rect 283840 463632 283892 463684
rect 284116 463632 284168 463684
rect 133144 462340 133196 462392
rect 579804 462340 579856 462392
rect 125968 456832 126020 456884
rect 299572 456764 299624 456816
rect 299756 456764 299808 456816
rect 125968 456696 126020 456748
rect 125968 453976 126020 454028
rect 126060 453976 126112 454028
rect 284024 454019 284076 454028
rect 284024 453985 284033 454019
rect 284033 453985 284067 454019
rect 284067 453985 284076 454019
rect 284024 453976 284076 453985
rect 299664 454019 299716 454028
rect 299664 453985 299673 454019
rect 299673 453985 299707 454019
rect 299707 453985 299716 454019
rect 299664 453976 299716 453985
rect 126060 452591 126112 452600
rect 126060 452557 126069 452591
rect 126069 452557 126103 452591
rect 126103 452557 126112 452591
rect 126060 452548 126112 452557
rect 3056 451324 3108 451376
rect 267280 451324 267332 451376
rect 133236 451256 133288 451308
rect 580172 451256 580224 451308
rect 299664 447083 299716 447092
rect 299664 447049 299673 447083
rect 299673 447049 299707 447083
rect 299707 447049 299716 447083
rect 299664 447040 299716 447049
rect 284116 444456 284168 444508
rect 153384 444363 153436 444372
rect 153384 444329 153393 444363
rect 153393 444329 153427 444363
rect 153427 444329 153436 444363
rect 153384 444320 153436 444329
rect 283840 444320 283892 444372
rect 284116 444320 284168 444372
rect 126060 443819 126112 443828
rect 126060 443785 126069 443819
rect 126069 443785 126103 443819
rect 126103 443785 126112 443819
rect 126060 443776 126112 443785
rect 436744 438880 436796 438932
rect 580172 438880 580224 438932
rect 299572 437452 299624 437504
rect 299756 437452 299808 437504
rect 153384 437427 153436 437436
rect 153384 437393 153393 437427
rect 153393 437393 153427 437427
rect 153427 437393 153436 437427
rect 153384 437384 153436 437393
rect 125968 434664 126020 434716
rect 284024 434707 284076 434716
rect 284024 434673 284033 434707
rect 284033 434673 284067 434707
rect 284067 434673 284076 434707
rect 284024 434664 284076 434673
rect 299664 434707 299716 434716
rect 299664 434673 299673 434707
rect 299673 434673 299707 434707
rect 299707 434673 299716 434707
rect 299664 434664 299716 434673
rect 125876 427771 125928 427780
rect 125876 427737 125885 427771
rect 125885 427737 125919 427771
rect 125919 427737 125928 427771
rect 125876 427728 125928 427737
rect 299664 427771 299716 427780
rect 299664 427737 299673 427771
rect 299673 427737 299707 427771
rect 299707 427737 299716 427771
rect 299664 427728 299716 427737
rect 284116 425144 284168 425196
rect 125876 425008 125928 425060
rect 125968 425008 126020 425060
rect 283840 425008 283892 425060
rect 284116 425008 284168 425060
rect 4068 423648 4120 423700
rect 5080 423648 5132 423700
rect 153292 418208 153344 418260
rect 299572 418140 299624 418192
rect 299756 418140 299808 418192
rect 153200 418072 153252 418124
rect 133052 415420 133104 415472
rect 579804 415420 579856 415472
rect 126152 415352 126204 415404
rect 128636 415352 128688 415404
rect 153200 415352 153252 415404
rect 153476 415352 153528 415404
rect 284024 415395 284076 415404
rect 284024 415361 284033 415395
rect 284033 415361 284067 415395
rect 284067 415361 284076 415395
rect 284024 415352 284076 415361
rect 299664 415395 299716 415404
rect 299664 415361 299673 415395
rect 299673 415361 299707 415395
rect 299707 415361 299716 415395
rect 299664 415352 299716 415361
rect 251732 410796 251784 410848
rect 266360 410796 266412 410848
rect 246028 410728 246080 410780
rect 267832 410728 267884 410780
rect 228916 410660 228968 410712
rect 267004 410660 267056 410712
rect 223396 410592 223448 410644
rect 266728 410592 266780 410644
rect 211988 410524 212040 410576
rect 267096 410524 267148 410576
rect 206284 410456 206336 410508
rect 266452 410456 266504 410508
rect 248972 410388 249024 410440
rect 267740 410388 267792 410440
rect 243268 410320 243320 410372
rect 266544 410320 266596 410372
rect 240324 410252 240376 410304
rect 266636 410252 266688 410304
rect 237564 410184 237616 410236
rect 267372 410184 267424 410236
rect 196900 410116 196952 410168
rect 200580 410116 200632 410168
rect 234620 410116 234672 410168
rect 266820 410116 266872 410168
rect 199752 410048 199804 410100
rect 217692 410048 217744 410100
rect 257436 410048 257488 410100
rect 267464 410048 267516 410100
rect 199844 409980 199896 410032
rect 220452 409980 220504 410032
rect 254676 409980 254728 410032
rect 268844 409980 268896 410032
rect 199936 409912 199988 409964
rect 214748 409912 214800 409964
rect 260380 409912 260432 409964
rect 267556 409912 267608 409964
rect 200028 409844 200080 409896
rect 209044 409844 209096 409896
rect 265900 409844 265952 409896
rect 268936 409844 268988 409896
rect 199568 409640 199620 409692
rect 202880 409640 202932 409692
rect 199660 409572 199712 409624
rect 205640 409572 205692 409624
rect 196808 409504 196860 409556
rect 209780 409504 209832 409556
rect 195612 409436 195664 409488
rect 212540 409436 212592 409488
rect 195796 409368 195848 409420
rect 215300 409368 215352 409420
rect 196716 409300 196768 409352
rect 222752 409300 222804 409352
rect 196624 409232 196676 409284
rect 222844 409232 222896 409284
rect 195704 409164 195756 409216
rect 222200 409164 222252 409216
rect 195520 409096 195572 409148
rect 222292 409096 222344 409148
rect 188344 407804 188396 407856
rect 377404 407804 377456 407856
rect 70216 407736 70268 407788
rect 104808 407736 104860 407788
rect 393320 407736 393372 407788
rect 198004 407192 198056 407244
rect 386420 407192 386472 407244
rect 130384 407124 130436 407176
rect 358084 407124 358136 407176
rect 197728 406580 197780 406632
rect 295340 406580 295392 406632
rect 70308 406512 70360 406564
rect 295984 406512 296036 406564
rect 153108 406444 153160 406496
rect 393412 406444 393464 406496
rect 295984 406376 296036 406428
rect 344284 406376 344336 406428
rect 152464 405968 152516 406020
rect 153108 405968 153160 406020
rect 126060 405739 126112 405748
rect 126060 405705 126069 405739
rect 126069 405705 126103 405739
rect 126103 405705 126112 405739
rect 126060 405696 126112 405705
rect 128544 405739 128596 405748
rect 128544 405705 128553 405739
rect 128553 405705 128587 405739
rect 128587 405705 128596 405739
rect 128544 405696 128596 405705
rect 284024 405739 284076 405748
rect 284024 405705 284033 405739
rect 284033 405705 284067 405739
rect 284067 405705 284076 405739
rect 284024 405696 284076 405705
rect 295340 405696 295392 405748
rect 296076 405696 296128 405748
rect 299756 405696 299808 405748
rect 128544 405603 128596 405612
rect 128544 405569 128553 405603
rect 128553 405569 128587 405603
rect 128587 405569 128596 405603
rect 128544 405560 128596 405569
rect 386420 402908 386472 402960
rect 387248 402908 387300 402960
rect 120908 399304 120960 399356
rect 121368 399304 121420 399356
rect 125692 399304 125744 399356
rect 153384 398939 153436 398948
rect 153384 398905 153393 398939
rect 153393 398905 153427 398939
rect 153427 398905 153436 398939
rect 153384 398896 153436 398905
rect 71688 398828 71740 398880
rect 85488 398828 85540 398880
rect 85488 398692 85540 398744
rect 90272 398692 90324 398744
rect 128636 398692 128688 398744
rect 379520 398624 379572 398676
rect 380624 398624 380676 398676
rect 380440 398488 380492 398540
rect 380624 398488 380676 398540
rect 380164 398352 380216 398404
rect 380440 398352 380492 398404
rect 129464 398148 129516 398200
rect 152464 398148 152516 398200
rect 75828 398080 75880 398132
rect 115940 398080 115992 398132
rect 127256 398080 127308 398132
rect 134156 398080 134208 398132
rect 191104 398080 191156 398132
rect 80796 397876 80848 397928
rect 124864 397876 124916 397928
rect 100668 397808 100720 397860
rect 113180 397808 113232 397860
rect 114468 397808 114520 397860
rect 110972 397740 111024 397792
rect 111708 397740 111760 397792
rect 127164 397740 127216 397792
rect 106004 397672 106056 397724
rect 127624 397672 127676 397724
rect 95884 397604 95936 397656
rect 134156 397604 134208 397656
rect 85948 397536 86000 397588
rect 129464 397536 129516 397588
rect 115848 397468 115900 397520
rect 126336 397468 126388 397520
rect 124864 397400 124916 397452
rect 126152 397400 126204 397452
rect 380072 397332 380124 397384
rect 380256 397332 380308 397384
rect 69940 396788 69992 396840
rect 117964 396788 118016 396840
rect 126520 396788 126572 396840
rect 114468 396720 114520 396772
rect 128268 396720 128320 396772
rect 198004 396720 198056 396772
rect 153384 396083 153436 396092
rect 153384 396049 153393 396083
rect 153393 396049 153427 396083
rect 153427 396049 153436 396083
rect 153384 396040 153436 396049
rect 134156 395972 134208 396024
rect 299572 396015 299624 396024
rect 299572 395981 299581 396015
rect 299581 395981 299615 396015
rect 299615 395981 299624 396015
rect 299572 395972 299624 395981
rect 153384 395904 153436 395956
rect 84016 395836 84068 395888
rect 84108 395700 84160 395752
rect 70032 395632 70084 395684
rect 108948 395632 109000 395684
rect 125876 395632 125928 395684
rect 168656 395564 168708 395616
rect 179512 395496 179564 395548
rect 349068 395428 349120 395480
rect 361856 395428 361908 395480
rect 344284 395360 344336 395412
rect 380256 395360 380308 395412
rect 296076 395292 296128 395344
rect 364248 395292 364300 395344
rect 344928 395224 344980 395276
rect 384856 395224 384908 395276
rect 355968 395156 356020 395208
rect 389456 395156 389508 395208
rect 355876 395088 355928 395140
rect 375656 395088 375708 395140
rect 353208 395020 353260 395072
rect 378048 395020 378100 395072
rect 382648 394952 382700 395004
rect 347688 394884 347740 394936
rect 373448 394884 373500 394936
rect 284024 394816 284076 394868
rect 343548 394816 343600 394868
rect 371056 394816 371108 394868
rect 360016 394748 360068 394800
rect 368848 394748 368900 394800
rect 284024 394680 284076 394732
rect 360108 394680 360160 394732
rect 366456 394680 366508 394732
rect 125784 394340 125836 394392
rect 126152 394340 126204 394392
rect 315948 394068 316000 394120
rect 380624 394068 380676 394120
rect 307668 394000 307720 394052
rect 379428 394000 379480 394052
rect 271788 393932 271840 393984
rect 380440 393932 380492 393984
rect 379428 393456 379480 393508
rect 379704 393456 379756 393508
rect 380164 393388 380216 393440
rect 379704 393320 379756 393372
rect 284024 393295 284076 393304
rect 284024 393261 284033 393295
rect 284033 393261 284067 393295
rect 284067 393261 284076 393295
rect 284024 393252 284076 393261
rect 302148 393252 302200 393304
rect 380348 393252 380400 393304
rect 300768 393184 300820 393236
rect 379796 393184 379848 393236
rect 298652 393116 298704 393168
rect 380532 393116 380584 393168
rect 380072 393048 380124 393100
rect 295156 392980 295208 393032
rect 379520 392980 379572 393032
rect 292396 392912 292448 392964
rect 377496 392912 377548 392964
rect 292304 392844 292356 392896
rect 378140 392844 378192 392896
rect 379428 392887 379480 392896
rect 379428 392853 379437 392887
rect 379437 392853 379471 392887
rect 379471 392853 379480 392887
rect 379428 392844 379480 392853
rect 379612 392887 379664 392896
rect 379612 392853 379621 392887
rect 379621 392853 379655 392887
rect 379655 392853 379664 392887
rect 379612 392844 379664 392853
rect 286876 392776 286928 392828
rect 377036 392776 377088 392828
rect 377220 392819 377272 392828
rect 377220 392785 377229 392819
rect 377229 392785 377263 392819
rect 377263 392785 377272 392819
rect 377220 392776 377272 392785
rect 379704 392819 379756 392828
rect 379704 392785 379713 392819
rect 379713 392785 379747 392819
rect 379747 392785 379756 392819
rect 379704 392776 379756 392785
rect 379888 392776 379940 392828
rect 288256 392708 288308 392760
rect 379980 392708 380032 392760
rect 281356 392640 281408 392692
rect 277216 392572 277268 392624
rect 302056 392504 302108 392556
rect 380716 392751 380768 392760
rect 380716 392717 380725 392751
rect 380725 392717 380759 392751
rect 380759 392717 380768 392751
rect 380716 392708 380768 392717
rect 380808 392708 380860 392760
rect 300676 392436 300728 392488
rect 308956 392368 309008 392420
rect 314568 392300 314620 392352
rect 322848 392232 322900 392284
rect 302884 391212 302936 391264
rect 357440 391212 357492 391264
rect 416596 389376 416648 389428
rect 464252 389376 464304 389428
rect 418068 389308 418120 389360
rect 487436 389308 487488 389360
rect 401508 389240 401560 389292
rect 475844 389240 475896 389292
rect 416688 389172 416740 389224
rect 499028 389172 499080 389224
rect 153292 389147 153344 389156
rect 153292 389113 153301 389147
rect 153301 389113 153335 389147
rect 153335 389113 153344 389147
rect 153292 389104 153344 389113
rect 351828 387812 351880 387864
rect 357440 387812 357492 387864
rect 357348 386563 357400 386572
rect 357348 386529 357357 386563
rect 357357 386529 357391 386563
rect 357391 386529 357400 386563
rect 357348 386520 357400 386529
rect 128636 386384 128688 386436
rect 128912 386384 128964 386436
rect 133972 386427 134024 386436
rect 133972 386393 133981 386427
rect 133981 386393 134015 386427
rect 134015 386393 134024 386427
rect 133972 386384 134024 386393
rect 297456 386427 297508 386436
rect 297456 386393 297465 386427
rect 297465 386393 297499 386427
rect 297499 386393 297508 386427
rect 297456 386384 297508 386393
rect 299664 386384 299716 386436
rect 357348 386359 357400 386368
rect 357348 386325 357357 386359
rect 357357 386325 357391 386359
rect 357391 386325 357400 386359
rect 357348 386316 357400 386325
rect 133972 386291 134024 386300
rect 133972 386257 133981 386291
rect 133981 386257 134015 386291
rect 134015 386257 134024 386291
rect 133972 386248 134024 386257
rect 284116 383664 284168 383716
rect 297456 383503 297508 383512
rect 297456 383469 297465 383503
rect 297465 383469 297499 383503
rect 297499 383469 297508 383503
rect 297456 383460 297508 383469
rect 351184 380876 351236 380928
rect 357440 380876 357492 380928
rect 153292 379448 153344 379500
rect 153476 379448 153528 379500
rect 134156 376728 134208 376780
rect 357164 376728 357216 376780
rect 357256 376592 357308 376644
rect 297640 375368 297692 375420
rect 128820 375343 128872 375352
rect 128820 375309 128829 375343
rect 128829 375309 128863 375343
rect 128863 375309 128872 375343
rect 128820 375300 128872 375309
rect 333888 374008 333940 374060
rect 357440 374008 357492 374060
rect 413928 374008 413980 374060
rect 456800 374008 456852 374060
rect 297548 370515 297600 370524
rect 297548 370481 297557 370515
rect 297557 370481 297591 370515
rect 297591 370481 297600 370515
rect 297548 370472 297600 370481
rect 357348 367115 357400 367124
rect 357348 367081 357357 367115
rect 357357 367081 357391 367115
rect 357391 367081 357400 367115
rect 357348 367072 357400 367081
rect 153568 367047 153620 367056
rect 153568 367013 153577 367047
rect 153577 367013 153611 367047
rect 153611 367013 153620 367047
rect 153568 367004 153620 367013
rect 284116 367004 284168 367056
rect 390560 367004 390612 367056
rect 390744 366936 390796 366988
rect 2780 365712 2832 365764
rect 5172 365712 5224 365764
rect 128820 365755 128872 365764
rect 128820 365721 128829 365755
rect 128829 365721 128863 365755
rect 128863 365721 128872 365755
rect 128820 365712 128872 365721
rect 129372 365644 129424 365696
rect 197728 365644 197780 365696
rect 358544 364352 358596 364404
rect 358728 364352 358780 364404
rect 299664 362287 299716 362296
rect 299664 362253 299673 362287
rect 299673 362253 299707 362287
rect 299707 362253 299716 362287
rect 299664 362244 299716 362253
rect 360016 360136 360068 360188
rect 364524 360136 364576 360188
rect 360108 360068 360160 360120
rect 365720 360068 365772 360120
rect 126520 358708 126572 358760
rect 128912 358708 128964 358760
rect 360108 358640 360160 358692
rect 367376 358640 367428 358692
rect 359464 358572 359516 358624
rect 369584 358572 369636 358624
rect 363696 358504 363748 358556
rect 374184 358504 374236 358556
rect 362868 358436 362920 358488
rect 378784 358436 378836 358488
rect 362224 358368 362276 358420
rect 383384 358368 383436 358420
rect 354588 358300 354640 358352
rect 376576 358300 376628 358352
rect 350448 358232 350500 358284
rect 371976 358232 372028 358284
rect 342168 358164 342220 358216
rect 364984 358164 365036 358216
rect 361488 358096 361540 358148
rect 390376 358096 390428 358148
rect 333796 358028 333848 358080
rect 387984 358028 388036 358080
rect 297732 357688 297784 357740
rect 153660 357416 153712 357468
rect 284024 357459 284076 357468
rect 284024 357425 284033 357459
rect 284033 357425 284067 357459
rect 284067 357425 284076 357459
rect 284024 357416 284076 357425
rect 297640 357416 297692 357468
rect 297732 357416 297784 357468
rect 299756 357416 299808 357468
rect 362776 357416 362828 357468
rect 363604 357416 363656 357468
rect 412548 357416 412600 357468
rect 456800 357416 456852 357468
rect 134248 357391 134300 357400
rect 134248 357357 134257 357391
rect 134257 357357 134291 357391
rect 134291 357357 134300 357391
rect 134248 357348 134300 357357
rect 390744 357348 390796 357400
rect 390928 357348 390980 357400
rect 185584 355988 185636 356040
rect 188344 355988 188396 356040
rect 297640 355988 297692 356040
rect 390928 356031 390980 356040
rect 390928 355997 390937 356031
rect 390937 355997 390971 356031
rect 390971 355997 390980 356031
rect 390928 355988 390980 355997
rect 267280 355308 267332 355360
rect 436100 355308 436152 355360
rect 129004 350956 129056 351008
rect 130384 350956 130436 351008
rect 134248 347803 134300 347812
rect 134248 347769 134257 347803
rect 134257 347769 134291 347803
rect 134291 347769 134300 347803
rect 134248 347760 134300 347769
rect 153476 347760 153528 347812
rect 153568 347760 153620 347812
rect 128820 347735 128872 347744
rect 128820 347701 128829 347735
rect 128829 347701 128863 347735
rect 128863 347701 128872 347735
rect 128820 347692 128872 347701
rect 284116 347692 284168 347744
rect 297548 346443 297600 346452
rect 297548 346409 297557 346443
rect 297557 346409 297591 346443
rect 297591 346409 297600 346443
rect 297548 346400 297600 346409
rect 390928 346443 390980 346452
rect 390928 346409 390937 346443
rect 390937 346409 390971 346443
rect 390971 346409 390980 346443
rect 390928 346400 390980 346409
rect 358544 345040 358596 345092
rect 358728 345040 358780 345092
rect 504824 345040 504876 345092
rect 579988 345040 580040 345092
rect 132960 342864 133012 342916
rect 192484 342864 192536 342916
rect 199292 342864 199344 342916
rect 200212 342864 200264 342916
rect 128820 342456 128872 342508
rect 132960 342456 133012 342508
rect 503812 341980 503864 342032
rect 504180 341980 504232 342032
rect 131948 341640 132000 341692
rect 580632 341640 580684 341692
rect 132040 341572 132092 341624
rect 580816 341572 580868 341624
rect 131672 341504 131724 341556
rect 580724 341504 580776 341556
rect 390928 340892 390980 340944
rect 127164 340824 127216 340876
rect 385040 340824 385092 340876
rect 390836 340824 390888 340876
rect 127256 340756 127308 340808
rect 380900 340756 380952 340808
rect 503904 340756 503956 340808
rect 504732 340824 504784 340876
rect 126888 340688 126940 340740
rect 358176 340688 358228 340740
rect 128820 340620 128872 340672
rect 360200 340620 360252 340672
rect 127716 340552 127768 340604
rect 358084 340552 358136 340604
rect 128912 340484 128964 340536
rect 111708 340212 111760 340264
rect 127164 340212 127216 340264
rect 110328 340144 110380 340196
rect 127256 340144 127308 340196
rect 126060 340076 126112 340128
rect 126888 340076 126940 340128
rect 198096 338988 198148 339040
rect 209964 338988 210016 339040
rect 199476 338920 199528 338972
rect 214104 338920 214156 338972
rect 257712 338920 257764 338972
rect 267556 338920 267608 338972
rect 199384 338852 199436 338904
rect 215300 338852 215352 338904
rect 253664 338852 253716 338904
rect 268844 338852 268896 338904
rect 198188 338784 198240 338836
rect 220820 338784 220872 338836
rect 244188 338784 244240 338836
rect 267464 338784 267516 338836
rect 198280 338716 198332 338768
rect 222200 338716 222252 338768
rect 237288 338716 237340 338768
rect 267372 338716 267424 338768
rect 262128 338376 262180 338428
rect 268936 338376 268988 338428
rect 284024 338215 284076 338224
rect 284024 338181 284033 338215
rect 284033 338181 284067 338215
rect 284067 338181 284076 338215
rect 284024 338172 284076 338181
rect 153384 338104 153436 338156
rect 153568 338104 153620 338156
rect 107568 338036 107620 338088
rect 284024 338036 284076 338088
rect 302884 338036 302936 338088
rect 97908 337968 97960 338020
rect 126980 337968 127032 338020
rect 128912 338011 128964 338020
rect 128912 337977 128921 338011
rect 128921 337977 128955 338011
rect 128955 337977 128964 338011
rect 128912 337968 128964 337977
rect 231860 337968 231912 338020
rect 248696 337968 248748 338020
rect 87788 337900 87840 337952
rect 113088 337900 113140 337952
rect 127072 337900 127124 337952
rect 220452 337900 220504 337952
rect 238116 337900 238168 337952
rect 122748 337832 122800 337884
rect 127716 337832 127768 337884
rect 209044 337832 209096 337884
rect 220084 337832 220136 337884
rect 226156 337832 226208 337884
rect 248512 337832 248564 337884
rect 250996 337832 251048 337884
rect 260196 337832 260248 337884
rect 203340 337764 203392 337816
rect 215944 337764 215996 337816
rect 217508 337764 217560 337816
rect 241428 337764 241480 337816
rect 246028 337764 246080 337816
rect 253756 337764 253808 337816
rect 263140 337764 263192 337816
rect 200580 337696 200632 337748
rect 238024 337696 238076 337748
rect 240048 337696 240100 337748
rect 243084 337696 243136 337748
rect 247684 337696 247736 337748
rect 257436 337696 257488 337748
rect 117228 337628 117280 337680
rect 126428 337628 126480 337680
rect 214748 337628 214800 337680
rect 258724 337628 258776 337680
rect 206100 337560 206152 337612
rect 255320 337560 255372 337612
rect 401416 337560 401468 337612
rect 460572 337560 460624 337612
rect 117964 337492 118016 337544
rect 132684 337492 132736 337544
rect 297364 337492 297416 337544
rect 411168 337492 411220 337544
rect 472164 337492 472216 337544
rect 72884 337424 72936 337476
rect 103428 337424 103480 337476
rect 299756 337424 299808 337476
rect 408408 337424 408460 337476
rect 483756 337424 483808 337476
rect 77852 337356 77904 337408
rect 100668 337356 100720 337408
rect 329840 337356 329892 337408
rect 413836 337356 413888 337408
rect 495348 337356 495400 337408
rect 228916 337288 228968 337340
rect 232504 337288 232556 337340
rect 244924 337288 244976 337340
rect 237564 337220 237616 337272
rect 243084 337220 243136 337272
rect 234620 337084 234672 337136
rect 237748 337084 237800 337136
rect 251732 337084 251784 337136
rect 252468 337084 252520 337136
rect 92756 336812 92808 336864
rect 93768 336812 93820 336864
rect 102876 336812 102928 336864
rect 103336 336812 103388 336864
rect 223212 336812 223264 336864
rect 229744 336812 229796 336864
rect 244096 336812 244148 336864
rect 248788 336812 248840 336864
rect 254492 336812 254544 336864
rect 258264 336812 258316 336864
rect 2964 336744 3016 336796
rect 434904 336744 434956 336796
rect 82728 336676 82780 336728
rect 125968 336676 126020 336728
rect 257712 336676 257764 336728
rect 257804 336676 257856 336728
rect 390928 336719 390980 336728
rect 390928 336685 390937 336719
rect 390937 336685 390971 336719
rect 390971 336685 390980 336719
rect 390928 336676 390980 336685
rect 257804 335248 257856 335300
rect 503536 333276 503588 333328
rect 503812 333276 503864 333328
rect 504364 333276 504416 333328
rect 504824 333276 504876 333328
rect 129004 332324 129056 332376
rect 214012 331304 214064 331356
rect 128728 331279 128780 331288
rect 128728 331245 128737 331279
rect 128737 331245 128771 331279
rect 128771 331245 128780 331279
rect 128728 331236 128780 331245
rect 503628 331168 503680 331220
rect 503996 331168 504048 331220
rect 134248 331100 134300 331152
rect 134248 330964 134300 331016
rect 284116 328559 284168 328568
rect 284116 328525 284125 328559
rect 284125 328525 284159 328559
rect 284159 328525 284168 328559
rect 284116 328516 284168 328525
rect 128728 328491 128780 328500
rect 128728 328457 128737 328491
rect 128737 328457 128771 328491
rect 128771 328457 128780 328491
rect 128728 328448 128780 328457
rect 209780 328448 209832 328500
rect 209964 328448 210016 328500
rect 213920 328491 213972 328500
rect 213920 328457 213929 328491
rect 213929 328457 213963 328491
rect 213963 328457 213972 328491
rect 213920 328448 213972 328457
rect 284116 328380 284168 328432
rect 390928 327131 390980 327140
rect 390928 327097 390937 327131
rect 390937 327097 390971 327131
rect 390971 327097 390980 327131
rect 390928 327088 390980 327097
rect 358544 325660 358596 325712
rect 358728 325660 358780 325712
rect 297640 323663 297692 323672
rect 297640 323629 297649 323663
rect 297649 323629 297683 323663
rect 297683 323629 297692 323663
rect 297640 323620 297692 323629
rect 503904 321759 503956 321768
rect 503904 321725 503913 321759
rect 503913 321725 503947 321759
rect 503947 321725 503956 321759
rect 503904 321716 503956 321725
rect 390928 321648 390980 321700
rect 503996 321691 504048 321700
rect 503996 321657 504005 321691
rect 504005 321657 504039 321691
rect 504039 321657 504048 321691
rect 503996 321648 504048 321657
rect 132776 321580 132828 321632
rect 579620 321580 579672 321632
rect 390836 321555 390888 321564
rect 390836 321521 390845 321555
rect 390845 321521 390879 321555
rect 390879 321521 390888 321555
rect 390836 321512 390888 321521
rect 503904 321555 503956 321564
rect 503904 321521 503913 321555
rect 503913 321521 503947 321555
rect 503947 321521 503956 321555
rect 503904 321512 503956 321521
rect 297640 318903 297692 318912
rect 297640 318869 297649 318903
rect 297649 318869 297683 318903
rect 297683 318869 297692 318903
rect 297640 318860 297692 318869
rect 153384 318792 153436 318844
rect 153476 318792 153528 318844
rect 284024 318835 284076 318844
rect 284024 318801 284033 318835
rect 284033 318801 284067 318835
rect 284067 318801 284076 318835
rect 284024 318792 284076 318801
rect 503996 318835 504048 318844
rect 503996 318801 504005 318835
rect 504005 318801 504039 318835
rect 504039 318801 504048 318835
rect 503996 318792 504048 318801
rect 128636 318724 128688 318776
rect 128728 318724 128780 318776
rect 134248 318724 134300 318776
rect 209780 318767 209832 318776
rect 209780 318733 209789 318767
rect 209789 318733 209823 318767
rect 209823 318733 209832 318767
rect 209780 318724 209832 318733
rect 503720 318767 503772 318776
rect 503720 318733 503729 318767
rect 503729 318733 503763 318767
rect 503763 318733 503772 318767
rect 503720 318724 503772 318733
rect 257712 317475 257764 317484
rect 257712 317441 257721 317475
rect 257721 317441 257755 317475
rect 257755 317441 257764 317475
rect 257712 317432 257764 317441
rect 128636 317407 128688 317416
rect 128636 317373 128645 317407
rect 128645 317373 128679 317407
rect 128679 317373 128688 317407
rect 128636 317364 128688 317373
rect 153384 311924 153436 311976
rect 153476 311924 153528 311976
rect 297548 311924 297600 311976
rect 503628 311856 503680 311908
rect 503996 311856 504048 311908
rect 297640 311788 297692 311840
rect 503628 311720 503680 311772
rect 503996 311720 504048 311772
rect 131856 310496 131908 310548
rect 579712 310496 579764 310548
rect 283932 309204 283984 309256
rect 284116 309204 284168 309256
rect 128728 309136 128780 309188
rect 134156 309179 134208 309188
rect 134156 309145 134165 309179
rect 134165 309145 134199 309179
rect 134199 309145 134208 309179
rect 134156 309136 134208 309145
rect 209780 309179 209832 309188
rect 209780 309145 209789 309179
rect 209789 309145 209823 309179
rect 209823 309145 209832 309179
rect 209780 309136 209832 309145
rect 503812 309136 503864 309188
rect 284116 309068 284168 309120
rect 390928 309068 390980 309120
rect 504364 309111 504416 309120
rect 504364 309077 504373 309111
rect 504373 309077 504407 309111
rect 504407 309077 504416 309111
rect 504364 309068 504416 309077
rect 132684 308252 132736 308304
rect 132868 308252 132920 308304
rect 297824 308048 297876 308100
rect 4068 307776 4120 307828
rect 5264 307776 5316 307828
rect 297824 307776 297876 307828
rect 128728 307751 128780 307760
rect 128728 307717 128737 307751
rect 128737 307717 128771 307751
rect 128771 307717 128780 307751
rect 128728 307708 128780 307717
rect 257804 307751 257856 307760
rect 257804 307717 257813 307751
rect 257813 307717 257847 307751
rect 257847 307717 257856 307751
rect 257804 307708 257856 307717
rect 297640 307708 297692 307760
rect 358544 306348 358596 306400
rect 358728 306348 358780 306400
rect 153292 302200 153344 302252
rect 153476 302200 153528 302252
rect 128728 302175 128780 302184
rect 128728 302141 128737 302175
rect 128737 302141 128771 302175
rect 128771 302141 128780 302175
rect 128728 302132 128780 302141
rect 134156 302132 134208 302184
rect 134340 302132 134392 302184
rect 284024 299591 284076 299600
rect 284024 299557 284033 299591
rect 284033 299557 284067 299591
rect 284067 299557 284076 299591
rect 284024 299548 284076 299557
rect 390836 299523 390888 299532
rect 390836 299489 390845 299523
rect 390845 299489 390879 299523
rect 390879 299489 390888 299523
rect 390836 299480 390888 299489
rect 504456 299480 504508 299532
rect 209780 299455 209832 299464
rect 209780 299421 209789 299455
rect 209789 299421 209823 299455
rect 209823 299421 209832 299455
rect 209780 299412 209832 299421
rect 284024 299455 284076 299464
rect 284024 299421 284033 299455
rect 284033 299421 284067 299455
rect 284067 299421 284076 299455
rect 284024 299412 284076 299421
rect 257896 298120 257948 298172
rect 297548 298163 297600 298172
rect 297548 298129 297557 298163
rect 297557 298129 297591 298163
rect 297591 298129 297600 298163
rect 297548 298120 297600 298129
rect 128728 298095 128780 298104
rect 128728 298061 128737 298095
rect 128737 298061 128771 298095
rect 128771 298061 128780 298095
rect 128728 298052 128780 298061
rect 134340 298052 134392 298104
rect 3332 293972 3384 294024
rect 434536 293972 434588 294024
rect 504272 292544 504324 292596
rect 504456 292544 504508 292596
rect 128728 292451 128780 292460
rect 128728 292417 128737 292451
rect 128737 292417 128771 292451
rect 128771 292417 128780 292451
rect 128728 292408 128780 292417
rect 284116 289892 284168 289944
rect 209780 289867 209832 289876
rect 209780 289833 209789 289867
rect 209789 289833 209823 289867
rect 209823 289833 209832 289867
rect 209780 289824 209832 289833
rect 284116 289756 284168 289808
rect 390928 289756 390980 289808
rect 134248 288439 134300 288448
rect 134248 288405 134257 288439
rect 134257 288405 134291 288439
rect 134291 288405 134300 288439
rect 134248 288396 134300 288405
rect 257804 288396 257856 288448
rect 257896 288396 257948 288448
rect 504272 288439 504324 288448
rect 504272 288405 504281 288439
rect 504281 288405 504315 288439
rect 504315 288405 504324 288439
rect 504272 288396 504324 288405
rect 297640 288328 297692 288380
rect 257804 288303 257856 288312
rect 257804 288269 257813 288303
rect 257813 288269 257847 288303
rect 257847 288269 257856 288303
rect 257804 288260 257856 288269
rect 358544 287036 358596 287088
rect 358728 287036 358780 287088
rect 503720 283024 503772 283076
rect 503812 282956 503864 283008
rect 128636 282931 128688 282940
rect 128636 282897 128645 282931
rect 128645 282897 128679 282931
rect 128679 282897 128688 282931
rect 128636 282888 128688 282897
rect 153292 282888 153344 282940
rect 153476 282888 153528 282940
rect 284024 280279 284076 280288
rect 284024 280245 284033 280279
rect 284033 280245 284067 280279
rect 284067 280245 284076 280279
rect 284024 280236 284076 280245
rect 357256 280236 357308 280288
rect 357348 280236 357400 280288
rect 504456 280236 504508 280288
rect 390836 280211 390888 280220
rect 390836 280177 390845 280211
rect 390845 280177 390879 280211
rect 390879 280177 390888 280211
rect 390836 280168 390888 280177
rect 153384 280143 153436 280152
rect 153384 280109 153393 280143
rect 153393 280109 153427 280143
rect 153427 280109 153436 280143
rect 153384 280100 153436 280109
rect 209780 280143 209832 280152
rect 209780 280109 209789 280143
rect 209789 280109 209823 280143
rect 209823 280109 209832 280143
rect 209780 280100 209832 280109
rect 284024 280143 284076 280152
rect 284024 280109 284033 280143
rect 284033 280109 284067 280143
rect 284067 280109 284076 280143
rect 284024 280100 284076 280109
rect 357256 280143 357308 280152
rect 357256 280109 357265 280143
rect 357265 280109 357299 280143
rect 357299 280109 357308 280143
rect 357256 280100 357308 280109
rect 134156 278808 134208 278860
rect 134248 278808 134300 278860
rect 128636 278783 128688 278792
rect 128636 278749 128645 278783
rect 128645 278749 128679 278783
rect 128679 278749 128688 278783
rect 128636 278740 128688 278749
rect 257896 278740 257948 278792
rect 134248 278715 134300 278724
rect 134248 278681 134257 278715
rect 134257 278681 134291 278715
rect 134291 278681 134300 278715
rect 134248 278672 134300 278681
rect 504456 278715 504508 278724
rect 504456 278681 504465 278715
rect 504465 278681 504499 278715
rect 504499 278681 504508 278715
rect 504456 278672 504508 278681
rect 132684 274660 132736 274712
rect 579620 274660 579672 274712
rect 128636 273343 128688 273352
rect 128636 273309 128645 273343
rect 128645 273309 128679 273343
rect 128679 273309 128688 273343
rect 128636 273300 128688 273309
rect 503628 273300 503680 273352
rect 503996 273300 504048 273352
rect 153568 273232 153620 273284
rect 503628 273164 503680 273216
rect 503996 273164 504048 273216
rect 209780 270555 209832 270564
rect 209780 270521 209789 270555
rect 209789 270521 209823 270555
rect 209823 270521 209832 270555
rect 209780 270512 209832 270521
rect 284024 270555 284076 270564
rect 284024 270521 284033 270555
rect 284033 270521 284067 270555
rect 284067 270521 284076 270555
rect 284024 270512 284076 270521
rect 297640 270512 297692 270564
rect 357348 270512 357400 270564
rect 128636 270487 128688 270496
rect 128636 270453 128645 270487
rect 128645 270453 128679 270487
rect 128679 270453 128688 270487
rect 128636 270444 128688 270453
rect 153568 270487 153620 270496
rect 153568 270453 153577 270487
rect 153577 270453 153611 270487
rect 153611 270453 153620 270487
rect 153568 270444 153620 270453
rect 257804 270487 257856 270496
rect 257804 270453 257813 270487
rect 257813 270453 257847 270487
rect 257847 270453 257856 270487
rect 257804 270444 257856 270453
rect 390928 270487 390980 270496
rect 390928 270453 390937 270487
rect 390937 270453 390971 270487
rect 390971 270453 390980 270487
rect 390928 270444 390980 270453
rect 134248 269127 134300 269136
rect 134248 269093 134257 269127
rect 134257 269093 134291 269127
rect 134291 269093 134300 269127
rect 134248 269084 134300 269093
rect 504640 269084 504692 269136
rect 358544 267724 358596 267776
rect 358728 267724 358780 267776
rect 2780 264936 2832 264988
rect 5448 264936 5500 264988
rect 284024 263687 284076 263696
rect 284024 263653 284033 263687
rect 284033 263653 284067 263687
rect 284067 263653 284076 263687
rect 284024 263644 284076 263653
rect 297548 263687 297600 263696
rect 297548 263653 297557 263687
rect 297557 263653 297591 263687
rect 297591 263653 297600 263687
rect 297548 263644 297600 263653
rect 503720 263644 503772 263696
rect 503996 263644 504048 263696
rect 131580 263576 131632 263628
rect 580172 263576 580224 263628
rect 257804 263551 257856 263560
rect 257804 263517 257813 263551
rect 257813 263517 257847 263551
rect 257847 263517 257856 263551
rect 257804 263508 257856 263517
rect 503720 263508 503772 263560
rect 503996 263508 504048 263560
rect 390928 263483 390980 263492
rect 390928 263449 390937 263483
rect 390937 263449 390971 263483
rect 390971 263449 390980 263483
rect 390928 263440 390980 263449
rect 284024 260967 284076 260976
rect 284024 260933 284033 260967
rect 284033 260933 284067 260967
rect 284067 260933 284076 260967
rect 284024 260924 284076 260933
rect 153660 260856 153712 260908
rect 297548 260899 297600 260908
rect 297548 260865 297557 260899
rect 297557 260865 297591 260899
rect 297591 260865 297600 260899
rect 297548 260856 297600 260865
rect 134340 260788 134392 260840
rect 209780 260831 209832 260840
rect 209780 260797 209789 260831
rect 209789 260797 209823 260831
rect 209823 260797 209832 260831
rect 209780 260788 209832 260797
rect 257804 260831 257856 260840
rect 257804 260797 257813 260831
rect 257813 260797 257847 260831
rect 257847 260797 257856 260831
rect 257804 260788 257856 260797
rect 284024 260788 284076 260840
rect 284300 260788 284352 260840
rect 390928 260831 390980 260840
rect 390928 260797 390937 260831
rect 390937 260797 390971 260831
rect 390971 260797 390980 260831
rect 390928 260788 390980 260797
rect 504272 260831 504324 260840
rect 504272 260797 504281 260831
rect 504281 260797 504315 260831
rect 504315 260797 504324 260831
rect 504272 260788 504324 260797
rect 128728 259360 128780 259412
rect 284116 254600 284168 254652
rect 284300 254600 284352 254652
rect 153660 253988 153712 254040
rect 503628 253988 503680 254040
rect 503996 253988 504048 254040
rect 153568 253852 153620 253904
rect 503628 253852 503680 253904
rect 503996 253852 504048 253904
rect 257804 253827 257856 253836
rect 257804 253793 257813 253827
rect 257813 253793 257847 253827
rect 257847 253793 257856 253827
rect 257804 253784 257856 253793
rect 390928 253827 390980 253836
rect 390928 253793 390937 253827
rect 390937 253793 390971 253827
rect 390971 253793 390980 253827
rect 390928 253784 390980 253793
rect 504272 253827 504324 253836
rect 504272 253793 504281 253827
rect 504281 253793 504315 253827
rect 504315 253793 504324 253827
rect 504272 253784 504324 253793
rect 284208 251404 284260 251456
rect 209780 251311 209832 251320
rect 209780 251277 209789 251311
rect 209789 251277 209823 251311
rect 209823 251277 209832 251311
rect 209780 251268 209832 251277
rect 297364 251268 297416 251320
rect 297640 251268 297692 251320
rect 3332 251200 3384 251252
rect 284208 251200 284260 251252
rect 435088 251200 435140 251252
rect 257804 251132 257856 251184
rect 357164 251132 357216 251184
rect 357348 251132 357400 251184
rect 358452 251132 358504 251184
rect 358636 251132 358688 251184
rect 390928 251175 390980 251184
rect 390928 251141 390937 251175
rect 390937 251141 390971 251175
rect 390971 251141 390980 251175
rect 390928 251132 390980 251141
rect 504272 251175 504324 251184
rect 504272 251141 504281 251175
rect 504281 251141 504315 251175
rect 504315 251141 504324 251175
rect 504272 251132 504324 251141
rect 134248 250631 134300 250640
rect 134248 250597 134257 250631
rect 134257 250597 134291 250631
rect 134291 250597 134300 250631
rect 134248 250588 134300 250597
rect 503720 244400 503772 244452
rect 297640 244332 297692 244384
rect 503812 244332 503864 244384
rect 297640 244196 297692 244248
rect 128636 241587 128688 241596
rect 128636 241553 128645 241587
rect 128645 241553 128679 241587
rect 128679 241553 128688 241587
rect 128636 241544 128688 241553
rect 257712 241519 257764 241528
rect 257712 241485 257721 241519
rect 257721 241485 257755 241519
rect 257755 241485 257764 241519
rect 257712 241476 257764 241485
rect 391020 241476 391072 241528
rect 504456 241476 504508 241528
rect 134064 240116 134116 240168
rect 134340 240116 134392 240168
rect 134340 235288 134392 235340
rect 153292 234676 153344 234728
rect 503628 234676 503680 234728
rect 503996 234676 504048 234728
rect 128728 234608 128780 234660
rect 257712 234608 257764 234660
rect 128636 234540 128688 234592
rect 153292 234540 153344 234592
rect 504456 234676 504508 234728
rect 503628 234540 503680 234592
rect 503996 234540 504048 234592
rect 504364 234540 504416 234592
rect 257804 234472 257856 234524
rect 357164 234472 357216 234524
rect 357348 234472 357400 234524
rect 358452 234472 358504 234524
rect 358636 234472 358688 234524
rect 209780 231820 209832 231872
rect 209964 231820 210016 231872
rect 284116 231820 284168 231872
rect 284300 231820 284352 231872
rect 390836 231820 390888 231872
rect 391020 231820 391072 231872
rect 504364 231795 504416 231804
rect 504364 231761 504373 231795
rect 504373 231761 504407 231795
rect 504407 231761 504416 231795
rect 504364 231752 504416 231761
rect 297364 230460 297416 230512
rect 297456 230460 297508 230512
rect 131304 227740 131356 227792
rect 580172 227740 580224 227792
rect 390560 226992 390612 227044
rect 390836 226992 390888 227044
rect 503720 225088 503772 225140
rect 503812 225020 503864 225072
rect 153200 224995 153252 225004
rect 153200 224961 153209 224995
rect 153209 224961 153243 224995
rect 153243 224961 153252 224995
rect 153200 224952 153252 224961
rect 257712 224995 257764 225004
rect 257712 224961 257721 224995
rect 257721 224961 257755 224995
rect 257755 224961 257764 224995
rect 257712 224952 257764 224961
rect 2964 222164 3016 222216
rect 14464 222164 14516 222216
rect 134248 222207 134300 222216
rect 134248 222173 134257 222207
rect 134257 222173 134291 222207
rect 134291 222173 134300 222207
rect 134248 222164 134300 222173
rect 153200 222207 153252 222216
rect 153200 222173 153209 222207
rect 153209 222173 153243 222207
rect 153243 222173 153252 222207
rect 153200 222164 153252 222173
rect 257712 222207 257764 222216
rect 257712 222173 257721 222207
rect 257721 222173 257755 222207
rect 257755 222173 257764 222207
rect 257712 222164 257764 222173
rect 297364 222164 297416 222216
rect 297456 222164 297508 222216
rect 504456 222164 504508 222216
rect 364524 222139 364576 222148
rect 364524 222105 364533 222139
rect 364533 222105 364567 222139
rect 364567 222105 364576 222139
rect 364524 222096 364576 222105
rect 390560 219376 390612 219428
rect 390744 219376 390796 219428
rect 131488 216656 131540 216708
rect 579620 216656 579672 216708
rect 283932 215364 283984 215416
rect 503628 215364 503680 215416
rect 503996 215364 504048 215416
rect 153200 215296 153252 215348
rect 257712 215296 257764 215348
rect 153292 215160 153344 215212
rect 504456 215364 504508 215416
rect 283932 215228 283984 215280
rect 308864 215228 308916 215280
rect 309048 215228 309100 215280
rect 503628 215228 503680 215280
rect 503996 215228 504048 215280
rect 504272 215228 504324 215280
rect 257804 215160 257856 215212
rect 209780 212508 209832 212560
rect 209964 212508 210016 212560
rect 297364 212508 297416 212560
rect 297640 212508 297692 212560
rect 357164 212508 357216 212560
rect 357256 212508 357308 212560
rect 364708 212508 364760 212560
rect 153292 212483 153344 212492
rect 153292 212449 153301 212483
rect 153301 212449 153335 212483
rect 153335 212449 153344 212483
rect 153292 212440 153344 212449
rect 298560 210400 298612 210452
rect 299020 210400 299072 210452
rect 297548 210264 297600 210316
rect 298008 210264 298060 210316
rect 390560 209788 390612 209840
rect 390744 209788 390796 209840
rect 244004 209720 244056 209772
rect 244188 209720 244240 209772
rect 301872 208496 301924 208548
rect 302148 208496 302200 208548
rect 2964 207000 3016 207052
rect 435180 207000 435232 207052
rect 503720 205776 503772 205828
rect 503812 205708 503864 205760
rect 257712 205683 257764 205692
rect 257712 205649 257721 205683
rect 257721 205649 257755 205683
rect 257755 205649 257764 205683
rect 257712 205640 257764 205649
rect 503720 205640 503772 205692
rect 503996 205640 504048 205692
rect 504180 205683 504232 205692
rect 504180 205649 504189 205683
rect 504189 205649 504223 205683
rect 504223 205649 504232 205683
rect 504180 205640 504232 205649
rect 196716 205300 196768 205352
rect 226892 205300 226944 205352
rect 196624 205232 196676 205284
rect 227904 205232 227956 205284
rect 195888 205164 195940 205216
rect 228640 205164 228692 205216
rect 195612 205096 195664 205148
rect 229560 205096 229612 205148
rect 195796 205028 195848 205080
rect 230480 205028 230532 205080
rect 195520 204960 195572 205012
rect 231216 204960 231268 205012
rect 195704 204892 195756 204944
rect 233240 204892 233292 204944
rect 266360 204892 266412 204944
rect 267464 204892 267516 204944
rect 255780 204144 255832 204196
rect 268292 204144 268344 204196
rect 253572 204076 253624 204128
rect 269028 204076 269080 204128
rect 250536 204008 250588 204060
rect 268016 204008 268068 204060
rect 199016 203940 199068 203992
rect 238760 203940 238812 203992
rect 247592 203940 247644 203992
rect 268200 203940 268252 203992
rect 197728 203872 197780 203924
rect 257160 203872 257212 203924
rect 198004 203804 198056 203856
rect 260380 203804 260432 203856
rect 198464 203736 198516 203788
rect 262772 203736 262824 203788
rect 197452 203668 197504 203720
rect 262956 203668 263008 203720
rect 197820 203600 197872 203652
rect 265256 203600 265308 203652
rect 198372 203532 198424 203584
rect 267372 203532 267424 203584
rect 153384 202852 153436 202904
rect 257712 202895 257764 202904
rect 199936 202784 199988 202836
rect 239680 202784 239732 202836
rect 240140 202784 240192 202836
rect 196900 202716 196952 202768
rect 200028 202648 200080 202700
rect 239220 202716 239272 202768
rect 240048 202716 240100 202768
rect 257712 202861 257721 202895
rect 257721 202861 257755 202895
rect 257755 202861 257764 202895
rect 257712 202852 257764 202861
rect 283656 202852 283708 202904
rect 283748 202852 283800 202904
rect 297456 202852 297508 202904
rect 297640 202852 297692 202904
rect 504180 202895 504232 202904
rect 504180 202861 504189 202895
rect 504189 202861 504223 202895
rect 504223 202861 504232 202895
rect 504180 202852 504232 202861
rect 240508 202784 240560 202836
rect 241428 202784 241480 202836
rect 241520 202648 241572 202700
rect 242072 202716 242124 202768
rect 247684 202716 247736 202768
rect 251824 202716 251876 202768
rect 267924 202784 267976 202836
rect 270960 202784 271012 202836
rect 271788 202784 271840 202836
rect 272248 202784 272300 202836
rect 273168 202784 273220 202836
rect 273996 202784 274048 202836
rect 274548 202784 274600 202836
rect 277032 202784 277084 202836
rect 277308 202784 277360 202836
rect 278688 202784 278740 202836
rect 279424 202784 279476 202836
rect 280528 202784 280580 202836
rect 281356 202784 281408 202836
rect 298652 202784 298704 202836
rect 299112 202784 299164 202836
rect 300124 202784 300176 202836
rect 300768 202784 300820 202836
rect 301412 202784 301464 202836
rect 302056 202784 302108 202836
rect 309140 202784 309192 202836
rect 309600 202784 309652 202836
rect 311900 202784 311952 202836
rect 312544 202784 312596 202836
rect 313556 202784 313608 202836
rect 314568 202784 314620 202836
rect 314752 202784 314804 202836
rect 315580 202784 315632 202836
rect 316684 202784 316736 202836
rect 321652 202784 321704 202836
rect 341340 202784 341392 202836
rect 342168 202784 342220 202836
rect 258724 202716 258776 202768
rect 263876 202716 263928 202768
rect 266360 202716 266412 202768
rect 267188 202716 267240 202768
rect 271420 202716 271472 202768
rect 272524 202716 272576 202768
rect 279240 202716 279292 202768
rect 280068 202716 280120 202768
rect 282276 202716 282328 202768
rect 284944 202716 284996 202768
rect 297916 202716 297968 202768
rect 298836 202716 298888 202768
rect 299480 202716 299532 202768
rect 313648 202716 313700 202768
rect 318616 202716 318668 202768
rect 333244 202716 333296 202768
rect 245200 202648 245252 202700
rect 250904 202648 250956 202700
rect 268384 202648 268436 202700
rect 299204 202648 299256 202700
rect 304356 202648 304408 202700
rect 304908 202648 304960 202700
rect 309140 202648 309192 202700
rect 311164 202648 311216 202700
rect 330484 202648 330536 202700
rect 358728 202648 358780 202700
rect 363420 202784 363472 202836
rect 375748 202784 375800 202836
rect 391204 202784 391256 202836
rect 400588 202784 400640 202836
rect 401416 202784 401468 202836
rect 413192 202784 413244 202836
rect 413928 202784 413980 202836
rect 415768 202784 415820 202836
rect 416596 202784 416648 202836
rect 417516 202784 417568 202836
rect 418068 202784 418120 202836
rect 374460 202716 374512 202768
rect 391296 202716 391348 202768
rect 504180 202716 504232 202768
rect 504456 202716 504508 202768
rect 361396 202648 361448 202700
rect 362224 202648 362276 202700
rect 376484 202648 376536 202700
rect 398104 202648 398156 202700
rect 160744 202580 160796 202632
rect 169116 202580 169168 202632
rect 197636 202580 197688 202632
rect 157984 202512 158036 202564
rect 176936 202512 176988 202564
rect 197544 202512 197596 202564
rect 244648 202580 244700 202632
rect 268108 202580 268160 202632
rect 299388 202580 299440 202632
rect 320640 202580 320692 202632
rect 359648 202580 359700 202632
rect 360108 202580 360160 202632
rect 360568 202580 360620 202632
rect 361488 202580 361540 202632
rect 362316 202580 362368 202632
rect 362868 202580 362920 202632
rect 363604 202580 363656 202632
rect 364340 202580 364392 202632
rect 367008 202580 367060 202632
rect 395344 202580 395396 202632
rect 244740 202512 244792 202564
rect 247500 202512 247552 202564
rect 267832 202512 267884 202564
rect 298928 202512 298980 202564
rect 303068 202512 303120 202564
rect 303160 202512 303212 202564
rect 304264 202512 304316 202564
rect 306656 202512 306708 202564
rect 307668 202512 307720 202564
rect 325700 202512 325752 202564
rect 346676 202512 346728 202564
rect 351184 202512 351236 202564
rect 357900 202512 357952 202564
rect 393320 202512 393372 202564
rect 159364 202444 159416 202496
rect 178040 202444 178092 202496
rect 197360 202444 197412 202496
rect 251916 202444 251968 202496
rect 252468 202444 252520 202496
rect 268476 202444 268528 202496
rect 286232 202444 286284 202496
rect 286876 202444 286928 202496
rect 287520 202444 287572 202496
rect 288256 202444 288308 202496
rect 289452 202444 289504 202496
rect 289728 202444 289780 202496
rect 290556 202444 290608 202496
rect 291016 202444 291068 202496
rect 292212 202444 292264 202496
rect 292396 202444 292448 202496
rect 153844 202376 153896 202428
rect 182180 202376 182232 202428
rect 199200 202376 199252 202428
rect 254032 202376 254084 202428
rect 255964 202376 256016 202428
rect 268568 202376 268620 202428
rect 275284 202376 275336 202428
rect 285036 202376 285088 202428
rect 289268 202376 289320 202428
rect 298744 202444 298796 202496
rect 299296 202444 299348 202496
rect 325148 202444 325200 202496
rect 352748 202444 352800 202496
rect 353208 202444 353260 202496
rect 358728 202444 358780 202496
rect 359464 202444 359516 202496
rect 393504 202444 393556 202496
rect 298008 202376 298060 202428
rect 310612 202376 310664 202428
rect 311256 202376 311308 202428
rect 325700 202376 325752 202428
rect 333152 202376 333204 202428
rect 333888 202376 333940 202428
rect 348332 202376 348384 202428
rect 390652 202376 390704 202428
rect 400956 202376 401008 202428
rect 401508 202376 401560 202428
rect 140044 202308 140096 202360
rect 168380 202308 168432 202360
rect 199108 202308 199160 202360
rect 258448 202308 258500 202360
rect 151084 202240 151136 202292
rect 181260 202240 181312 202292
rect 198924 202240 198976 202292
rect 261944 202308 261996 202360
rect 265164 202308 265216 202360
rect 266912 202308 266964 202360
rect 280988 202308 281040 202360
rect 281448 202308 281500 202360
rect 282736 202308 282788 202360
rect 294604 202308 294656 202360
rect 298560 202308 298612 202360
rect 305000 202308 305052 202360
rect 334624 202308 334676 202360
rect 345756 202308 345808 202360
rect 392032 202308 392084 202360
rect 103336 202172 103388 202224
rect 142528 202172 142580 202224
rect 146944 202172 146996 202224
rect 180340 202172 180392 202224
rect 198832 202172 198884 202224
rect 266820 202240 266872 202292
rect 283564 202240 283616 202292
rect 337384 202240 337436 202292
rect 344008 202240 344060 202292
rect 390560 202240 390612 202292
rect 414940 202240 414992 202292
rect 503904 202240 503956 202292
rect 260196 202172 260248 202224
rect 275744 202172 275796 202224
rect 287704 202172 287756 202224
rect 288808 202172 288860 202224
rect 322204 202172 322256 202224
rect 332508 202172 332560 202224
rect 391940 202172 391992 202224
rect 411076 202172 411128 202224
rect 503812 202172 503864 202224
rect 93768 202104 93820 202156
rect 134708 202104 134760 202156
rect 144184 202104 144236 202156
rect 178684 202104 178736 202156
rect 197912 202104 197964 202156
rect 269488 202104 269540 202156
rect 271696 202104 271748 202156
rect 337476 202104 337528 202156
rect 342076 202104 342128 202156
rect 393412 202104 393464 202156
rect 409236 202104 409288 202156
rect 503720 202104 503772 202156
rect 200028 202036 200080 202088
rect 236644 202036 236696 202088
rect 237288 202036 237340 202088
rect 240968 202036 241020 202088
rect 267280 202036 267332 202088
rect 299020 202036 299072 202088
rect 311992 202036 312044 202088
rect 315304 202036 315356 202088
rect 319444 202036 319496 202088
rect 351736 202036 351788 202088
rect 362868 202036 362920 202088
rect 363696 202036 363748 202088
rect 199936 201968 199988 202020
rect 198648 201900 198700 201952
rect 198740 201832 198792 201884
rect 211712 201832 211764 201884
rect 232504 201968 232556 202020
rect 236736 201968 236788 202020
rect 238116 201968 238168 202020
rect 258356 201968 258408 202020
rect 216036 201900 216088 201952
rect 215944 201832 215996 201884
rect 247776 201900 247828 201952
rect 251456 201900 251508 201952
rect 268660 201968 268712 202020
rect 291384 201968 291436 202020
rect 292488 201968 292540 202020
rect 296168 201968 296220 202020
rect 301504 201968 301556 202020
rect 315396 201968 315448 202020
rect 242164 201832 242216 201884
rect 248972 201832 249024 201884
rect 266544 201900 266596 201952
rect 298376 201900 298428 201952
rect 196808 201764 196860 201816
rect 199292 201696 199344 201748
rect 219532 201696 219584 201748
rect 220820 201764 220872 201816
rect 221280 201764 221332 201816
rect 229744 201764 229796 201816
rect 237380 201764 237432 201816
rect 238024 201764 238076 201816
rect 223028 201696 223080 201748
rect 199568 201628 199620 201680
rect 218612 201628 218664 201680
rect 241060 201628 241112 201680
rect 242992 201696 243044 201748
rect 244096 201696 244148 201748
rect 244924 201696 244976 201748
rect 246028 201696 246080 201748
rect 250076 201696 250128 201748
rect 250996 201696 251048 201748
rect 253112 201696 253164 201748
rect 253756 201696 253808 201748
rect 255228 201764 255280 201816
rect 259460 201696 259512 201748
rect 266268 201832 266320 201884
rect 269120 201832 269172 201884
rect 297732 201832 297784 201884
rect 264888 201764 264940 201816
rect 267740 201764 267792 201816
rect 298652 201764 298704 201816
rect 314936 201764 314988 201816
rect 315948 201764 316000 201816
rect 266636 201696 266688 201748
rect 267096 201696 267148 201748
rect 268200 201696 268252 201748
rect 297824 201696 297876 201748
rect 303896 201696 303948 201748
rect 306472 201696 306524 201748
rect 307300 201696 307352 201748
rect 351000 201696 351052 201748
rect 351828 201696 351880 201748
rect 355324 201696 355376 201748
rect 355968 201696 356020 201748
rect 243176 201628 243228 201680
rect 252376 201628 252428 201680
rect 263600 201628 263652 201680
rect 273628 201628 273680 201680
rect 279516 201628 279568 201680
rect 297548 201628 297600 201680
rect 305644 201628 305696 201680
rect 353576 201628 353628 201680
rect 356704 201628 356756 201680
rect 126336 201560 126388 201612
rect 134156 201560 134208 201612
rect 199660 201560 199712 201612
rect 216864 201560 216916 201612
rect 238208 201560 238260 201612
rect 245660 201560 245712 201612
rect 260840 201560 260892 201612
rect 266728 201560 266780 201612
rect 267004 201560 267056 201612
rect 267740 201560 267792 201612
rect 293776 201560 293828 201612
rect 294696 201560 294748 201612
rect 308404 201560 308456 201612
rect 308956 201560 309008 201612
rect 127624 201492 127676 201544
rect 134340 201492 134392 201544
rect 198556 201492 198608 201544
rect 202880 201492 202932 201544
rect 212448 201492 212500 201544
rect 220084 201492 220136 201544
rect 246488 201492 246540 201544
rect 254860 201492 254912 201544
rect 260104 201492 260156 201544
rect 267648 201492 267700 201544
rect 293040 201492 293092 201544
rect 293868 201492 293920 201544
rect 294420 201492 294472 201544
rect 295248 201492 295300 201544
rect 295800 201492 295852 201544
rect 296628 201492 296680 201544
rect 307024 201492 307076 201544
rect 314660 201560 314712 201612
rect 316040 201492 316092 201544
rect 317144 201492 317196 201544
rect 319076 201492 319128 201544
rect 320088 201492 320140 201544
rect 320548 201492 320600 201544
rect 321468 201492 321520 201544
rect 324044 201492 324096 201544
rect 327080 201492 327132 201544
rect 410156 201492 410208 201544
rect 411168 201492 411220 201544
rect 133512 201152 133564 201204
rect 153384 201152 153436 201204
rect 3884 201084 3936 201136
rect 436560 201084 436612 201136
rect 3608 201016 3660 201068
rect 436468 201016 436520 201068
rect 3424 200948 3476 201000
rect 436376 200948 436428 201000
rect 132408 200880 132460 200932
rect 580264 200880 580316 200932
rect 132224 200812 132276 200864
rect 580448 200812 580500 200864
rect 131396 200744 131448 200796
rect 580356 200744 580408 200796
rect 209872 200200 209924 200252
rect 210286 200200 210338 200252
rect 213920 200200 213972 200252
rect 214610 200200 214662 200252
rect 3240 200132 3292 200184
rect 436652 200132 436704 200184
rect 134248 200064 134300 200116
rect 238760 199860 238812 199912
rect 239496 199860 239548 199912
rect 243084 199860 243136 199912
rect 243820 199860 243872 199912
rect 133604 199792 133656 199844
rect 580264 199792 580316 199844
rect 131396 198296 131448 198348
rect 3424 197344 3476 197396
rect 131396 197344 131448 197396
rect 5356 196256 5408 196308
rect 131396 196256 131448 196308
rect 17224 196052 17276 196104
rect 130844 196052 130896 196104
rect 131764 196095 131816 196104
rect 131764 196061 131773 196095
rect 131773 196061 131807 196095
rect 131807 196061 131816 196095
rect 131764 196052 131816 196061
rect 132868 196095 132920 196104
rect 132868 196061 132877 196095
rect 132877 196061 132911 196095
rect 132911 196061 132920 196095
rect 132868 196052 132920 196061
rect 128544 195984 128596 196036
rect 131396 195984 131448 196036
rect 131764 195959 131816 195968
rect 131764 195925 131773 195959
rect 131773 195925 131807 195959
rect 131807 195925 131816 195959
rect 131764 195916 131816 195925
rect 132868 195959 132920 195968
rect 132868 195925 132877 195959
rect 132877 195925 132911 195959
rect 132911 195925 132920 195959
rect 132868 195916 132920 195925
rect 134064 195959 134116 195968
rect 134064 195925 134073 195959
rect 134073 195925 134107 195959
rect 134107 195925 134116 195959
rect 134064 195916 134116 195925
rect 128636 195848 128688 195900
rect 15844 194624 15896 194676
rect 130844 194624 130896 194676
rect 14464 194488 14516 194540
rect 130844 194488 130896 194540
rect 5264 193128 5316 193180
rect 130752 193128 130804 193180
rect 5448 193060 5500 193112
rect 130844 193060 130896 193112
rect 5172 191768 5224 191820
rect 130844 191768 130896 191820
rect 128636 191743 128688 191752
rect 128636 191709 128645 191743
rect 128645 191709 128679 191743
rect 128679 191709 128688 191743
rect 128636 191700 128688 191709
rect 129004 191743 129056 191752
rect 129004 191709 129013 191743
rect 129013 191709 129047 191743
rect 129047 191709 129056 191743
rect 129004 191700 129056 191709
rect 5080 190408 5132 190460
rect 130844 190408 130896 190460
rect 3516 188980 3568 189032
rect 130752 188980 130804 189032
rect 4988 188912 5040 188964
rect 130844 188912 130896 188964
rect 4896 187620 4948 187672
rect 130844 187620 130896 187672
rect 4804 186260 4856 186312
rect 128636 186235 128688 186244
rect 128636 186201 128645 186235
rect 128645 186201 128679 186235
rect 128679 186201 128688 186235
rect 128636 186192 128688 186201
rect 131212 186260 131264 186312
rect 131212 186124 131264 186176
rect 13084 184832 13136 184884
rect 131212 184832 131264 184884
rect 129004 183923 129056 183932
rect 129004 183889 129013 183923
rect 129013 183889 129047 183923
rect 129047 183889 129056 183923
rect 129004 183880 129056 183889
rect 72424 183472 72476 183524
rect 131212 183472 131264 183524
rect 131212 183336 131264 183388
rect 128820 182112 128872 182164
rect 128728 182044 128780 182096
rect 128912 182044 128964 182096
rect 132868 181432 132920 181484
rect 133328 181432 133380 181484
rect 2872 180752 2924 180804
rect 15844 180752 15896 180804
rect 133972 180387 134024 180396
rect 133972 180353 133981 180387
rect 133981 180353 134015 180387
rect 134015 180353 134024 180387
rect 133972 180344 134024 180353
rect 133880 176604 133932 176656
rect 134064 176604 134116 176656
rect 504456 173884 504508 173936
rect 504640 173884 504692 173936
rect 128636 172567 128688 172576
rect 128636 172533 128645 172567
rect 128645 172533 128679 172567
rect 128679 172533 128688 172567
rect 128636 172524 128688 172533
rect 133972 172567 134024 172576
rect 133972 172533 133981 172567
rect 133981 172533 134015 172567
rect 134015 172533 134024 172567
rect 133972 172524 134024 172533
rect 128912 167016 128964 167068
rect 128912 166880 128964 166932
rect 132592 164704 132644 164756
rect 133328 164704 133380 164756
rect 128636 164160 128688 164212
rect 128728 164160 128780 164212
rect 132592 164160 132644 164212
rect 504180 164160 504232 164212
rect 504364 164160 504416 164212
rect 132776 164092 132828 164144
rect 128636 162843 128688 162852
rect 128636 162809 128645 162843
rect 128645 162809 128679 162843
rect 128679 162809 128688 162843
rect 128636 162800 128688 162809
rect 133972 162800 134024 162852
rect 436836 157360 436888 157412
rect 580172 157360 580224 157412
rect 131120 156272 131172 156324
rect 3516 156068 3568 156120
rect 131304 156068 131356 156120
rect 3240 156000 3292 156052
rect 131120 156000 131172 156052
rect 131304 155932 131356 155984
rect 3608 155864 3660 155916
rect 131120 155864 131172 155916
rect 436100 155184 436152 155236
rect 438124 155184 438176 155236
rect 131212 155048 131264 155100
rect 132684 155048 132736 155100
rect 131120 154368 131172 154420
rect 3332 154300 3384 154352
rect 128636 153255 128688 153264
rect 128636 153221 128645 153255
rect 128645 153221 128679 153255
rect 128679 153221 128688 153255
rect 128636 153212 128688 153221
rect 4068 153144 4120 153196
rect 131120 153144 131172 153196
rect 437388 153144 437440 153196
rect 447784 153144 447836 153196
rect 131304 153119 131356 153128
rect 131304 153085 131313 153119
rect 131313 153085 131347 153119
rect 131347 153085 131356 153119
rect 131304 153076 131356 153085
rect 3976 152872 4028 152924
rect 131304 152940 131356 152992
rect 131304 151895 131356 151904
rect 131304 151861 131313 151895
rect 131313 151861 131347 151895
rect 131347 151861 131356 151895
rect 131304 151852 131356 151861
rect 3792 151716 3844 151768
rect 131120 151716 131172 151768
rect 3700 150356 3752 150408
rect 131120 150356 131172 150408
rect 437388 150356 437440 150408
rect 446404 150356 446456 150408
rect 28264 148996 28316 149048
rect 31024 148928 31076 148980
rect 131120 148928 131172 148980
rect 436100 148996 436152 149048
rect 445024 148996 445076 149048
rect 131120 148588 131172 148640
rect 128636 147747 128688 147756
rect 128636 147713 128645 147747
rect 128645 147713 128679 147747
rect 128679 147713 128688 147747
rect 128636 147704 128688 147713
rect 21364 147568 21416 147620
rect 131212 147611 131264 147620
rect 128636 147543 128688 147552
rect 128636 147509 128645 147543
rect 128645 147509 128679 147543
rect 128679 147509 128688 147543
rect 128636 147500 128688 147509
rect 131212 147577 131221 147611
rect 131221 147577 131255 147611
rect 131255 147577 131264 147611
rect 131212 147568 131264 147577
rect 131212 147432 131264 147484
rect 19984 146208 20036 146260
rect 131120 146208 131172 146260
rect 437388 146140 437440 146192
rect 442264 146140 442316 146192
rect 128912 144916 128964 144968
rect 128820 144848 128872 144900
rect 437020 144848 437072 144900
rect 514024 144848 514076 144900
rect 24768 144644 24820 144696
rect 128176 144712 128228 144764
rect 126244 144372 126296 144424
rect 131120 144372 131172 144424
rect 133972 143556 134024 143608
rect 132684 142103 132736 142112
rect 132684 142069 132693 142103
rect 132693 142069 132727 142103
rect 132727 142069 132736 142103
rect 132684 142060 132736 142069
rect 436100 142060 436152 142112
rect 438216 142060 438268 142112
rect 133880 138703 133932 138712
rect 133880 138669 133889 138703
rect 133889 138669 133923 138703
rect 133923 138669 133932 138703
rect 133880 138660 133932 138669
rect 437388 137912 437440 137964
rect 580540 137912 580592 137964
rect 3332 136552 3384 136604
rect 17224 136552 17276 136604
rect 437020 136552 437072 136604
rect 504456 136552 504508 136604
rect 132776 135192 132828 135244
rect 437388 133832 437440 133884
rect 580632 133832 580684 133884
rect 128636 132812 128688 132864
rect 128820 132812 128872 132864
rect 131212 132515 131264 132524
rect 131212 132481 131221 132515
rect 131221 132481 131255 132515
rect 131255 132481 131264 132515
rect 131212 132472 131264 132481
rect 132776 132404 132828 132456
rect 437388 132404 437440 132456
rect 580724 132404 580776 132456
rect 437388 129684 437440 129736
rect 580816 129684 580868 129736
rect 131120 125604 131172 125656
rect 131212 125604 131264 125656
rect 133880 125647 133932 125656
rect 133880 125613 133889 125647
rect 133889 125613 133923 125647
rect 133923 125613 133932 125647
rect 133880 125604 133932 125613
rect 131120 124151 131172 124160
rect 131120 124117 131129 124151
rect 131129 124117 131163 124151
rect 131163 124117 131172 124151
rect 131120 124108 131172 124117
rect 133880 121184 133932 121236
rect 580540 121184 580592 121236
rect 132408 121116 132460 121168
rect 580356 121116 580408 121168
rect 133972 121048 134024 121100
rect 580264 121048 580316 121100
rect 3056 120980 3108 121032
rect 436284 120980 436336 121032
rect 134064 120912 134116 120964
rect 180984 119756 181036 119808
rect 182042 119756 182094 119808
rect 185124 119756 185176 119808
rect 185722 119756 185774 119808
rect 138296 119348 138348 119400
rect 138848 119348 138900 119400
rect 143632 119348 143684 119400
rect 144368 119348 144420 119400
rect 67548 119076 67600 119128
rect 70308 119076 70360 119128
rect 130936 118872 130988 118924
rect 142252 118872 142304 118924
rect 142528 118872 142580 118924
rect 129648 118804 129700 118856
rect 145104 118804 145156 118856
rect 131028 118736 131080 118788
rect 147772 118736 147824 118788
rect 128728 118668 128780 118720
rect 128912 118668 128964 118720
rect 129556 118668 129608 118720
rect 149060 118668 149112 118720
rect 168380 118600 168432 118652
rect 178684 118600 178736 118652
rect 216680 118600 216732 118652
rect 217324 118600 217376 118652
rect 242256 118600 242308 118652
rect 75920 118532 75972 118584
rect 97908 118532 97960 118584
rect 181076 118532 181128 118584
rect 195888 118532 195940 118584
rect 234620 118532 234672 118584
rect 428464 118668 428516 118720
rect 258264 118600 258316 118652
rect 306012 118600 306064 118652
rect 332876 118600 332928 118652
rect 82728 118464 82780 118516
rect 164516 118464 164568 118516
rect 190368 118464 190420 118516
rect 231308 118464 231360 118516
rect 85488 118396 85540 118448
rect 71504 118328 71556 118380
rect 88340 118328 88392 118380
rect 113088 118396 113140 118448
rect 175556 118396 175608 118448
rect 186228 118396 186280 118448
rect 229468 118396 229520 118448
rect 230388 118396 230440 118448
rect 236184 118396 236236 118448
rect 238668 118396 238720 118448
rect 252744 118532 252796 118584
rect 257620 118532 257672 118584
rect 309692 118532 309744 118584
rect 339592 118600 339644 118652
rect 345848 118600 345900 118652
rect 396724 118600 396776 118652
rect 400864 118600 400916 118652
rect 480904 118600 480956 118652
rect 255320 118464 255372 118516
rect 257344 118464 257396 118516
rect 264336 118464 264388 118516
rect 310888 118464 310940 118516
rect 255780 118396 255832 118448
rect 308496 118396 308548 118448
rect 338396 118532 338448 118584
rect 362316 118532 362368 118584
rect 443000 118532 443052 118584
rect 341340 118464 341392 118516
rect 347596 118464 347648 118516
rect 376024 118464 376076 118516
rect 393596 118464 393648 118516
rect 475384 118464 475436 118516
rect 334808 118396 334860 118448
rect 335268 118396 335320 118448
rect 342168 118396 342220 118448
rect 389824 118396 389876 118448
rect 397276 118396 397328 118448
rect 478144 118396 478196 118448
rect 149888 118328 149940 118380
rect 194508 118328 194560 118380
rect 233240 118328 233292 118380
rect 234528 118328 234580 118380
rect 253940 118328 253992 118380
rect 256608 118328 256660 118380
rect 265532 118328 265584 118380
rect 311532 118328 311584 118380
rect 343916 118328 343968 118380
rect 365996 118328 366048 118380
rect 449900 118328 449952 118380
rect 71688 118260 71740 118312
rect 73896 118260 73948 118312
rect 82636 118260 82688 118312
rect 31668 118192 31720 118244
rect 107568 118192 107620 118244
rect 108304 118192 108356 118244
rect 125876 118260 125928 118312
rect 126888 118260 126940 118312
rect 129280 118260 129332 118312
rect 182916 118260 182968 118312
rect 184848 118260 184900 118312
rect 229192 118260 229244 118312
rect 231768 118260 231820 118312
rect 126244 118192 126296 118244
rect 126980 118192 127032 118244
rect 129188 118192 129240 118244
rect 177396 118192 177448 118244
rect 180064 118192 180116 118244
rect 225144 118192 225196 118244
rect 236828 118192 236880 118244
rect 237196 118192 237248 118244
rect 249800 118260 249852 118312
rect 251456 118260 251508 118312
rect 251548 118260 251600 118312
rect 256976 118260 257028 118312
rect 257988 118260 258040 118312
rect 266360 118260 266412 118312
rect 296168 118260 296220 118312
rect 305644 118260 305696 118312
rect 307208 118260 307260 118312
rect 334624 118260 334676 118312
rect 336648 118260 336700 118312
rect 374644 118260 374696 118312
rect 377036 118260 377088 118312
rect 469864 118260 469916 118312
rect 254676 118192 254728 118244
rect 263692 118192 263744 118244
rect 293776 118192 293828 118244
rect 302884 118192 302936 118244
rect 307668 118192 307720 118244
rect 336924 118192 336976 118244
rect 338488 118192 338540 118244
rect 384212 118192 384264 118244
rect 386236 118192 386288 118244
rect 389916 118192 389968 118244
rect 474004 118192 474056 118244
rect 28908 118124 28960 118176
rect 111708 118124 111760 118176
rect 23388 118056 23440 118108
rect 110328 118056 110380 118108
rect 113088 118056 113140 118108
rect 125692 118056 125744 118108
rect 126980 118056 127032 118108
rect 129648 118056 129700 118108
rect 173900 118124 173952 118176
rect 174544 118124 174596 118176
rect 220084 118124 220136 118176
rect 170036 118056 170088 118108
rect 179328 118056 179380 118108
rect 225788 118056 225840 118108
rect 227628 118056 227680 118108
rect 247224 118056 247276 118108
rect 250260 118056 250312 118108
rect 60648 117988 60700 118040
rect 88340 117988 88392 118040
rect 179420 117988 179472 118040
rect 183468 117988 183520 118040
rect 227720 117988 227772 118040
rect 229008 117988 229060 118040
rect 9588 117920 9640 117972
rect 70216 117920 70268 117972
rect 73896 117920 73948 117972
rect 107568 117920 107620 117972
rect 128912 117920 128964 117972
rect 129648 117920 129700 117972
rect 142160 117920 142212 117972
rect 143080 117920 143132 117972
rect 156512 117920 156564 117972
rect 156880 117920 156932 117972
rect 171876 117920 171928 117972
rect 176568 117920 176620 117972
rect 223948 117920 224000 117972
rect 226248 117920 226300 117972
rect 244280 117920 244332 117972
rect 122104 117852 122156 117904
rect 122564 117852 122616 117904
rect 160836 117852 160888 117904
rect 197268 117852 197320 117904
rect 234988 117852 235040 117904
rect 235356 117852 235408 117904
rect 245476 117988 245528 118040
rect 260012 118124 260064 118176
rect 295616 118124 295668 118176
rect 308404 118124 308456 118176
rect 345112 118124 345164 118176
rect 349436 118124 349488 118176
rect 369676 118124 369728 118176
rect 456800 118124 456852 118176
rect 252100 117988 252152 118040
rect 252468 118056 252520 118108
rect 263140 118056 263192 118108
rect 263416 118056 263468 118108
rect 269212 118056 269264 118108
rect 284576 118056 284628 118108
rect 291384 118056 291436 118108
rect 296628 118056 296680 118108
rect 314844 118056 314896 118108
rect 354312 118056 354364 118108
rect 369216 118056 369268 118108
rect 373356 118056 373408 118108
rect 463700 118056 463752 118108
rect 255228 117988 255280 118040
rect 264980 117988 265032 118040
rect 283932 117988 283984 118040
rect 290096 117988 290148 118040
rect 298652 117988 298704 118040
rect 318984 117988 319036 118040
rect 321928 117988 321980 118040
rect 363512 117988 363564 118040
rect 470600 117988 470652 118040
rect 251088 117920 251140 117972
rect 262496 117920 262548 117972
rect 263508 117920 263560 117972
rect 268660 117920 268712 117972
rect 294328 117920 294380 117972
rect 295248 117920 295300 117972
rect 297456 117920 297508 117972
rect 298008 117920 298060 117972
rect 300492 117920 300544 117972
rect 321744 117920 321796 117972
rect 354312 117920 354364 117972
rect 358176 117920 358228 117972
rect 380716 117920 380768 117972
rect 477500 117920 477552 117972
rect 120724 117716 120776 117768
rect 126888 117716 126940 117768
rect 162860 117784 162912 117836
rect 201408 117784 201460 117836
rect 233884 117784 233936 117836
rect 238852 117784 238904 117836
rect 240048 117784 240100 117836
rect 248972 117784 249024 117836
rect 256700 117852 256752 117904
rect 262128 117852 262180 117904
rect 268016 117852 268068 117904
rect 288900 117852 288952 117904
rect 251272 117784 251324 117836
rect 293132 117852 293184 117904
rect 293868 117852 293920 117904
rect 304816 117852 304868 117904
rect 297364 117784 297416 117836
rect 311808 117852 311860 117904
rect 333980 117852 334032 117904
rect 353116 117852 353168 117904
rect 425060 117852 425112 117904
rect 425152 117852 425204 117904
rect 511264 117852 511316 117904
rect 331312 117784 331364 117836
rect 332968 117784 333020 117836
rect 333888 117784 333940 117836
rect 416780 117784 416832 117836
rect 419264 117784 419316 117836
rect 420184 117784 420236 117836
rect 129096 117716 129148 117768
rect 166356 117716 166408 117768
rect 208308 117716 208360 117768
rect 240416 117716 240468 117768
rect 243544 117716 243596 117768
rect 244188 117716 244240 117768
rect 258816 117716 258868 117768
rect 302148 117716 302200 117768
rect 329288 117716 329340 117768
rect 357992 117716 358044 117768
rect 364064 117716 364116 117768
rect 402244 117716 402296 117768
rect 411904 117716 411956 117768
rect 415308 117716 415360 117768
rect 500224 117784 500276 117836
rect 422944 117716 422996 117768
rect 424324 117716 424376 117768
rect 426348 117716 426400 117768
rect 507124 117716 507176 117768
rect 157340 117648 157392 117700
rect 185584 117648 185636 117700
rect 209228 117648 209280 117700
rect 211068 117648 211120 117700
rect 241704 117648 241756 117700
rect 245568 117648 245620 117700
rect 259460 117648 259512 117700
rect 304172 117648 304224 117700
rect 329840 117648 329892 117700
rect 130384 117580 130436 117632
rect 158996 117580 159048 117632
rect 192484 117580 192536 117632
rect 211160 117580 211212 117632
rect 213828 117580 213880 117632
rect 238024 117580 238076 117632
rect 129464 117512 129516 117564
rect 152004 117512 152056 117564
rect 155316 117512 155368 117564
rect 198004 117512 198056 117564
rect 209964 117512 210016 117564
rect 220268 117512 220320 117564
rect 224224 117512 224276 117564
rect 129372 117444 129424 117496
rect 135444 117444 135496 117496
rect 141884 117444 141936 117496
rect 213184 117444 213236 117496
rect 226984 117444 227036 117496
rect 228364 117444 228416 117496
rect 243636 117512 243688 117564
rect 247684 117580 247736 117632
rect 260840 117580 260892 117632
rect 294972 117580 295024 117632
rect 311900 117580 311952 117632
rect 314568 117580 314620 117632
rect 247776 117512 247828 117564
rect 245936 117444 245988 117496
rect 249708 117512 249760 117564
rect 262220 117512 262272 117564
rect 266268 117512 266320 117564
rect 270500 117512 270552 117564
rect 280068 117512 280120 117564
rect 283104 117512 283156 117564
rect 299848 117512 299900 117564
rect 315304 117512 315356 117564
rect 325424 117580 325476 117632
rect 356796 117648 356848 117700
rect 393964 117648 394016 117700
rect 404268 117648 404320 117700
rect 482284 117648 482336 117700
rect 330484 117580 330536 117632
rect 331036 117580 331088 117632
rect 354956 117580 355008 117632
rect 320824 117512 320876 117564
rect 358084 117512 358136 117564
rect 358636 117512 358688 117564
rect 359280 117580 359332 117632
rect 360108 117580 360160 117632
rect 360476 117580 360528 117632
rect 398104 117580 398156 117632
rect 408224 117580 408276 117632
rect 486424 117580 486476 117632
rect 369124 117512 369176 117564
rect 384396 117512 384448 117564
rect 413284 117512 413336 117564
rect 248328 117444 248380 117496
rect 261300 117444 261352 117496
rect 267648 117444 267700 117496
rect 271052 117444 271104 117496
rect 282736 117444 282788 117496
rect 284944 117444 284996 117496
rect 289452 117444 289504 117496
rect 294604 117444 294656 117496
rect 306656 117444 306708 117496
rect 320088 117444 320140 117496
rect 324964 117444 325016 117496
rect 326344 117444 326396 117496
rect 328092 117444 328144 117496
rect 328276 117444 328328 117496
rect 367836 117444 367888 117496
rect 377404 117444 377456 117496
rect 399668 117444 399720 117496
rect 400036 117444 400088 117496
rect 408868 117444 408920 117496
rect 409696 117444 409748 117496
rect 111708 117376 111760 117428
rect 148048 117376 148100 117428
rect 229744 117376 229796 117428
rect 235264 117376 235316 117428
rect 92388 117308 92440 117360
rect 97908 117308 97960 117360
rect 190276 117308 190328 117360
rect 190552 117308 190604 117360
rect 195980 117308 196032 117360
rect 225604 117308 225656 117360
rect 232412 117308 232464 117360
rect 132960 117240 133012 117292
rect 237288 117240 237340 117292
rect 241428 117308 241480 117360
rect 253296 117376 253348 117428
rect 261484 117376 261536 117428
rect 267740 117376 267792 117428
rect 269764 117376 269816 117428
rect 271880 117376 271932 117428
rect 272524 117376 272576 117428
rect 273536 117376 273588 117428
rect 278412 117376 278464 117428
rect 279148 117376 279200 117428
rect 282092 117376 282144 117428
rect 283564 117376 283616 117428
rect 290004 117376 290056 117428
rect 291108 117376 291160 117428
rect 316408 117376 316460 117428
rect 317328 117376 317380 117428
rect 318248 117376 318300 117428
rect 322204 117376 322256 117428
rect 344008 117376 344060 117428
rect 344928 117376 344980 117428
rect 371516 117376 371568 117428
rect 372528 117376 372580 117428
rect 405188 117376 405240 117428
rect 405648 117376 405700 117428
rect 410708 117376 410760 117428
rect 411168 117376 411220 117428
rect 413744 117376 413796 117428
rect 416044 117376 416096 117428
rect 250444 117308 250496 117360
rect 254584 117308 254636 117360
rect 259368 117308 259420 117360
rect 266820 117308 266872 117360
rect 268384 117308 268436 117360
rect 269856 117308 269908 117360
rect 273168 117308 273220 117360
rect 274180 117308 274232 117360
rect 277860 117308 277912 117360
rect 278872 117308 278924 117360
rect 279056 117308 279108 117360
rect 280344 117308 280396 117360
rect 280896 117308 280948 117360
rect 281356 117308 281408 117360
rect 283380 117308 283432 117360
rect 284208 117308 284260 117360
rect 285220 117308 285272 117360
rect 285588 117308 285640 117360
rect 286416 117308 286468 117360
rect 286876 117308 286928 117360
rect 287612 117308 287664 117360
rect 288348 117308 288400 117360
rect 290740 117308 290792 117360
rect 291016 117308 291068 117360
rect 291936 117308 291988 117360
rect 292488 117308 292540 117360
rect 301136 117308 301188 117360
rect 302148 117308 302200 117360
rect 302976 117308 303028 117360
rect 303528 117308 303580 117360
rect 305368 117308 305420 117360
rect 306288 117308 306340 117360
rect 312728 117308 312780 117360
rect 313188 117308 313240 117360
rect 313924 117308 313976 117360
rect 314568 117308 314620 117360
rect 315212 117308 315264 117360
rect 315856 117308 315908 117360
rect 317052 117308 317104 117360
rect 317236 117308 317288 117360
rect 319444 117308 319496 117360
rect 320088 117308 320140 117360
rect 320732 117308 320784 117360
rect 321376 117308 321428 117360
rect 323768 117308 323820 117360
rect 324228 117308 324280 117360
rect 326252 117308 326304 117360
rect 326988 117308 327040 117360
rect 327448 117308 327500 117360
rect 328368 117308 328420 117360
rect 331680 117308 331732 117360
rect 332508 117308 332560 117360
rect 333520 117308 333572 117360
rect 333796 117308 333848 117360
rect 336004 117308 336056 117360
rect 336648 117308 336700 117360
rect 337200 117308 337252 117360
rect 338028 117308 338080 117360
rect 339040 117308 339092 117360
rect 339408 117308 339460 117360
rect 340328 117308 340380 117360
rect 340788 117308 340840 117360
rect 341524 117308 341576 117360
rect 342168 117308 342220 117360
rect 342720 117308 342772 117360
rect 343548 117308 343600 117360
rect 344560 117308 344612 117360
rect 344836 117308 344888 117360
rect 347044 117308 347096 117360
rect 347688 117308 347740 117360
rect 348240 117308 348292 117360
rect 349068 117308 349120 117360
rect 350080 117308 350132 117360
rect 350448 117308 350500 117360
rect 351276 117308 351328 117360
rect 351828 117308 351880 117360
rect 352564 117308 352616 117360
rect 353208 117308 353260 117360
rect 353760 117308 353812 117360
rect 354588 117308 354640 117360
rect 355600 117308 355652 117360
rect 355968 117308 356020 117360
rect 361120 117308 361172 117360
rect 361488 117308 361540 117360
rect 363604 117308 363656 117360
rect 364248 117308 364300 117360
rect 364800 117308 364852 117360
rect 365628 117308 365680 117360
rect 366640 117308 366692 117360
rect 367008 117308 367060 117360
rect 369032 117308 369084 117360
rect 369768 117308 369820 117360
rect 370320 117308 370372 117360
rect 371148 117308 371200 117360
rect 372160 117308 372212 117360
rect 372436 117308 372488 117360
rect 374552 117308 374604 117360
rect 375196 117308 375248 117360
rect 375840 117308 375892 117360
rect 376668 117308 376720 117360
rect 377680 117308 377732 117360
rect 378048 117308 378100 117360
rect 378876 117308 378928 117360
rect 379428 117308 379480 117360
rect 380072 117308 380124 117360
rect 380808 117308 380860 117360
rect 381360 117308 381412 117360
rect 382188 117308 382240 117360
rect 382556 117308 382608 117360
rect 383568 117308 383620 117360
rect 385592 117308 385644 117360
rect 386328 117308 386380 117360
rect 386788 117308 386840 117360
rect 387616 117308 387668 117360
rect 388076 117308 388128 117360
rect 389088 117308 389140 117360
rect 391112 117308 391164 117360
rect 391756 117308 391808 117360
rect 392308 117308 392360 117360
rect 393136 117308 393188 117360
rect 395436 117308 395488 117360
rect 395988 117308 396040 117360
rect 396632 117308 396684 117360
rect 397368 117308 397420 117360
rect 397828 117308 397880 117360
rect 398748 117308 398800 117360
rect 399116 117308 399168 117360
rect 400128 117308 400180 117360
rect 402152 117308 402204 117360
rect 402796 117308 402848 117360
rect 403348 117308 403400 117360
rect 404268 117308 404320 117360
rect 406384 117308 406436 117360
rect 407028 117308 407080 117360
rect 407672 117308 407724 117360
rect 408408 117308 408460 117360
rect 413192 117308 413244 117360
rect 413928 117308 413980 117360
rect 414388 117308 414440 117360
rect 415308 117308 415360 117360
rect 417424 117512 417476 117564
rect 420828 117512 420880 117564
rect 427268 117512 427320 117564
rect 427728 117512 427780 117564
rect 429844 117512 429896 117564
rect 430304 117512 430356 117564
rect 431224 117512 431276 117564
rect 431776 117512 431828 117564
rect 416228 117376 416280 117428
rect 416688 117376 416740 117428
rect 418620 117376 418672 117428
rect 419448 117376 419500 117428
rect 419908 117376 419960 117428
rect 420828 117376 420880 117428
rect 421748 117376 421800 117428
rect 422208 117376 422260 117428
rect 424140 117376 424192 117428
rect 424968 117376 425020 117428
rect 429660 117444 429712 117496
rect 430488 117444 430540 117496
rect 430948 117444 431000 117496
rect 431868 117444 431920 117496
rect 502984 117512 503036 117564
rect 432788 117444 432840 117496
rect 433248 117444 433300 117496
rect 425428 117376 425480 117428
rect 426348 117376 426400 117428
rect 493324 117376 493376 117428
rect 489184 117308 489236 117360
rect 192024 117104 192076 117156
rect 496084 116900 496136 116952
rect 190552 116764 190604 116816
rect 202972 116628 203024 116680
rect 203156 116628 203208 116680
rect 197360 116560 197412 116612
rect 198188 116560 198240 116612
rect 198740 116560 198792 116612
rect 199476 116560 199528 116612
rect 201500 116560 201552 116612
rect 201868 116560 201920 116612
rect 202880 116560 202932 116612
rect 203708 116560 203760 116612
rect 204260 116560 204312 116612
rect 204904 116560 204956 116612
rect 403716 116016 403768 116068
rect 403992 116016 404044 116068
rect 221464 115948 221516 116000
rect 221648 115948 221700 116000
rect 272248 115948 272300 116000
rect 272432 115948 272484 116000
rect 301412 115948 301464 116000
rect 301596 115948 301648 116000
rect 322388 115948 322440 116000
rect 322572 115948 322624 116000
rect 382924 115948 382976 116000
rect 383108 115948 383160 116000
rect 420276 115948 420328 116000
rect 420460 115948 420512 116000
rect 425888 115948 425940 116000
rect 425980 115948 426032 116000
rect 431316 115948 431368 116000
rect 431500 115948 431552 116000
rect 73896 115923 73948 115932
rect 73896 115889 73905 115923
rect 73905 115889 73939 115923
rect 73939 115889 73948 115923
rect 73896 115880 73948 115889
rect 133052 115923 133104 115932
rect 133052 115889 133061 115923
rect 133061 115889 133095 115923
rect 133095 115889 133104 115923
rect 133052 115880 133104 115889
rect 183744 115880 183796 115932
rect 183928 115880 183980 115932
rect 184756 115880 184808 115932
rect 185032 115880 185084 115932
rect 233424 115880 233476 115932
rect 233608 115880 233660 115932
rect 243636 115880 243688 115932
rect 243912 115880 243964 115932
rect 248328 115923 248380 115932
rect 248328 115889 248337 115923
rect 248337 115889 248371 115923
rect 248371 115889 248380 115923
rect 248328 115880 248380 115889
rect 341064 115880 341116 115932
rect 341340 115880 341392 115932
rect 388720 115880 388772 115932
rect 388904 115880 388956 115932
rect 403992 115880 404044 115932
rect 414848 115880 414900 115932
rect 414940 115880 414992 115932
rect 420460 115855 420512 115864
rect 420460 115821 420469 115855
rect 420469 115821 420503 115855
rect 420503 115821 420512 115855
rect 420460 115812 420512 115821
rect 131212 114520 131264 114572
rect 150900 114520 150952 114572
rect 151176 114520 151228 114572
rect 157432 114520 157484 114572
rect 157800 114520 157852 114572
rect 325700 114563 325752 114572
rect 325700 114529 325709 114563
rect 325709 114529 325743 114563
rect 325743 114529 325752 114563
rect 325700 114520 325752 114529
rect 243912 114452 243964 114504
rect 272248 114495 272300 114504
rect 272248 114461 272257 114495
rect 272257 114461 272291 114495
rect 272291 114461 272300 114495
rect 272248 114452 272300 114461
rect 213920 113976 213972 114028
rect 214196 113976 214248 114028
rect 133880 113840 133932 113892
rect 134524 113840 134576 113892
rect 135260 113840 135312 113892
rect 135720 113840 135772 113892
rect 136732 113840 136784 113892
rect 137560 113840 137612 113892
rect 139492 113840 139544 113892
rect 140044 113840 140096 113892
rect 140780 113840 140832 113892
rect 141240 113840 141292 113892
rect 146300 113840 146352 113892
rect 146760 113840 146812 113892
rect 153200 113840 153252 113892
rect 154120 113840 154172 113892
rect 161480 113840 161532 113892
rect 162124 113840 162176 113892
rect 167000 113840 167052 113892
rect 167644 113840 167696 113892
rect 169852 113840 169904 113892
rect 170680 113840 170732 113892
rect 189172 113840 189224 113892
rect 189632 113840 189684 113892
rect 191840 113840 191892 113892
rect 192668 113840 192720 113892
rect 213920 113840 213972 113892
rect 214104 113840 214156 113892
rect 215300 113840 215352 113892
rect 215944 113840 215996 113892
rect 218060 113840 218112 113892
rect 218428 113840 218480 113892
rect 219532 113840 219584 113892
rect 219716 113840 219768 113892
rect 222200 113840 222252 113892
rect 222660 113840 222712 113892
rect 231860 113840 231912 113892
rect 232504 113840 232556 113892
rect 248512 113840 248564 113892
rect 249064 113840 249116 113892
rect 173900 113160 173952 113212
rect 174360 113160 174412 113212
rect 175556 113160 175608 113212
rect 176200 113160 176252 113212
rect 178132 113160 178184 113212
rect 178592 113160 178644 113212
rect 179420 113160 179472 113212
rect 179880 113160 179932 113212
rect 180984 113135 181036 113144
rect 180984 113101 180993 113135
rect 180993 113101 181027 113135
rect 181027 113101 181036 113135
rect 180984 113092 181036 113101
rect 200212 113092 200264 113144
rect 200396 113092 200448 113144
rect 436928 111732 436980 111784
rect 579804 111732 579856 111784
rect 172520 111596 172572 111648
rect 173072 111596 173124 111648
rect 212632 110415 212684 110424
rect 212632 110381 212641 110415
rect 212641 110381 212675 110415
rect 212675 110381 212684 110415
rect 212632 110372 212684 110381
rect 194784 109692 194836 109744
rect 205916 109080 205968 109132
rect 207112 109080 207164 109132
rect 214104 109012 214156 109064
rect 214564 109012 214616 109064
rect 234712 109012 234764 109064
rect 235448 109012 235500 109064
rect 387524 109012 387576 109064
rect 387708 109012 387760 109064
rect 393044 109012 393096 109064
rect 393228 109012 393280 109064
rect 73896 108987 73948 108996
rect 73896 108953 73905 108987
rect 73905 108953 73939 108987
rect 73939 108953 73948 108987
rect 73896 108944 73948 108953
rect 205916 108944 205968 108996
rect 207112 108944 207164 108996
rect 420644 108944 420696 108996
rect 238852 106292 238904 106344
rect 238944 106292 238996 106344
rect 248328 106335 248380 106344
rect 248328 106301 248337 106335
rect 248337 106301 248371 106335
rect 248371 106301 248380 106335
rect 248328 106292 248380 106301
rect 403900 106335 403952 106344
rect 403900 106301 403909 106335
rect 403909 106301 403943 106335
rect 403943 106301 403952 106335
rect 403900 106292 403952 106301
rect 131304 106267 131356 106276
rect 131304 106233 131313 106267
rect 131313 106233 131347 106267
rect 131347 106233 131356 106267
rect 131304 106224 131356 106233
rect 301964 106267 302016 106276
rect 301964 106233 301973 106267
rect 301973 106233 302007 106267
rect 302007 106233 302016 106267
rect 301964 106224 302016 106233
rect 322664 106267 322716 106276
rect 322664 106233 322673 106267
rect 322673 106233 322707 106267
rect 322707 106233 322716 106267
rect 322664 106224 322716 106233
rect 388720 106224 388772 106276
rect 388812 106224 388864 106276
rect 394424 106267 394476 106276
rect 394424 106233 394433 106267
rect 394433 106233 394467 106267
rect 394467 106233 394476 106267
rect 394424 106224 394476 106233
rect 431684 106267 431736 106276
rect 431684 106233 431693 106267
rect 431693 106233 431727 106267
rect 431727 106233 431736 106267
rect 431684 106224 431736 106233
rect 183652 106156 183704 106208
rect 183928 106156 183980 106208
rect 148232 104864 148284 104916
rect 148508 104864 148560 104916
rect 194692 104907 194744 104916
rect 194692 104873 194701 104907
rect 194701 104873 194735 104907
rect 194735 104873 194744 104907
rect 194692 104864 194744 104873
rect 243728 104907 243780 104916
rect 243728 104873 243737 104907
rect 243737 104873 243771 104907
rect 243771 104873 243780 104907
rect 243728 104864 243780 104873
rect 274916 104864 274968 104916
rect 275376 104864 275428 104916
rect 133420 104796 133472 104848
rect 233424 104839 233476 104848
rect 233424 104805 233433 104839
rect 233433 104805 233467 104839
rect 233467 104805 233476 104839
rect 233424 104796 233476 104805
rect 248328 104796 248380 104848
rect 325700 104839 325752 104848
rect 325700 104805 325709 104839
rect 325709 104805 325743 104839
rect 325743 104805 325752 104839
rect 325700 104796 325752 104805
rect 415032 104839 415084 104848
rect 415032 104805 415041 104839
rect 415041 104805 415075 104839
rect 415075 104805 415084 104839
rect 415032 104796 415084 104805
rect 420644 104839 420696 104848
rect 420644 104805 420653 104839
rect 420653 104805 420687 104839
rect 420687 104805 420696 104839
rect 420644 104796 420696 104805
rect 181076 104728 181128 104780
rect 157248 103504 157300 103556
rect 157432 103504 157484 103556
rect 272064 103504 272116 103556
rect 173900 103436 173952 103488
rect 178132 103436 178184 103488
rect 178316 103436 178368 103488
rect 179420 103436 179472 103488
rect 279792 103436 279844 103488
rect 279976 103436 280028 103488
rect 173992 103368 174044 103420
rect 179512 103368 179564 103420
rect 212724 100716 212776 100768
rect 221096 100079 221148 100088
rect 221096 100045 221105 100079
rect 221105 100045 221139 100079
rect 221139 100045 221148 100079
rect 221096 100036 221148 100045
rect 73804 99356 73856 99408
rect 73988 99356 74040 99408
rect 150716 99424 150768 99476
rect 209872 99424 209924 99476
rect 229192 99424 229244 99476
rect 234712 99424 234764 99476
rect 240232 99424 240284 99476
rect 216772 99356 216824 99408
rect 243636 99356 243688 99408
rect 244372 99356 244424 99408
rect 244556 99356 244608 99408
rect 245844 99356 245896 99408
rect 246028 99356 246080 99408
rect 272064 99424 272116 99476
rect 341248 99356 341300 99408
rect 131304 99331 131356 99340
rect 131304 99297 131313 99331
rect 131313 99297 131347 99331
rect 131347 99297 131356 99331
rect 131304 99288 131356 99297
rect 150624 99288 150676 99340
rect 209872 99288 209924 99340
rect 229192 99288 229244 99340
rect 234712 99288 234764 99340
rect 240232 99288 240284 99340
rect 271972 99288 272024 99340
rect 301964 99331 302016 99340
rect 301964 99297 301973 99331
rect 301973 99297 302007 99331
rect 302007 99297 302016 99331
rect 301964 99288 302016 99297
rect 322664 99331 322716 99340
rect 322664 99297 322673 99331
rect 322673 99297 322707 99331
rect 322707 99297 322716 99331
rect 322664 99288 322716 99297
rect 383292 99424 383344 99476
rect 403900 99356 403952 99408
rect 341340 99288 341392 99340
rect 383200 99288 383252 99340
rect 394424 99331 394476 99340
rect 394424 99297 394433 99331
rect 394433 99297 394467 99331
rect 394467 99297 394476 99331
rect 394424 99288 394476 99297
rect 403992 99288 404044 99340
rect 431684 99331 431736 99340
rect 431684 99297 431693 99331
rect 431693 99297 431727 99331
rect 431727 99297 431736 99331
rect 431684 99288 431736 99297
rect 227720 96611 227772 96620
rect 227720 96577 227729 96611
rect 227729 96577 227763 96611
rect 227763 96577 227772 96611
rect 227720 96568 227772 96577
rect 238852 96611 238904 96620
rect 238852 96577 238861 96611
rect 238861 96577 238895 96611
rect 238895 96577 238904 96611
rect 238852 96568 238904 96577
rect 341064 96568 341116 96620
rect 341340 96568 341392 96620
rect 383200 96568 383252 96620
rect 388720 96568 388772 96620
rect 403992 96568 404044 96620
rect 145104 95344 145156 95396
rect 133144 95251 133196 95260
rect 133144 95217 133153 95251
rect 133153 95217 133187 95251
rect 133187 95217 133196 95251
rect 133144 95208 133196 95217
rect 145104 95208 145156 95260
rect 147956 95208 148008 95260
rect 148232 95208 148284 95260
rect 181076 95208 181128 95260
rect 221188 95208 221240 95260
rect 233516 95208 233568 95260
rect 243728 95251 243780 95260
rect 243728 95217 243737 95251
rect 243737 95217 243771 95251
rect 243771 95217 243780 95251
rect 243728 95208 243780 95217
rect 248236 95251 248288 95260
rect 248236 95217 248245 95251
rect 248245 95217 248279 95251
rect 248279 95217 248288 95251
rect 248236 95208 248288 95217
rect 325700 95251 325752 95260
rect 325700 95217 325709 95251
rect 325709 95217 325743 95251
rect 325743 95217 325752 95251
rect 325700 95208 325752 95217
rect 415216 95208 415268 95260
rect 420644 95251 420696 95260
rect 420644 95217 420653 95251
rect 420653 95217 420687 95251
rect 420687 95217 420696 95251
rect 420644 95208 420696 95217
rect 426256 95140 426308 95192
rect 181168 95072 181220 95124
rect 162860 93848 162912 93900
rect 163044 93848 163096 93900
rect 206008 93916 206060 93968
rect 156052 93823 156104 93832
rect 156052 93789 156061 93823
rect 156061 93789 156095 93823
rect 156095 93789 156104 93823
rect 156052 93780 156104 93789
rect 205916 93780 205968 93832
rect 279700 93823 279752 93832
rect 279700 93789 279709 93823
rect 279709 93789 279743 93823
rect 279743 93789 279752 93823
rect 279700 93780 279752 93789
rect 2780 93304 2832 93356
rect 5356 93304 5408 93356
rect 181168 92463 181220 92472
rect 181168 92429 181177 92463
rect 181177 92429 181211 92463
rect 181211 92429 181220 92463
rect 181168 92420 181220 92429
rect 212724 91060 212776 91112
rect 212908 91060 212960 91112
rect 216680 91103 216732 91112
rect 216680 91069 216689 91103
rect 216689 91069 216723 91103
rect 216723 91069 216732 91103
rect 216680 91060 216732 91069
rect 207112 91035 207164 91044
rect 207112 91001 207121 91035
rect 207121 91001 207155 91035
rect 207155 91001 207164 91035
rect 207112 90992 207164 91001
rect 145104 90380 145156 90432
rect 73804 89836 73856 89888
rect 194784 89700 194836 89752
rect 243728 89700 243780 89752
rect 322572 89700 322624 89752
rect 322756 89700 322808 89752
rect 394332 89700 394384 89752
rect 394516 89700 394568 89752
rect 227812 89632 227864 89684
rect 238852 89675 238904 89684
rect 238852 89641 238861 89675
rect 238861 89641 238895 89675
rect 238895 89641 238904 89675
rect 238852 89632 238904 89641
rect 415216 89768 415268 89820
rect 420644 89700 420696 89752
rect 415124 89632 415176 89684
rect 194876 89564 194928 89616
rect 243728 89564 243780 89616
rect 420644 89564 420696 89616
rect 179512 88995 179564 89004
rect 179512 88961 179521 88995
rect 179521 88961 179555 88995
rect 179555 88961 179564 88995
rect 179512 88952 179564 88961
rect 131396 88272 131448 88324
rect 580172 88272 580224 88324
rect 248236 87116 248288 87168
rect 73712 87023 73764 87032
rect 73712 86989 73721 87023
rect 73721 86989 73755 87023
rect 73755 86989 73764 87023
rect 73712 86980 73764 86989
rect 233424 86980 233476 87032
rect 233516 86980 233568 87032
rect 248328 86980 248380 87032
rect 271880 86980 271932 87032
rect 383108 87023 383160 87032
rect 383108 86989 383117 87023
rect 383117 86989 383151 87023
rect 383151 86989 383160 87023
rect 383108 86980 383160 86989
rect 388628 87023 388680 87032
rect 388628 86989 388637 87023
rect 388637 86989 388671 87023
rect 388671 86989 388680 87023
rect 388628 86980 388680 86989
rect 403900 87023 403952 87032
rect 403900 86989 403909 87023
rect 403909 86989 403943 87023
rect 403943 86989 403952 87023
rect 403900 86980 403952 86989
rect 183744 86912 183796 86964
rect 183928 86912 183980 86964
rect 190736 86955 190788 86964
rect 190736 86921 190745 86955
rect 190745 86921 190779 86955
rect 190779 86921 190788 86955
rect 190736 86912 190788 86921
rect 243728 86955 243780 86964
rect 243728 86921 243737 86955
rect 243737 86921 243771 86955
rect 243771 86921 243780 86955
rect 243728 86912 243780 86921
rect 245936 86912 245988 86964
rect 274916 86912 274968 86964
rect 322664 86955 322716 86964
rect 322664 86921 322673 86955
rect 322673 86921 322707 86955
rect 322707 86921 322716 86955
rect 322664 86912 322716 86921
rect 394424 86955 394476 86964
rect 394424 86921 394433 86955
rect 394433 86921 394467 86955
rect 394467 86921 394476 86955
rect 394424 86912 394476 86921
rect 233424 86887 233476 86896
rect 233424 86853 233433 86887
rect 233433 86853 233467 86887
rect 233467 86853 233476 86887
rect 233424 86844 233476 86853
rect 271880 86844 271932 86896
rect 150624 85620 150676 85672
rect 144920 85595 144972 85604
rect 144920 85561 144929 85595
rect 144929 85561 144963 85595
rect 144963 85561 144972 85595
rect 144920 85552 144972 85561
rect 150532 85552 150584 85604
rect 426164 85595 426216 85604
rect 426164 85561 426173 85595
rect 426173 85561 426207 85595
rect 426207 85561 426216 85595
rect 426164 85552 426216 85561
rect 194876 85527 194928 85536
rect 194876 85493 194885 85527
rect 194885 85493 194919 85527
rect 194919 85493 194928 85527
rect 194876 85484 194928 85493
rect 200304 85527 200356 85536
rect 200304 85493 200313 85527
rect 200313 85493 200347 85527
rect 200347 85493 200356 85527
rect 200304 85484 200356 85493
rect 248328 85527 248380 85536
rect 248328 85493 248337 85527
rect 248337 85493 248371 85527
rect 248371 85493 248380 85527
rect 248328 85484 248380 85493
rect 325700 85527 325752 85536
rect 325700 85493 325709 85527
rect 325709 85493 325743 85527
rect 325743 85493 325752 85527
rect 325700 85484 325752 85493
rect 279700 84303 279752 84312
rect 279700 84269 279709 84303
rect 279709 84269 279743 84303
rect 279743 84269 279752 84303
rect 279700 84260 279752 84269
rect 156144 84192 156196 84244
rect 179604 84192 179656 84244
rect 162860 84167 162912 84176
rect 162860 84133 162869 84167
rect 162869 84133 162903 84167
rect 162903 84133 162912 84167
rect 162860 84124 162912 84133
rect 279700 84167 279752 84176
rect 279700 84133 279709 84167
rect 279709 84133 279743 84167
rect 279743 84133 279752 84167
rect 279700 84124 279752 84133
rect 426164 84124 426216 84176
rect 181260 82832 181312 82884
rect 227904 82127 227956 82136
rect 227904 82093 227913 82127
rect 227913 82093 227947 82127
rect 227947 82093 227956 82127
rect 227904 82084 227956 82093
rect 420276 82084 420328 82136
rect 420644 82084 420696 82136
rect 205916 81404 205968 81456
rect 206100 81404 206152 81456
rect 207204 81404 207256 81456
rect 211344 81404 211396 81456
rect 211436 81404 211488 81456
rect 238944 81447 238996 81456
rect 238944 81413 238953 81447
rect 238953 81413 238987 81447
rect 238987 81413 238996 81447
rect 238944 81404 238996 81413
rect 150532 80724 150584 80776
rect 150716 80724 150768 80776
rect 205916 80155 205968 80164
rect 205916 80121 205925 80155
rect 205925 80121 205959 80155
rect 205959 80121 205968 80155
rect 205916 80112 205968 80121
rect 207204 80155 207256 80164
rect 207204 80121 207213 80155
rect 207213 80121 207247 80155
rect 207247 80121 207256 80155
rect 207204 80112 207256 80121
rect 221096 80112 221148 80164
rect 229284 80112 229336 80164
rect 357992 80155 358044 80164
rect 357992 80121 358001 80155
rect 358001 80121 358035 80155
rect 358035 80121 358044 80155
rect 357992 80112 358044 80121
rect 229192 80044 229244 80096
rect 431592 80044 431644 80096
rect 431776 80044 431828 80096
rect 3240 79976 3292 80028
rect 434996 79976 435048 80028
rect 221004 79951 221056 79960
rect 221004 79917 221013 79951
rect 221013 79917 221047 79951
rect 221047 79917 221056 79951
rect 221004 79908 221056 79917
rect 357992 79951 358044 79960
rect 357992 79917 358001 79951
rect 358001 79917 358035 79951
rect 358035 79917 358044 79951
rect 357992 79908 358044 79917
rect 184848 77367 184900 77376
rect 184848 77333 184857 77367
rect 184857 77333 184891 77367
rect 184891 77333 184900 77367
rect 184848 77324 184900 77333
rect 301872 77324 301924 77376
rect 302056 77324 302108 77376
rect 128820 77256 128872 77308
rect 129004 77256 129056 77308
rect 190828 77256 190880 77308
rect 227996 77256 228048 77308
rect 233424 77299 233476 77308
rect 233424 77265 233433 77299
rect 233433 77265 233467 77299
rect 233467 77265 233476 77299
rect 233424 77256 233476 77265
rect 238944 77299 238996 77308
rect 238944 77265 238953 77299
rect 238953 77265 238987 77299
rect 238987 77265 238996 77299
rect 238944 77256 238996 77265
rect 243728 77299 243780 77308
rect 243728 77265 243737 77299
rect 243737 77265 243771 77299
rect 243771 77265 243780 77299
rect 243728 77256 243780 77265
rect 245752 77299 245804 77308
rect 245752 77265 245761 77299
rect 245761 77265 245795 77299
rect 245795 77265 245804 77299
rect 245752 77256 245804 77265
rect 274824 77299 274876 77308
rect 274824 77265 274833 77299
rect 274833 77265 274867 77299
rect 274867 77265 274876 77299
rect 274824 77256 274876 77265
rect 322756 77256 322808 77308
rect 394516 77256 394568 77308
rect 132132 77188 132184 77240
rect 580172 77188 580224 77240
rect 184848 77163 184900 77172
rect 184848 77129 184857 77163
rect 184857 77129 184891 77163
rect 184891 77129 184900 77163
rect 184848 77120 184900 77129
rect 302056 77120 302108 77172
rect 341340 77163 341392 77172
rect 341340 77129 341349 77163
rect 341349 77129 341383 77163
rect 341383 77129 341392 77163
rect 341340 77120 341392 77129
rect 383200 77163 383252 77172
rect 383200 77129 383209 77163
rect 383209 77129 383243 77163
rect 383243 77129 383252 77163
rect 383200 77120 383252 77129
rect 388720 77163 388772 77172
rect 388720 77129 388729 77163
rect 388729 77129 388763 77163
rect 388763 77129 388772 77163
rect 388720 77120 388772 77129
rect 403992 77163 404044 77172
rect 403992 77129 404001 77163
rect 404001 77129 404035 77163
rect 404035 77129 404044 77163
rect 403992 77120 404044 77129
rect 184756 77052 184808 77104
rect 185032 77052 185084 77104
rect 207204 76619 207256 76628
rect 207204 76585 207213 76619
rect 207213 76585 207247 76619
rect 207247 76585 207256 76619
rect 207204 76576 207256 76585
rect 173992 75896 174044 75948
rect 174084 75896 174136 75948
rect 181260 75964 181312 76016
rect 194876 75939 194928 75948
rect 194876 75905 194885 75939
rect 194885 75905 194919 75939
rect 194919 75905 194928 75939
rect 194876 75896 194928 75905
rect 200304 75939 200356 75948
rect 200304 75905 200313 75939
rect 200313 75905 200347 75939
rect 200347 75905 200356 75939
rect 200304 75896 200356 75905
rect 248328 75939 248380 75948
rect 248328 75905 248337 75939
rect 248337 75905 248371 75939
rect 248371 75905 248380 75939
rect 248328 75896 248380 75905
rect 325700 75939 325752 75948
rect 325700 75905 325709 75939
rect 325709 75905 325743 75939
rect 325743 75905 325752 75939
rect 325700 75896 325752 75905
rect 415032 75896 415084 75948
rect 415124 75896 415176 75948
rect 157432 75871 157484 75880
rect 157432 75837 157441 75871
rect 157441 75837 157475 75871
rect 157475 75837 157484 75871
rect 157432 75828 157484 75837
rect 178132 75828 178184 75880
rect 178316 75828 178368 75880
rect 181076 75828 181128 75880
rect 183928 75828 183980 75880
rect 211344 75828 211396 75880
rect 244280 75871 244332 75880
rect 244280 75837 244289 75871
rect 244289 75837 244323 75871
rect 244323 75837 244332 75871
rect 244280 75828 244332 75837
rect 245752 75871 245804 75880
rect 245752 75837 245761 75871
rect 245761 75837 245795 75871
rect 245795 75837 245804 75871
rect 245752 75828 245804 75837
rect 271880 75871 271932 75880
rect 271880 75837 271889 75871
rect 271889 75837 271923 75871
rect 271923 75837 271932 75871
rect 271880 75828 271932 75837
rect 431592 75871 431644 75880
rect 431592 75837 431601 75871
rect 431601 75837 431635 75871
rect 431635 75837 431644 75871
rect 431592 75828 431644 75837
rect 156052 74536 156104 74588
rect 156236 74536 156288 74588
rect 162860 74579 162912 74588
rect 162860 74545 162869 74579
rect 162869 74545 162903 74579
rect 162903 74545 162912 74579
rect 162860 74536 162912 74545
rect 279792 74536 279844 74588
rect 174084 74468 174136 74520
rect 205916 74103 205968 74112
rect 205916 74069 205925 74103
rect 205925 74069 205959 74103
rect 205959 74069 205968 74103
rect 205916 74060 205968 74069
rect 212816 73244 212868 73296
rect 212724 73176 212776 73228
rect 181076 73151 181128 73160
rect 181076 73117 181085 73151
rect 181085 73117 181119 73151
rect 181119 73117 181128 73151
rect 181076 73108 181128 73117
rect 150716 70456 150768 70508
rect 194876 70456 194928 70508
rect 209872 70499 209924 70508
rect 209872 70465 209881 70499
rect 209881 70465 209915 70499
rect 209915 70465 209924 70499
rect 209872 70456 209924 70465
rect 240232 70499 240284 70508
rect 240232 70465 240241 70499
rect 240241 70465 240275 70499
rect 240275 70465 240284 70499
rect 240232 70456 240284 70465
rect 279792 70388 279844 70440
rect 150624 70320 150676 70372
rect 194784 70320 194836 70372
rect 271972 70252 272024 70304
rect 279792 70252 279844 70304
rect 426072 69683 426124 69692
rect 426072 69649 426081 69683
rect 426081 69649 426115 69683
rect 426115 69649 426124 69683
rect 426072 69640 426124 69649
rect 212724 68391 212776 68400
rect 212724 68357 212733 68391
rect 212733 68357 212767 68391
rect 212767 68357 212776 68391
rect 212724 68348 212776 68357
rect 128728 67668 128780 67720
rect 190828 67668 190880 67720
rect 234712 67711 234764 67720
rect 234712 67677 234721 67711
rect 234721 67677 234755 67711
rect 234755 67677 234764 67711
rect 234712 67668 234764 67677
rect 128912 67600 128964 67652
rect 184756 67600 184808 67652
rect 184940 67600 184992 67652
rect 190736 67600 190788 67652
rect 200304 67600 200356 67652
rect 200396 67600 200448 67652
rect 209872 67643 209924 67652
rect 209872 67609 209881 67643
rect 209881 67609 209915 67643
rect 209915 67609 209924 67643
rect 209872 67600 209924 67609
rect 240232 67643 240284 67652
rect 240232 67609 240241 67643
rect 240241 67609 240275 67643
rect 240275 67609 240284 67643
rect 240232 67600 240284 67609
rect 301964 67643 302016 67652
rect 301964 67609 301973 67643
rect 301973 67609 302007 67643
rect 302007 67609 302016 67643
rect 301964 67600 302016 67609
rect 341432 67600 341484 67652
rect 383292 67600 383344 67652
rect 388812 67600 388864 67652
rect 394424 67600 394476 67652
rect 394516 67600 394568 67652
rect 404084 67600 404136 67652
rect 233424 67575 233476 67584
rect 233424 67541 233433 67575
rect 233433 67541 233467 67575
rect 233467 67541 233476 67575
rect 233424 67532 233476 67541
rect 145104 66308 145156 66360
rect 145288 66308 145340 66360
rect 183744 66351 183796 66360
rect 183744 66317 183753 66351
rect 183753 66317 183787 66351
rect 183787 66317 183796 66351
rect 183744 66308 183796 66317
rect 73804 66240 73856 66292
rect 73896 66240 73948 66292
rect 157432 66283 157484 66292
rect 157432 66249 157441 66283
rect 157441 66249 157475 66283
rect 157475 66249 157484 66283
rect 157432 66240 157484 66249
rect 179512 66240 179564 66292
rect 179604 66240 179656 66292
rect 211252 66283 211304 66292
rect 211252 66249 211261 66283
rect 211261 66249 211295 66283
rect 211295 66249 211304 66283
rect 211252 66240 211304 66249
rect 234712 66283 234764 66292
rect 234712 66249 234721 66283
rect 234721 66249 234755 66283
rect 234755 66249 234764 66283
rect 234712 66240 234764 66249
rect 244372 66240 244424 66292
rect 245844 66240 245896 66292
rect 322664 66240 322716 66292
rect 322756 66240 322808 66292
rect 420460 66240 420512 66292
rect 420552 66240 420604 66292
rect 431592 66283 431644 66292
rect 431592 66249 431601 66283
rect 431601 66249 431635 66283
rect 431635 66249 431644 66283
rect 431592 66240 431644 66249
rect 128912 66215 128964 66224
rect 128912 66181 128921 66215
rect 128921 66181 128955 66215
rect 128955 66181 128964 66215
rect 128912 66172 128964 66181
rect 183744 66215 183796 66224
rect 183744 66181 183753 66215
rect 183753 66181 183787 66215
rect 183787 66181 183796 66215
rect 183744 66172 183796 66181
rect 190736 66172 190788 66224
rect 190828 66172 190880 66224
rect 194784 66172 194836 66224
rect 207204 66172 207256 66224
rect 248328 66215 248380 66224
rect 248328 66181 248337 66215
rect 248337 66181 248371 66215
rect 248371 66181 248380 66215
rect 248328 66172 248380 66181
rect 325700 66172 325752 66224
rect 415032 66215 415084 66224
rect 415032 66181 415041 66215
rect 415041 66181 415075 66215
rect 415075 66181 415084 66215
rect 415032 66172 415084 66181
rect 420460 66104 420512 66156
rect 420644 66104 420696 66156
rect 173992 64923 174044 64932
rect 173992 64889 174001 64923
rect 174001 64889 174035 64923
rect 174035 64889 174044 64923
rect 173992 64880 174044 64889
rect 3332 64812 3384 64864
rect 131672 64812 131724 64864
rect 145104 64855 145156 64864
rect 145104 64821 145113 64855
rect 145113 64821 145147 64855
rect 145147 64821 145156 64855
rect 145104 64812 145156 64821
rect 147956 64855 148008 64864
rect 147956 64821 147965 64855
rect 147965 64821 147999 64855
rect 147999 64821 148008 64855
rect 147956 64812 148008 64821
rect 159088 64855 159140 64864
rect 159088 64821 159097 64855
rect 159097 64821 159131 64855
rect 159131 64821 159140 64855
rect 159088 64812 159140 64821
rect 162860 64812 162912 64864
rect 163136 64812 163188 64864
rect 178132 64812 178184 64864
rect 178316 64812 178368 64864
rect 436836 64812 436888 64864
rect 579804 64812 579856 64864
rect 181076 63563 181128 63572
rect 181076 63529 181085 63563
rect 181085 63529 181119 63563
rect 181119 63529 181128 63563
rect 181076 63520 181128 63529
rect 233424 62815 233476 62824
rect 233424 62781 233433 62815
rect 233433 62781 233467 62815
rect 233467 62781 233476 62815
rect 233424 62772 233476 62781
rect 181076 61004 181128 61056
rect 184940 60843 184992 60852
rect 184940 60809 184949 60843
rect 184949 60809 184983 60843
rect 184983 60809 184992 60843
rect 184940 60800 184992 60809
rect 205916 60800 205968 60852
rect 227996 60800 228048 60852
rect 243728 60800 243780 60852
rect 227904 60732 227956 60784
rect 150532 60664 150584 60716
rect 150716 60664 150768 60716
rect 156052 60664 156104 60716
rect 156236 60664 156288 60716
rect 216772 60664 216824 60716
rect 216956 60664 217008 60716
rect 221004 60664 221056 60716
rect 221188 60664 221240 60716
rect 383292 60800 383344 60852
rect 388812 60800 388864 60852
rect 404084 60800 404136 60852
rect 244372 60664 244424 60716
rect 244556 60664 244608 60716
rect 245844 60664 245896 60716
rect 246028 60664 246080 60716
rect 271972 60664 272024 60716
rect 272156 60664 272208 60716
rect 279884 60664 279936 60716
rect 280068 60664 280120 60716
rect 383200 60664 383252 60716
rect 388720 60664 388772 60716
rect 403992 60664 404044 60716
rect 243728 60596 243780 60648
rect 178224 59848 178276 59900
rect 178316 59848 178368 59900
rect 240232 58012 240284 58064
rect 73896 57944 73948 57996
rect 205824 57987 205876 57996
rect 205824 57953 205833 57987
rect 205833 57953 205867 57987
rect 205867 57953 205876 57987
rect 205824 57944 205876 57953
rect 133236 57876 133288 57928
rect 150716 57919 150768 57928
rect 150716 57885 150725 57919
rect 150725 57885 150759 57919
rect 150759 57885 150768 57919
rect 150716 57876 150768 57885
rect 184940 57919 184992 57928
rect 184940 57885 184949 57919
rect 184949 57885 184983 57919
rect 184983 57885 184992 57919
rect 184940 57876 184992 57885
rect 200396 57876 200448 57928
rect 212540 57919 212592 57928
rect 212540 57885 212549 57919
rect 212549 57885 212583 57919
rect 212583 57885 212592 57919
rect 212724 57919 212776 57928
rect 212540 57876 212592 57885
rect 212724 57885 212733 57919
rect 212733 57885 212767 57919
rect 212767 57885 212776 57919
rect 212724 57876 212776 57885
rect 216956 57876 217008 57928
rect 276112 57876 276164 57928
rect 276296 57876 276348 57928
rect 280068 57876 280120 57928
rect 301780 57919 301832 57928
rect 301780 57885 301789 57919
rect 301789 57885 301823 57919
rect 301823 57885 301832 57919
rect 301780 57876 301832 57885
rect 322756 57876 322808 57928
rect 383200 57919 383252 57928
rect 383200 57885 383209 57919
rect 383209 57885 383243 57919
rect 383243 57885 383252 57919
rect 383200 57876 383252 57885
rect 388720 57919 388772 57928
rect 388720 57885 388729 57919
rect 388729 57885 388763 57919
rect 388763 57885 388772 57919
rect 388720 57876 388772 57885
rect 403992 57919 404044 57928
rect 403992 57885 404001 57919
rect 404001 57885 404035 57919
rect 404035 57885 404044 57919
rect 403992 57876 404044 57885
rect 73988 57808 74040 57860
rect 129004 57808 129056 57860
rect 183744 56627 183796 56636
rect 183744 56593 183753 56627
rect 183753 56593 183787 56627
rect 183787 56593 183796 56627
rect 183744 56584 183796 56593
rect 195152 56627 195204 56636
rect 195152 56593 195161 56627
rect 195161 56593 195195 56627
rect 195195 56593 195204 56627
rect 207112 56627 207164 56636
rect 195152 56584 195204 56593
rect 207112 56593 207121 56627
rect 207121 56593 207155 56627
rect 207155 56593 207164 56627
rect 207112 56584 207164 56593
rect 240140 56627 240192 56636
rect 240140 56593 240149 56627
rect 240149 56593 240183 56627
rect 240183 56593 240192 56627
rect 248328 56627 248380 56636
rect 240140 56584 240192 56593
rect 248328 56593 248337 56627
rect 248337 56593 248371 56627
rect 248371 56593 248380 56627
rect 248328 56584 248380 56593
rect 325516 56627 325568 56636
rect 325516 56593 325525 56627
rect 325525 56593 325559 56627
rect 325559 56593 325568 56627
rect 325516 56584 325568 56593
rect 415032 56627 415084 56636
rect 415032 56593 415041 56627
rect 415041 56593 415075 56627
rect 415075 56593 415084 56627
rect 415032 56584 415084 56593
rect 145104 56559 145156 56568
rect 145104 56525 145113 56559
rect 145113 56525 145147 56559
rect 145147 56525 145156 56559
rect 145104 56516 145156 56525
rect 234712 56559 234764 56568
rect 234712 56525 234721 56559
rect 234721 56525 234755 56559
rect 234755 56525 234764 56559
rect 234712 56516 234764 56525
rect 431592 56516 431644 56568
rect 431776 56516 431828 56568
rect 147956 55267 148008 55276
rect 147956 55233 147965 55267
rect 147965 55233 147999 55267
rect 147999 55233 148008 55267
rect 147956 55224 148008 55233
rect 159088 55267 159140 55276
rect 159088 55233 159097 55267
rect 159097 55233 159131 55267
rect 159131 55233 159140 55267
rect 159088 55224 159140 55233
rect 173992 55224 174044 55276
rect 174084 55224 174136 55276
rect 175648 55224 175700 55276
rect 175832 55224 175884 55276
rect 227904 53159 227956 53168
rect 227904 53125 227913 53159
rect 227913 53125 227947 53159
rect 227947 53125 227956 53159
rect 227904 53116 227956 53125
rect 238852 53116 238904 53168
rect 239036 53116 239088 53168
rect 243452 53116 243504 53168
rect 243728 53116 243780 53168
rect 426072 53116 426124 53168
rect 426256 53116 426308 53168
rect 147956 51756 148008 51808
rect 148140 51756 148192 51808
rect 415032 51280 415084 51332
rect 415216 51280 415268 51332
rect 209872 51187 209924 51196
rect 209872 51153 209881 51187
rect 209881 51153 209915 51187
rect 209915 51153 209924 51187
rect 209872 51144 209924 51153
rect 341524 51187 341576 51196
rect 341524 51153 341533 51187
rect 341533 51153 341567 51187
rect 341567 51153 341576 51187
rect 341524 51144 341576 51153
rect 159088 51076 159140 51128
rect 179512 51076 179564 51128
rect 184940 51119 184992 51128
rect 184940 51085 184949 51119
rect 184949 51085 184983 51119
rect 184983 51085 184992 51119
rect 184940 51076 184992 51085
rect 212540 51119 212592 51128
rect 212540 51085 212549 51119
rect 212549 51085 212583 51119
rect 212583 51085 212592 51119
rect 212540 51076 212592 51085
rect 221188 51076 221240 51128
rect 244556 51076 244608 51128
rect 272156 51076 272208 51128
rect 179420 51008 179472 51060
rect 221096 51008 221148 51060
rect 244464 51008 244516 51060
rect 272064 51008 272116 51060
rect 357900 51008 357952 51060
rect 358084 51008 358136 51060
rect 159088 50940 159140 50992
rect 181168 50643 181220 50652
rect 181168 50609 181177 50643
rect 181177 50609 181211 50643
rect 181211 50609 181220 50643
rect 181168 50600 181220 50609
rect 133144 48331 133196 48340
rect 133144 48297 133153 48331
rect 133153 48297 133187 48331
rect 133187 48297 133196 48331
rect 133144 48288 133196 48297
rect 150808 48288 150860 48340
rect 184940 48331 184992 48340
rect 184940 48297 184949 48331
rect 184949 48297 184983 48331
rect 184983 48297 184992 48331
rect 184940 48288 184992 48297
rect 200304 48331 200356 48340
rect 200304 48297 200313 48331
rect 200313 48297 200347 48331
rect 200347 48297 200356 48331
rect 200304 48288 200356 48297
rect 216864 48331 216916 48340
rect 216864 48297 216873 48331
rect 216873 48297 216907 48331
rect 216907 48297 216916 48331
rect 216864 48288 216916 48297
rect 227996 48288 228048 48340
rect 240140 48288 240192 48340
rect 240232 48288 240284 48340
rect 248328 48331 248380 48340
rect 248328 48297 248337 48331
rect 248337 48297 248371 48331
rect 248371 48297 248380 48331
rect 248328 48288 248380 48297
rect 279884 48331 279936 48340
rect 279884 48297 279893 48331
rect 279893 48297 279927 48331
rect 279927 48297 279936 48331
rect 279884 48288 279936 48297
rect 301872 48288 301924 48340
rect 322664 48331 322716 48340
rect 322664 48297 322673 48331
rect 322673 48297 322707 48331
rect 322707 48297 322716 48331
rect 322664 48288 322716 48297
rect 383292 48288 383344 48340
rect 388812 48288 388864 48340
rect 394424 48288 394476 48340
rect 394516 48288 394568 48340
rect 404084 48288 404136 48340
rect 73620 48220 73672 48272
rect 358084 48220 358136 48272
rect 178224 47608 178276 47660
rect 178408 47608 178460 47660
rect 207112 46996 207164 47048
rect 207204 46928 207256 46980
rect 209872 46971 209924 46980
rect 209872 46937 209881 46971
rect 209881 46937 209915 46971
rect 209915 46937 209924 46971
rect 209872 46928 209924 46937
rect 211252 46971 211304 46980
rect 211252 46937 211261 46971
rect 211261 46937 211295 46971
rect 211295 46937 211304 46971
rect 211252 46928 211304 46937
rect 234712 46971 234764 46980
rect 234712 46937 234721 46971
rect 234721 46937 234755 46971
rect 234755 46937 234764 46971
rect 234712 46928 234764 46937
rect 248328 46971 248380 46980
rect 248328 46937 248337 46971
rect 248337 46937 248371 46971
rect 248371 46937 248380 46971
rect 248328 46928 248380 46937
rect 157432 46860 157484 46912
rect 190828 46860 190880 46912
rect 194968 46860 195020 46912
rect 276112 46903 276164 46912
rect 276112 46869 276121 46903
rect 276121 46869 276155 46903
rect 276155 46869 276164 46903
rect 276112 46860 276164 46869
rect 325700 46903 325752 46912
rect 325700 46869 325709 46903
rect 325709 46869 325743 46903
rect 325743 46869 325752 46903
rect 325700 46860 325752 46869
rect 420460 46860 420512 46912
rect 420644 46860 420696 46912
rect 425980 46903 426032 46912
rect 425980 46869 425989 46903
rect 425989 46869 426023 46903
rect 426023 46869 426032 46903
rect 425980 46860 426032 46869
rect 431592 46903 431644 46912
rect 431592 46869 431601 46903
rect 431601 46869 431635 46903
rect 431635 46869 431644 46903
rect 431592 46860 431644 46869
rect 238852 45883 238904 45892
rect 238852 45849 238861 45883
rect 238861 45849 238895 45883
rect 238895 45849 238904 45883
rect 238852 45840 238904 45849
rect 211252 45611 211304 45620
rect 211252 45577 211261 45611
rect 211261 45577 211295 45611
rect 211295 45577 211304 45611
rect 211252 45568 211304 45577
rect 341524 45611 341576 45620
rect 341524 45577 341533 45611
rect 341533 45577 341567 45611
rect 341567 45577 341576 45611
rect 341524 45568 341576 45577
rect 207204 45543 207256 45552
rect 207204 45509 207213 45543
rect 207213 45509 207247 45543
rect 207247 45509 207256 45543
rect 207204 45500 207256 45509
rect 414940 45543 414992 45552
rect 414940 45509 414949 45543
rect 414949 45509 414983 45543
rect 414983 45509 414992 45543
rect 414940 45500 414992 45509
rect 341524 45432 341576 45484
rect 181168 44115 181220 44124
rect 181168 44081 181177 44115
rect 181177 44081 181211 44115
rect 181211 44081 181220 44115
rect 181168 44072 181220 44081
rect 147864 42032 147916 42084
rect 148140 42032 148192 42084
rect 243452 41828 243504 41880
rect 243820 41828 243872 41880
rect 150808 41463 150860 41472
rect 150808 41429 150817 41463
rect 150817 41429 150851 41463
rect 150851 41429 150860 41463
rect 150808 41420 150860 41429
rect 133604 41352 133656 41404
rect 580172 41352 580224 41404
rect 238944 41284 238996 41336
rect 211344 40672 211396 40724
rect 211528 40672 211580 40724
rect 173900 39312 173952 39364
rect 174084 39312 174136 39364
rect 212632 38632 212684 38684
rect 212724 38632 212776 38684
rect 216680 38632 216732 38684
rect 216772 38632 216824 38684
rect 220912 38632 220964 38684
rect 221096 38632 221148 38684
rect 244280 38632 244332 38684
rect 244372 38632 244424 38684
rect 245752 38632 245804 38684
rect 245844 38632 245896 38684
rect 357992 38675 358044 38684
rect 357992 38641 358001 38675
rect 358001 38641 358035 38675
rect 358035 38641 358044 38675
rect 357992 38632 358044 38641
rect 129004 38564 129056 38616
rect 133236 38564 133288 38616
rect 150808 38607 150860 38616
rect 150808 38573 150817 38607
rect 150817 38573 150851 38607
rect 150851 38573 150860 38607
rect 150808 38564 150860 38573
rect 200488 38564 200540 38616
rect 322756 38564 322808 38616
rect 383200 38607 383252 38616
rect 383200 38573 383209 38607
rect 383209 38573 383243 38607
rect 383243 38573 383252 38607
rect 383200 38564 383252 38573
rect 403992 38607 404044 38616
rect 403992 38573 404001 38607
rect 404001 38573 404035 38607
rect 404035 38573 404044 38607
rect 403992 38564 404044 38573
rect 341432 38267 341484 38276
rect 341432 38233 341441 38267
rect 341441 38233 341475 38267
rect 341475 38233 341484 38267
rect 341432 38224 341484 38233
rect 157340 37315 157392 37324
rect 157340 37281 157349 37315
rect 157349 37281 157383 37315
rect 157383 37281 157392 37315
rect 157340 37272 157392 37281
rect 194692 37315 194744 37324
rect 194692 37281 194701 37315
rect 194701 37281 194735 37315
rect 194735 37281 194744 37315
rect 194692 37272 194744 37281
rect 276112 37315 276164 37324
rect 276112 37281 276121 37315
rect 276121 37281 276155 37315
rect 276155 37281 276164 37315
rect 276112 37272 276164 37281
rect 426072 37272 426124 37324
rect 431592 37315 431644 37324
rect 431592 37281 431601 37315
rect 431601 37281 431635 37315
rect 431635 37281 431644 37315
rect 431592 37272 431644 37281
rect 150808 37204 150860 37256
rect 234712 37247 234764 37256
rect 234712 37213 234721 37247
rect 234721 37213 234755 37247
rect 234755 37213 234764 37247
rect 234712 37204 234764 37213
rect 238944 37204 238996 37256
rect 244280 37247 244332 37256
rect 244280 37213 244289 37247
rect 244289 37213 244323 37247
rect 244323 37213 244332 37247
rect 244280 37204 244332 37213
rect 245752 37247 245804 37256
rect 245752 37213 245761 37247
rect 245761 37213 245795 37247
rect 245795 37213 245804 37247
rect 245752 37204 245804 37213
rect 248328 37247 248380 37256
rect 248328 37213 248337 37247
rect 248337 37213 248371 37247
rect 248371 37213 248380 37247
rect 248328 37204 248380 37213
rect 271880 37247 271932 37256
rect 271880 37213 271889 37247
rect 271889 37213 271923 37247
rect 271923 37213 271932 37247
rect 271880 37204 271932 37213
rect 431592 37179 431644 37188
rect 431592 37145 431601 37179
rect 431601 37145 431635 37179
rect 431635 37145 431644 37179
rect 431592 37136 431644 37145
rect 207204 35955 207256 35964
rect 207204 35921 207213 35955
rect 207213 35921 207247 35955
rect 207247 35921 207256 35955
rect 207204 35912 207256 35921
rect 415032 35912 415084 35964
rect 3424 35844 3476 35896
rect 436192 35844 436244 35896
rect 73804 35343 73856 35352
rect 73804 35309 73813 35343
rect 73813 35309 73847 35343
rect 73847 35309 73856 35343
rect 73804 35300 73856 35309
rect 229192 31875 229244 31884
rect 229192 31841 229201 31875
rect 229201 31841 229235 31875
rect 229235 31841 229244 31875
rect 229192 31832 229244 31841
rect 301964 31832 302016 31884
rect 145012 31764 145064 31816
rect 145196 31764 145248 31816
rect 178224 31696 178276 31748
rect 178408 31696 178460 31748
rect 245844 31696 245896 31748
rect 279884 31696 279936 31748
rect 280068 31696 280120 31748
rect 302056 31696 302108 31748
rect 388720 31696 388772 31748
rect 388904 31696 388956 31748
rect 181168 31671 181220 31680
rect 181168 31637 181177 31671
rect 181177 31637 181211 31671
rect 181211 31637 181220 31671
rect 181168 31628 181220 31637
rect 244372 31628 244424 31680
rect 341432 31628 341484 31680
rect 341524 31628 341576 31680
rect 431684 31628 431736 31680
rect 133144 31059 133196 31068
rect 133144 31025 133153 31059
rect 133153 31025 133187 31059
rect 133187 31025 133196 31059
rect 133144 31016 133196 31025
rect 132408 30268 132460 30320
rect 580172 30268 580224 30320
rect 325700 29087 325752 29096
rect 325700 29053 325709 29087
rect 325709 29053 325743 29087
rect 325743 29053 325752 29087
rect 325700 29044 325752 29053
rect 357992 29044 358044 29096
rect 128912 29019 128964 29028
rect 128912 28985 128921 29019
rect 128921 28985 128955 29019
rect 128955 28985 128964 29019
rect 128912 28976 128964 28985
rect 157340 28976 157392 29028
rect 157432 28976 157484 29028
rect 159088 28976 159140 29028
rect 159272 28976 159324 29028
rect 190736 29019 190788 29028
rect 190736 28985 190745 29019
rect 190745 28985 190779 29019
rect 190779 28985 190788 29019
rect 190736 28976 190788 28985
rect 200396 29019 200448 29028
rect 200396 28985 200405 29019
rect 200405 28985 200439 29019
rect 200439 28985 200448 29019
rect 200396 28976 200448 28985
rect 229192 29019 229244 29028
rect 229192 28985 229201 29019
rect 229201 28985 229235 29019
rect 229235 28985 229244 29019
rect 229192 28976 229244 28985
rect 322664 29019 322716 29028
rect 322664 28985 322673 29019
rect 322673 28985 322707 29019
rect 322707 28985 322716 29019
rect 322664 28976 322716 28985
rect 383292 28976 383344 29028
rect 394424 28976 394476 29028
rect 394516 28976 394568 29028
rect 404084 28976 404136 29028
rect 183744 28908 183796 28960
rect 185032 28908 185084 28960
rect 207204 28908 207256 28960
rect 207296 28908 207348 28960
rect 280068 28908 280120 28960
rect 183744 28772 183796 28824
rect 388720 28772 388772 28824
rect 388904 28772 388956 28824
rect 150716 27659 150768 27668
rect 150716 27625 150725 27659
rect 150725 27625 150759 27659
rect 150759 27625 150768 27659
rect 150716 27616 150768 27625
rect 211160 27616 211212 27668
rect 211344 27616 211396 27668
rect 234712 27659 234764 27668
rect 234712 27625 234721 27659
rect 234721 27625 234755 27659
rect 234755 27625 234764 27659
rect 234712 27616 234764 27625
rect 238852 27659 238904 27668
rect 238852 27625 238861 27659
rect 238861 27625 238895 27659
rect 238895 27625 238904 27659
rect 238852 27616 238904 27625
rect 243728 27659 243780 27668
rect 243728 27625 243737 27659
rect 243737 27625 243771 27659
rect 243771 27625 243780 27659
rect 243728 27616 243780 27625
rect 248328 27659 248380 27668
rect 248328 27625 248337 27659
rect 248337 27625 248371 27659
rect 248371 27625 248380 27659
rect 248328 27616 248380 27625
rect 272156 27616 272208 27668
rect 157432 27548 157484 27600
rect 276112 27591 276164 27600
rect 276112 27557 276121 27591
rect 276121 27557 276155 27591
rect 276155 27557 276164 27591
rect 276112 27548 276164 27557
rect 325700 27591 325752 27600
rect 325700 27557 325709 27591
rect 325709 27557 325743 27591
rect 325743 27557 325752 27591
rect 325700 27548 325752 27557
rect 420460 27591 420512 27600
rect 420460 27557 420469 27591
rect 420469 27557 420503 27591
rect 420503 27557 420512 27591
rect 420460 27548 420512 27557
rect 357716 26367 357768 26376
rect 357716 26333 357725 26367
rect 357725 26333 357759 26367
rect 357759 26333 357768 26367
rect 357716 26324 357768 26333
rect 175556 26299 175608 26308
rect 175556 26265 175565 26299
rect 175565 26265 175599 26299
rect 175599 26265 175608 26299
rect 175556 26256 175608 26265
rect 179420 26256 179472 26308
rect 179512 26256 179564 26308
rect 243728 26299 243780 26308
rect 243728 26265 243737 26299
rect 243737 26265 243771 26299
rect 243771 26265 243780 26299
rect 243728 26256 243780 26265
rect 301872 26231 301924 26240
rect 301872 26197 301881 26231
rect 301881 26197 301915 26231
rect 301915 26197 301924 26231
rect 301872 26188 301924 26197
rect 357716 26188 357768 26240
rect 415032 26231 415084 26240
rect 415032 26197 415041 26231
rect 415041 26197 415075 26231
rect 415075 26197 415084 26231
rect 415032 26188 415084 26197
rect 431684 26188 431736 26240
rect 383384 25279 383436 25288
rect 383384 25245 383393 25279
rect 383393 25245 383427 25279
rect 383427 25245 383436 25279
rect 383384 25236 383436 25245
rect 178040 25075 178092 25084
rect 178040 25041 178049 25075
rect 178049 25041 178083 25075
rect 178083 25041 178092 25075
rect 178040 25032 178092 25041
rect 73620 24828 73672 24880
rect 73896 24828 73948 24880
rect 175556 24871 175608 24880
rect 175556 24837 175565 24871
rect 175565 24837 175599 24871
rect 175599 24837 175608 24871
rect 175556 24828 175608 24837
rect 179512 24760 179564 24812
rect 178040 24735 178092 24744
rect 178040 24701 178049 24735
rect 178049 24701 178083 24735
rect 178083 24701 178092 24735
rect 178040 24692 178092 24701
rect 147864 24148 147916 24200
rect 148048 24148 148100 24200
rect 220912 24148 220964 24200
rect 221096 24148 221148 24200
rect 234712 22788 234764 22840
rect 394516 22244 394568 22296
rect 205916 22176 205968 22228
rect 394424 22176 394476 22228
rect 181168 22108 181220 22160
rect 212724 22108 212776 22160
rect 233332 22151 233384 22160
rect 233332 22117 233341 22151
rect 233341 22117 233375 22151
rect 233375 22117 233384 22151
rect 233332 22108 233384 22117
rect 243728 22108 243780 22160
rect 3148 22040 3200 22092
rect 132224 22040 132276 22092
rect 181076 22040 181128 22092
rect 200212 22040 200264 22092
rect 200396 22040 200448 22092
rect 214104 22040 214156 22092
rect 212724 21972 212776 22024
rect 404084 22108 404136 22160
rect 244372 22040 244424 22092
rect 244556 22040 244608 22092
rect 245844 22040 245896 22092
rect 246028 22040 246080 22092
rect 403992 22040 404044 22092
rect 214196 21972 214248 22024
rect 243728 21972 243780 22024
rect 357900 22015 357952 22024
rect 357900 21981 357909 22015
rect 357909 21981 357943 22015
rect 357943 21981 357952 22015
rect 357900 21972 357952 21981
rect 73896 20000 73948 20052
rect 173900 20000 173952 20052
rect 190736 19388 190788 19440
rect 159088 19320 159140 19372
rect 159272 19320 159324 19372
rect 162952 19320 163004 19372
rect 163136 19320 163188 19372
rect 184940 19363 184992 19372
rect 184940 19329 184949 19363
rect 184949 19329 184983 19363
rect 184983 19329 184992 19363
rect 184940 19320 184992 19329
rect 205732 19363 205784 19372
rect 205732 19329 205741 19363
rect 205741 19329 205775 19363
rect 205775 19329 205784 19363
rect 205732 19320 205784 19329
rect 211160 19320 211212 19372
rect 211344 19320 211396 19372
rect 216680 19320 216732 19372
rect 216956 19320 217008 19372
rect 229100 19320 229152 19372
rect 229284 19320 229336 19372
rect 279976 19363 280028 19372
rect 279976 19329 279985 19363
rect 279985 19329 280019 19363
rect 280019 19329 280028 19363
rect 279976 19320 280028 19329
rect 383384 19363 383436 19372
rect 383384 19329 383393 19363
rect 383393 19329 383427 19363
rect 383427 19329 383436 19363
rect 383384 19320 383436 19329
rect 143632 19295 143684 19304
rect 143632 19261 143641 19295
rect 143641 19261 143675 19295
rect 143675 19261 143684 19295
rect 143632 19252 143684 19261
rect 200396 19295 200448 19304
rect 200396 19261 200405 19295
rect 200405 19261 200439 19295
rect 200439 19261 200448 19295
rect 200396 19252 200448 19261
rect 233332 19295 233384 19304
rect 233332 19261 233341 19295
rect 233341 19261 233375 19295
rect 233375 19261 233384 19295
rect 233332 19252 233384 19261
rect 244556 19295 244608 19304
rect 244556 19261 244565 19295
rect 244565 19261 244599 19295
rect 244599 19261 244608 19295
rect 244556 19252 244608 19261
rect 394332 19295 394384 19304
rect 394332 19261 394341 19295
rect 394341 19261 394375 19295
rect 394375 19261 394384 19295
rect 394332 19252 394384 19261
rect 425980 19252 426032 19304
rect 426072 19252 426124 19304
rect 274824 18139 274876 18148
rect 274824 18105 274833 18139
rect 274833 18105 274867 18139
rect 274867 18105 274876 18139
rect 274824 18096 274876 18105
rect 190644 18003 190696 18012
rect 190644 17969 190653 18003
rect 190653 17969 190687 18003
rect 190687 17969 190696 18003
rect 190644 17960 190696 17969
rect 234620 18003 234672 18012
rect 234620 17969 234629 18003
rect 234629 17969 234663 18003
rect 234663 17969 234672 18003
rect 234620 17960 234672 17969
rect 276112 18003 276164 18012
rect 276112 17969 276121 18003
rect 276121 17969 276155 18003
rect 276155 17969 276164 18003
rect 276112 17960 276164 17969
rect 420552 17960 420604 18012
rect 436744 17892 436796 17944
rect 579804 17892 579856 17944
rect 415032 16643 415084 16652
rect 415032 16609 415041 16643
rect 415041 16609 415075 16643
rect 415075 16609 415084 16643
rect 415032 16600 415084 16609
rect 431500 16643 431552 16652
rect 431500 16609 431509 16643
rect 431509 16609 431543 16643
rect 431543 16609 431552 16643
rect 431500 16600 431552 16609
rect 383292 12563 383344 12572
rect 383292 12529 383301 12563
rect 383301 12529 383335 12563
rect 383335 12529 383344 12563
rect 383292 12520 383344 12529
rect 168472 12452 168524 12504
rect 183744 12452 183796 12504
rect 211344 12452 211396 12504
rect 276112 12452 276164 12504
rect 183652 12384 183704 12436
rect 211252 12384 211304 12436
rect 74264 12359 74316 12368
rect 74264 12325 74273 12359
rect 74273 12325 74307 12359
rect 74307 12325 74316 12359
rect 74264 12316 74316 12325
rect 178132 12359 178184 12368
rect 178132 12325 178141 12359
rect 178141 12325 178175 12359
rect 178175 12325 178184 12359
rect 178132 12316 178184 12325
rect 415032 12452 415084 12504
rect 420552 12452 420604 12504
rect 280344 12384 280396 12436
rect 281264 12384 281316 12436
rect 321744 12384 321796 12436
rect 414940 12384 414992 12436
rect 420460 12384 420512 12436
rect 463700 12384 463752 12436
rect 464344 12384 464396 12436
rect 276480 12316 276532 12368
rect 322756 12316 322808 12368
rect 200396 12291 200448 12300
rect 200396 12257 200405 12291
rect 200405 12257 200439 12291
rect 200439 12257 200448 12291
rect 200396 12248 200448 12257
rect 205548 12112 205600 12164
rect 205732 12112 205784 12164
rect 246028 11908 246080 11960
rect 244556 11883 244608 11892
rect 244556 11849 244565 11883
rect 244565 11849 244599 11883
rect 244599 11849 244608 11883
rect 244556 11840 244608 11849
rect 246028 11772 246080 11824
rect 371056 10684 371108 10736
rect 459652 10684 459704 10736
rect 372344 10616 372396 10668
rect 463240 10616 463292 10668
rect 375196 10548 375248 10600
rect 466828 10548 466880 10600
rect 376576 10480 376628 10532
rect 470324 10480 470376 10532
rect 377956 10412 378008 10464
rect 473360 10412 473412 10464
rect 380808 10344 380860 10396
rect 477592 10344 477644 10396
rect 382096 10276 382148 10328
rect 481088 10276 481140 10328
rect 143724 9664 143776 9716
rect 157340 9707 157392 9716
rect 157340 9673 157349 9707
rect 157349 9673 157383 9707
rect 157383 9673 157392 9707
rect 157340 9664 157392 9673
rect 168380 9707 168432 9716
rect 168380 9673 168389 9707
rect 168389 9673 168423 9707
rect 168423 9673 168432 9707
rect 168380 9664 168432 9673
rect 190644 9664 190696 9716
rect 190736 9664 190788 9716
rect 228916 9664 228968 9716
rect 229192 9664 229244 9716
rect 234620 9664 234672 9716
rect 234712 9664 234764 9716
rect 275284 9664 275336 9716
rect 326252 9664 326304 9716
rect 383292 9707 383344 9716
rect 383292 9673 383301 9707
rect 383301 9673 383335 9707
rect 383335 9673 383344 9707
rect 383292 9664 383344 9673
rect 394424 9664 394476 9716
rect 87328 9596 87380 9648
rect 183652 9639 183704 9648
rect 183652 9605 183661 9639
rect 183661 9605 183695 9639
rect 183695 9605 183704 9639
rect 183652 9596 183704 9605
rect 368388 9596 368440 9648
rect 454868 9596 454920 9648
rect 75460 9528 75512 9580
rect 371148 9528 371200 9580
rect 458456 9528 458508 9580
rect 68284 9460 68336 9512
rect 168380 9460 168432 9512
rect 183560 9503 183612 9512
rect 183560 9469 183569 9503
rect 183569 9469 183603 9503
rect 183603 9469 183612 9503
rect 183560 9460 183612 9469
rect 372436 9460 372488 9512
rect 462044 9460 462096 9512
rect 61200 9392 61252 9444
rect 164424 9392 164476 9444
rect 172612 9392 172664 9444
rect 419448 9392 419500 9444
rect 552388 9392 552440 9444
rect 55220 9324 55272 9376
rect 161480 9324 161532 9376
rect 420460 9324 420512 9376
rect 555976 9324 556028 9376
rect 58808 9256 58860 9308
rect 164332 9256 164384 9308
rect 422116 9256 422168 9308
rect 559564 9256 559616 9308
rect 54024 9188 54076 9240
rect 161572 9188 161624 9240
rect 409512 9188 409564 9240
rect 409788 9188 409840 9240
rect 424968 9188 425020 9240
rect 563152 9188 563204 9240
rect 46940 9120 46992 9172
rect 157340 9120 157392 9172
rect 350356 9120 350408 9172
rect 420368 9120 420420 9172
rect 425980 9120 426032 9172
rect 566740 9120 566792 9172
rect 40960 9052 41012 9104
rect 154672 9052 154724 9104
rect 353208 9052 353260 9104
rect 423956 9052 424008 9104
rect 427636 9052 427688 9104
rect 570236 9052 570288 9104
rect 26700 8984 26752 9036
rect 147772 8984 147824 9036
rect 354496 8984 354548 9036
rect 427544 8984 427596 9036
rect 431500 8984 431552 9036
rect 577412 8984 577464 9036
rect 6460 8916 6512 8968
rect 136824 8916 136876 8968
rect 355876 8916 355928 8968
rect 431132 8916 431184 8968
rect 433156 8916 433208 8968
rect 581000 8916 581052 8968
rect 106372 8848 106424 8900
rect 187792 8848 187844 8900
rect 369768 8848 369820 8900
rect 456064 8848 456116 8900
rect 119436 8780 119488 8832
rect 194784 8780 194836 8832
rect 366916 8780 366968 8832
rect 452476 8780 452528 8832
rect 120632 8712 120684 8764
rect 190552 8712 190604 8764
rect 365536 8712 365588 8764
rect 448980 8712 449032 8764
rect 361396 8644 361448 8696
rect 441804 8644 441856 8696
rect 364248 8576 364300 8628
rect 445392 8576 445444 8628
rect 360016 8508 360068 8560
rect 438216 8508 438268 8560
rect 358636 8440 358688 8492
rect 434628 8440 434680 8492
rect 247960 8304 248012 8356
rect 248328 8304 248380 8356
rect 302056 8304 302108 8356
rect 357808 8304 357860 8356
rect 357900 8304 357952 8356
rect 3424 8236 3476 8288
rect 131764 8236 131816 8288
rect 133788 8236 133840 8288
rect 203064 8236 203116 8288
rect 384948 8236 385000 8288
rect 486976 8236 487028 8288
rect 34980 8168 35032 8220
rect 127624 8168 127676 8220
rect 127808 8168 127860 8220
rect 198740 8168 198792 8220
rect 387616 8168 387668 8220
rect 490564 8168 490616 8220
rect 51632 8100 51684 8152
rect 160192 8100 160244 8152
rect 388904 8100 388956 8152
rect 494152 8100 494204 8152
rect 48136 8032 48188 8084
rect 158812 8032 158864 8084
rect 390468 8032 390520 8084
rect 497740 8032 497792 8084
rect 20720 7964 20772 8016
rect 143724 7964 143776 8016
rect 144460 7964 144512 8016
rect 208492 7964 208544 8016
rect 393136 7964 393188 8016
rect 501236 7964 501288 8016
rect 13636 7896 13688 7948
rect 140872 7896 140924 7948
rect 143264 7896 143316 7948
rect 207204 7896 207256 7948
rect 394332 7896 394384 7948
rect 504824 7896 504876 7948
rect 7656 7828 7708 7880
rect 136732 7828 136784 7880
rect 140964 7828 141016 7880
rect 205548 7828 205600 7880
rect 395896 7828 395948 7880
rect 508412 7828 508464 7880
rect 1676 7760 1728 7812
rect 133880 7760 133932 7812
rect 136088 7760 136140 7812
rect 202880 7760 202932 7812
rect 413928 7760 413980 7812
rect 541716 7760 541768 7812
rect 5264 7692 5316 7744
rect 136640 7692 136692 7744
rect 139676 7692 139728 7744
rect 205640 7692 205692 7744
rect 344744 7692 344796 7744
rect 409696 7692 409748 7744
rect 414940 7692 414992 7744
rect 545304 7692 545356 7744
rect 2872 7624 2924 7676
rect 135352 7624 135404 7676
rect 137284 7624 137336 7676
rect 204352 7624 204404 7676
rect 347688 7624 347740 7676
rect 413284 7624 413336 7676
rect 416596 7624 416648 7676
rect 548892 7624 548944 7676
rect 572 7556 624 7608
rect 134156 7556 134208 7608
rect 134892 7556 134944 7608
rect 202972 7556 203024 7608
rect 348976 7556 349028 7608
rect 416780 7556 416832 7608
rect 417976 7556 418028 7608
rect 430488 7556 430540 7608
rect 573824 7556 573876 7608
rect 115940 7488 115992 7540
rect 117136 7488 117188 7540
rect 118240 7488 118292 7540
rect 194600 7488 194652 7540
rect 383292 7488 383344 7540
rect 121828 7420 121880 7472
rect 196072 7420 196124 7472
rect 367008 7420 367060 7472
rect 451280 7420 451332 7472
rect 477500 7488 477552 7540
rect 478696 7488 478748 7540
rect 483480 7420 483532 7472
rect 126612 7352 126664 7404
rect 198832 7352 198884 7404
rect 365628 7352 365680 7404
rect 447784 7352 447836 7404
rect 77852 7284 77904 7336
rect 84936 7216 84988 7268
rect 129004 7284 129056 7336
rect 200120 7284 200172 7336
rect 362868 7284 362920 7336
rect 444196 7284 444248 7336
rect 95700 7148 95752 7200
rect 129096 7216 129148 7268
rect 130200 7216 130252 7268
rect 200396 7216 200448 7268
rect 361488 7216 361540 7268
rect 440608 7216 440660 7268
rect 129188 7148 129240 7200
rect 131396 7148 131448 7200
rect 201592 7148 201644 7200
rect 358728 7148 358780 7200
rect 435824 7148 435876 7200
rect 109960 7080 110012 7132
rect 133052 7080 133104 7132
rect 133144 7080 133196 7132
rect 201500 7080 201552 7132
rect 360108 7080 360160 7132
rect 437020 7080 437072 7132
rect 129280 7012 129332 7064
rect 416872 7012 416924 7064
rect 173992 6919 174044 6928
rect 173992 6885 174001 6919
rect 174001 6885 174035 6919
rect 174035 6885 174044 6919
rect 173992 6876 174044 6885
rect 179420 6919 179472 6928
rect 179420 6885 179429 6919
rect 179429 6885 179463 6919
rect 179463 6885 179472 6919
rect 179420 6876 179472 6885
rect 96896 6808 96948 6860
rect 317144 6808 317196 6860
rect 356152 6808 356204 6860
rect 391756 6808 391808 6860
rect 498936 6808 498988 6860
rect 94504 6740 94556 6792
rect 182272 6740 182324 6792
rect 326896 6740 326948 6792
rect 374000 6740 374052 6792
rect 393228 6740 393280 6792
rect 502432 6740 502484 6792
rect 89720 6672 89772 6724
rect 179420 6672 179472 6724
rect 328184 6672 328236 6724
rect 377588 6672 377640 6724
rect 394608 6672 394660 6724
rect 506020 6672 506072 6724
rect 90916 6604 90968 6656
rect 180892 6604 180944 6656
rect 331036 6604 331088 6656
rect 381176 6604 381228 6656
rect 397368 6604 397420 6656
rect 509608 6604 509660 6656
rect 86132 6536 86184 6588
rect 178040 6536 178092 6588
rect 332416 6536 332468 6588
rect 384672 6536 384724 6588
rect 398656 6536 398708 6588
rect 513196 6536 513248 6588
rect 79048 6468 79100 6520
rect 173992 6468 174044 6520
rect 336648 6468 336700 6520
rect 391848 6468 391900 6520
rect 399944 6468 399996 6520
rect 516784 6468 516836 6520
rect 71872 6400 71924 6452
rect 169852 6400 169904 6452
rect 333704 6400 333756 6452
rect 388260 6400 388312 6452
rect 402796 6400 402848 6452
rect 520280 6400 520332 6452
rect 64788 6332 64840 6384
rect 167092 6332 167144 6384
rect 337936 6332 337988 6384
rect 395436 6332 395488 6384
rect 404176 6332 404228 6384
rect 523868 6332 523920 6384
rect 57612 6264 57664 6316
rect 162860 6264 162912 6316
rect 177488 6264 177540 6316
rect 214196 6264 214248 6316
rect 342168 6264 342220 6316
rect 402520 6264 402572 6316
rect 408408 6264 408460 6316
rect 531044 6264 531096 6316
rect 36176 6196 36228 6248
rect 151820 6196 151872 6248
rect 183560 6196 183612 6248
rect 222292 6196 222344 6248
rect 339316 6196 339368 6248
rect 399024 6196 399076 6248
rect 405556 6196 405608 6248
rect 527456 6196 527508 6248
rect 29092 6128 29144 6180
rect 148048 6128 148100 6180
rect 153936 6128 153988 6180
rect 212724 6128 212776 6180
rect 343456 6128 343508 6180
rect 406108 6128 406160 6180
rect 409604 6128 409656 6180
rect 534540 6128 534592 6180
rect 98092 6060 98144 6112
rect 318708 6060 318760 6112
rect 358544 6060 358596 6112
rect 388996 6060 389048 6112
rect 495348 6060 495400 6112
rect 101588 5992 101640 6044
rect 186320 5992 186372 6044
rect 317236 5992 317288 6044
rect 354956 5992 355008 6044
rect 387708 5992 387760 6044
rect 491760 5992 491812 6044
rect 103980 5924 104032 5976
rect 186504 5924 186556 5976
rect 315948 5924 316000 5976
rect 352564 5924 352616 5976
rect 383476 5924 383528 5976
rect 484584 5924 484636 5976
rect 105176 5856 105228 5908
rect 187700 5856 187752 5908
rect 315856 5856 315908 5908
rect 351368 5856 351420 5908
rect 386328 5856 386380 5908
rect 488172 5856 488224 5908
rect 56416 5788 56468 5840
rect 108304 5788 108356 5840
rect 108764 5788 108816 5840
rect 189172 5788 189224 5840
rect 379336 5788 379388 5840
rect 476304 5788 476356 5840
rect 112352 5720 112404 5772
rect 191932 5720 191984 5772
rect 382188 5720 382240 5772
rect 479892 5720 479944 5772
rect 111156 5652 111208 5704
rect 190552 5652 190604 5704
rect 378048 5652 378100 5704
rect 472716 5652 472768 5704
rect 115940 5584 115992 5636
rect 193220 5584 193272 5636
rect 373908 5584 373960 5636
rect 465632 5584 465684 5636
rect 123024 5516 123076 5568
rect 197452 5516 197504 5568
rect 376668 5516 376720 5568
rect 469128 5516 469180 5568
rect 69480 5448 69532 5500
rect 169944 5448 169996 5500
rect 174176 5448 174228 5500
rect 223672 5448 223724 5500
rect 335176 5448 335228 5500
rect 390652 5448 390704 5500
rect 415308 5448 415360 5500
rect 544108 5448 544160 5500
rect 65984 5380 66036 5432
rect 167000 5380 167052 5432
rect 170588 5380 170640 5432
rect 221096 5380 221148 5432
rect 339408 5380 339460 5432
rect 397828 5380 397880 5432
rect 416688 5380 416740 5432
rect 547696 5380 547748 5432
rect 62396 5312 62448 5364
rect 165712 5312 165764 5364
rect 167092 5312 167144 5364
rect 219532 5312 219584 5364
rect 340696 5312 340748 5364
rect 401324 5312 401376 5364
rect 418068 5312 418120 5364
rect 551192 5312 551244 5364
rect 44548 5244 44600 5296
rect 156236 5244 156288 5296
rect 158720 5244 158772 5296
rect 215392 5244 215444 5296
rect 343548 5244 343600 5296
rect 404912 5244 404964 5296
rect 420828 5244 420880 5296
rect 554780 5244 554832 5296
rect 37372 5176 37424 5228
rect 153292 5176 153344 5228
rect 156328 5176 156380 5228
rect 213920 5176 213972 5228
rect 344836 5176 344888 5228
rect 408684 5176 408736 5228
rect 422208 5176 422260 5228
rect 558368 5176 558420 5228
rect 33876 5108 33928 5160
rect 150716 5108 150768 5160
rect 155132 5108 155184 5160
rect 214012 5108 214064 5160
rect 346308 5108 346360 5160
rect 412088 5108 412140 5160
rect 423588 5108 423640 5160
rect 561956 5108 562008 5160
rect 18328 5040 18380 5092
rect 135444 5040 135496 5092
rect 138480 5040 138532 5092
rect 204260 5040 204312 5092
rect 204352 5040 204404 5092
rect 237472 5040 237524 5092
rect 349068 5040 349120 5092
rect 415676 5040 415728 5092
rect 426348 5040 426400 5092
rect 565544 5040 565596 5092
rect 21916 4972 21968 5024
rect 145104 4972 145156 5024
rect 152740 4972 152792 5024
rect 212540 4972 212592 5024
rect 350448 4972 350500 5024
rect 419172 4972 419224 5024
rect 427728 4972 427780 5024
rect 569040 4972 569092 5024
rect 17224 4904 17276 4956
rect 142252 4904 142304 4956
rect 149244 4904 149296 4956
rect 209872 4904 209924 4956
rect 215852 4904 215904 4956
rect 244556 4904 244608 4956
rect 310428 4904 310480 4956
rect 341892 4904 341944 4956
rect 354588 4904 354640 4956
rect 426348 4904 426400 4956
rect 429108 4904 429160 4956
rect 572628 4904 572680 4956
rect 12440 4836 12492 4888
rect 139492 4836 139544 4888
rect 145656 4836 145708 4888
rect 208584 4836 208636 4888
rect 212264 4836 212316 4888
rect 242992 4836 243044 4888
rect 314568 4836 314620 4888
rect 349068 4836 349120 4888
rect 351736 4836 351788 4888
rect 422760 4836 422812 4888
rect 431868 4836 431920 4888
rect 576216 4836 576268 4888
rect 4068 4768 4120 4820
rect 135260 4768 135312 4820
rect 142068 4768 142120 4820
rect 207020 4768 207072 4820
rect 208216 4768 208268 4820
rect 238944 4768 238996 4820
rect 313096 4768 313148 4820
rect 347872 4768 347924 4820
rect 355968 4768 356020 4820
rect 429936 4768 429988 4820
rect 433248 4768 433300 4820
rect 579804 4768 579856 4820
rect 73068 4700 73120 4752
rect 171232 4700 171284 4752
rect 173900 4700 173952 4752
rect 211252 4700 211304 4752
rect 338028 4700 338080 4752
rect 394240 4700 394292 4752
rect 412548 4700 412600 4752
rect 540520 4700 540572 4752
rect 76656 4632 76708 4684
rect 172520 4632 172572 4684
rect 208676 4632 208728 4684
rect 240140 4632 240192 4684
rect 333796 4632 333848 4684
rect 387064 4632 387116 4684
rect 411168 4632 411220 4684
rect 536932 4632 536984 4684
rect 80244 4564 80296 4616
rect 175372 4564 175424 4616
rect 202880 4564 202932 4616
rect 233332 4564 233384 4616
rect 329748 4564 329800 4616
rect 379980 4564 380032 4616
rect 409788 4564 409840 4616
rect 533436 4564 533488 4616
rect 83832 4496 83884 4548
rect 176752 4496 176804 4548
rect 204260 4496 204312 4548
rect 234712 4496 234764 4548
rect 332508 4496 332560 4548
rect 383568 4496 383620 4548
rect 406936 4496 406988 4548
rect 529848 4496 529900 4548
rect 49332 4428 49384 4480
rect 130384 4428 130436 4480
rect 163504 4428 163556 4480
rect 218152 4428 218204 4480
rect 328276 4428 328328 4480
rect 376392 4428 376444 4480
rect 405648 4428 405700 4480
rect 526260 4428 526312 4480
rect 45744 4360 45796 4412
rect 126244 4360 126296 4412
rect 326988 4360 327040 4412
rect 372804 4360 372856 4412
rect 401508 4360 401560 4412
rect 519084 4360 519136 4412
rect 52828 4292 52880 4344
rect 122104 4292 122156 4344
rect 164700 4292 164752 4344
rect 218060 4292 218112 4344
rect 324136 4292 324188 4344
rect 369124 4292 369176 4344
rect 404268 4292 404320 4344
rect 522672 4292 522724 4344
rect 63592 4224 63644 4276
rect 128820 4224 128872 4276
rect 215300 4224 215352 4276
rect 322572 4224 322624 4276
rect 365720 4224 365772 4276
rect 400036 4224 400088 4276
rect 515588 4224 515640 4276
rect 67548 4156 67600 4208
rect 70676 4156 70728 4208
rect 120724 4156 120776 4208
rect 42156 4088 42208 4140
rect 151912 4088 151964 4140
rect 159916 4088 159968 4140
rect 321376 4156 321428 4208
rect 362132 4156 362184 4208
rect 398748 4156 398800 4208
rect 512000 4156 512052 4208
rect 168196 4088 168248 4140
rect 174544 4088 174596 4140
rect 175372 4088 175424 4140
rect 176568 4088 176620 4140
rect 177764 4088 177816 4140
rect 180064 4088 180116 4140
rect 182548 4088 182600 4140
rect 183468 4088 183520 4140
rect 190828 4088 190880 4140
rect 43352 4020 43404 4072
rect 155960 4020 156012 4072
rect 187240 4020 187292 4072
rect 39764 3952 39816 4004
rect 153200 3952 153252 4004
rect 171784 3952 171836 4004
rect 183560 3952 183612 4004
rect 188436 3952 188488 4004
rect 225328 4088 225380 4140
rect 226248 4088 226300 4140
rect 226524 4088 226576 4140
rect 227628 4088 227680 4140
rect 227720 4088 227772 4140
rect 229008 4088 229060 4140
rect 231308 4088 231360 4140
rect 231768 4088 231820 4140
rect 233700 4088 233752 4140
rect 234528 4088 234580 4140
rect 239588 4088 239640 4140
rect 240048 4088 240100 4140
rect 243176 4088 243228 4140
rect 244188 4088 244240 4140
rect 244372 4088 244424 4140
rect 245568 4088 245620 4140
rect 246764 4088 246816 4140
rect 247684 4088 247736 4140
rect 249156 4088 249208 4140
rect 249708 4088 249760 4140
rect 251456 4088 251508 4140
rect 252468 4088 252520 4140
rect 265808 4088 265860 4140
rect 266268 4088 266320 4140
rect 268108 4088 268160 4140
rect 269764 4088 269816 4140
rect 271696 4088 271748 4140
rect 272524 4088 272576 4140
rect 274088 4088 274140 4140
rect 274548 4088 274600 4140
rect 277308 4088 277360 4140
rect 277676 4088 277728 4140
rect 280068 4088 280120 4140
rect 282460 4088 282512 4140
rect 292396 4088 292448 4140
rect 307392 4088 307444 4140
rect 315304 4088 315356 4140
rect 315856 4088 315908 4140
rect 321468 4088 321520 4140
rect 363328 4088 363380 4140
rect 363604 4088 363656 4140
rect 364524 4088 364576 4140
rect 391756 4088 391808 4140
rect 500132 4088 500184 4140
rect 502984 4088 503036 4140
rect 507124 4088 507176 4140
rect 571432 4088 571484 4140
rect 241980 4020 242032 4072
rect 243728 4020 243780 4072
rect 284208 4020 284260 4072
rect 289544 4020 289596 4072
rect 297916 4020 297968 4072
rect 298008 4020 298060 4072
rect 316960 4020 317012 4072
rect 322848 4020 322900 4072
rect 395988 4020 396040 4072
rect 507216 4020 507268 4072
rect 578608 4020 578660 4072
rect 231952 3952 232004 4004
rect 269304 3952 269356 4004
rect 272156 3952 272208 4004
rect 285588 3952 285640 4004
rect 293132 3952 293184 4004
rect 318064 3952 318116 4004
rect 324228 3952 324280 4004
rect 368020 3952 368072 4004
rect 400128 3952 400180 4004
rect 514392 3952 514444 4004
rect 32680 3884 32732 3936
rect 150440 3884 150492 3936
rect 161112 3884 161164 3936
rect 178684 3884 178736 3936
rect 183744 3884 183796 3936
rect 227904 3884 227956 3936
rect 236000 3884 236052 3936
rect 237288 3884 237340 3936
rect 283564 3884 283616 3936
rect 287152 3884 287204 3936
rect 288348 3884 288400 3936
rect 297916 3884 297968 3936
rect 302148 3884 302200 3936
rect 324044 3884 324096 3936
rect 326344 3884 326396 3936
rect 370412 3884 370464 3936
rect 374644 3884 374696 3936
rect 25504 3816 25556 3868
rect 146300 3816 146352 3868
rect 157524 3816 157576 3868
rect 177488 3816 177540 3868
rect 180156 3816 180208 3868
rect 226432 3816 226484 3868
rect 228916 3816 228968 3868
rect 235264 3816 235316 3868
rect 286876 3816 286928 3868
rect 295524 3816 295576 3868
rect 299388 3816 299440 3868
rect 320456 3816 320508 3868
rect 328368 3816 328420 3868
rect 375196 3816 375248 3868
rect 384304 3884 384356 3936
rect 396632 3884 396684 3936
rect 402888 3884 402940 3936
rect 521476 3884 521528 3936
rect 393044 3816 393096 3868
rect 24308 3748 24360 3800
rect 146392 3748 146444 3800
rect 151544 3748 151596 3800
rect 173900 3748 173952 3800
rect 176476 3748 176528 3800
rect 19524 3680 19576 3732
rect 143540 3680 143592 3732
rect 172980 3680 173032 3732
rect 230572 3748 230624 3800
rect 286968 3748 287020 3800
rect 296720 3748 296772 3800
rect 302056 3748 302108 3800
rect 325240 3748 325292 3800
rect 326160 3748 326212 3800
rect 334624 3748 334676 3800
rect 335912 3748 335964 3800
rect 382372 3748 382424 3800
rect 389824 3748 389876 3800
rect 403716 3748 403768 3800
rect 407028 3816 407080 3868
rect 528652 3816 528704 3868
rect 409512 3748 409564 3800
rect 535736 3748 535788 3800
rect 218152 3680 218204 3732
rect 224224 3680 224276 3732
rect 229192 3680 229244 3732
rect 288256 3680 288308 3732
rect 299112 3680 299164 3732
rect 303528 3680 303580 3732
rect 327632 3680 327684 3732
rect 333888 3680 333940 3732
rect 385868 3680 385920 3732
rect 396724 3680 396776 3732
rect 410892 3680 410944 3732
rect 418160 3680 418212 3732
rect 542912 3680 542964 3732
rect 14832 3612 14884 3664
rect 140780 3612 140832 3664
rect 148048 3612 148100 3664
rect 196808 3612 196860 3664
rect 197268 3612 197320 3664
rect 200396 3612 200448 3664
rect 201408 3612 201460 3664
rect 201500 3612 201552 3664
rect 204352 3612 204404 3664
rect 207480 3612 207532 3664
rect 208308 3612 208360 3664
rect 209872 3612 209924 3664
rect 211068 3612 211120 3664
rect 233884 3612 233936 3664
rect 234804 3612 234856 3664
rect 250444 3612 250496 3664
rect 284944 3612 284996 3664
rect 288348 3612 288400 3664
rect 291016 3612 291068 3664
rect 303804 3612 303856 3664
rect 306288 3612 306340 3664
rect 332416 3612 332468 3664
rect 335268 3612 335320 3664
rect 389456 3612 389508 3664
rect 393964 3612 394016 3664
rect 413192 3612 413244 3664
rect 420184 3612 420236 3664
rect 553584 3612 553636 3664
rect 16028 3544 16080 3596
rect 142344 3544 142396 3596
rect 169392 3544 169444 3596
rect 214656 3544 214708 3596
rect 220084 3544 220136 3596
rect 224132 3544 224184 3596
rect 248512 3544 248564 3596
rect 291108 3544 291160 3596
rect 302608 3544 302660 3596
rect 303436 3544 303488 3596
rect 328828 3544 328880 3596
rect 331128 3544 331180 3596
rect 341616 3544 341668 3596
rect 343088 3544 343140 3596
rect 358176 3544 358228 3596
rect 360936 3544 360988 3596
rect 366916 3544 366968 3596
rect 369216 3544 369268 3596
rect 371608 3544 371660 3596
rect 398104 3544 398156 3596
rect 408316 3544 408368 3596
rect 408500 3544 408552 3596
rect 8852 3476 8904 3528
rect 9588 3476 9640 3528
rect 10048 3476 10100 3528
rect 138020 3476 138072 3528
rect 165896 3476 165948 3528
rect 219624 3476 219676 3528
rect 222200 3476 222252 3528
rect 222936 3476 222988 3528
rect 248604 3476 248656 3528
rect 257436 3476 257488 3528
rect 257988 3476 258040 3528
rect 259828 3476 259880 3528
rect 261484 3476 261536 3528
rect 262220 3476 262272 3528
rect 263508 3476 263560 3528
rect 290924 3476 290976 3528
rect 305000 3476 305052 3528
rect 305644 3476 305696 3528
rect 306288 3476 306340 3528
rect 309048 3476 309100 3528
rect 339500 3476 339552 3528
rect 344928 3476 344980 3528
rect 407304 3476 407356 3528
rect 417884 3476 417936 3528
rect 11244 3408 11296 3460
rect 139584 3408 139636 3460
rect 27896 3340 27948 3392
rect 28908 3340 28960 3392
rect 50528 3340 50580 3392
rect 159088 3340 159140 3392
rect 60004 3272 60056 3324
rect 60648 3272 60700 3324
rect 38568 3204 38620 3256
rect 81440 3272 81492 3324
rect 82544 3272 82596 3324
rect 82636 3272 82688 3324
rect 132592 3272 132644 3324
rect 133144 3272 133196 3324
rect 162308 3408 162360 3460
rect 219348 3408 219400 3460
rect 246028 3408 246080 3460
rect 270500 3408 270552 3460
rect 273352 3408 273404 3460
rect 285496 3408 285548 3460
rect 294328 3408 294380 3460
rect 295248 3408 295300 3460
rect 310980 3408 311032 3460
rect 313188 3408 313240 3460
rect 346676 3408 346728 3460
rect 351828 3408 351880 3460
rect 421564 3476 421616 3528
rect 424324 3544 424376 3596
rect 560760 3544 560812 3596
rect 439412 3476 439464 3528
rect 567844 3476 567896 3528
rect 418344 3408 418396 3460
rect 432328 3408 432380 3460
rect 442172 3408 442224 3460
rect 582196 3408 582248 3460
rect 189632 3340 189684 3392
rect 190368 3340 190420 3392
rect 197912 3340 197964 3392
rect 231860 3340 231912 3392
rect 250352 3340 250404 3392
rect 251088 3340 251140 3392
rect 293868 3340 293920 3392
rect 308588 3340 308640 3392
rect 320088 3340 320140 3392
rect 359740 3340 359792 3392
rect 389088 3340 389140 3392
rect 492956 3340 493008 3392
rect 493324 3340 493376 3392
rect 496084 3340 496136 3392
rect 510804 3340 510856 3392
rect 511264 3340 511316 3392
rect 564348 3340 564400 3392
rect 175648 3272 175700 3324
rect 93308 3204 93360 3256
rect 181076 3272 181128 3324
rect 198004 3272 198056 3324
rect 204260 3272 204312 3324
rect 217048 3272 217100 3324
rect 76012 3136 76064 3188
rect 99288 3136 99340 3188
rect 100024 3136 100076 3188
rect 100484 3136 100536 3188
rect 184940 3204 184992 3256
rect 192024 3204 192076 3256
rect 199200 3204 199252 3256
rect 181352 3136 181404 3188
rect 202696 3204 202748 3256
rect 229744 3204 229796 3256
rect 240784 3272 240836 3324
rect 241428 3272 241480 3324
rect 253848 3272 253900 3324
rect 257344 3272 257396 3324
rect 267004 3272 267056 3324
rect 267648 3272 267700 3324
rect 292488 3272 292540 3324
rect 306196 3272 306248 3324
rect 306288 3272 306340 3324
rect 314568 3272 314620 3324
rect 317328 3272 317380 3324
rect 353760 3272 353812 3324
rect 357808 3272 357860 3324
rect 378784 3272 378836 3324
rect 383476 3272 383528 3324
rect 482284 3272 482336 3324
rect 486424 3272 486476 3324
rect 500224 3272 500276 3324
rect 557172 3272 557224 3324
rect 243544 3204 243596 3256
rect 261024 3204 261076 3256
rect 262128 3204 262180 3256
rect 281448 3204 281500 3256
rect 285956 3204 286008 3256
rect 294604 3204 294656 3256
rect 301412 3204 301464 3256
rect 315856 3204 315908 3256
rect 321652 3204 321704 3256
rect 322204 3204 322256 3256
rect 357348 3204 357400 3256
rect 379428 3204 379480 3256
rect 475108 3204 475160 3256
rect 225604 3136 225656 3188
rect 281356 3136 281408 3188
rect 284760 3136 284812 3188
rect 297364 3136 297416 3188
rect 300308 3136 300360 3188
rect 302884 3136 302936 3188
rect 309784 3136 309836 3188
rect 320824 3136 320876 3188
rect 350264 3136 350316 3188
rect 375288 3136 375340 3188
rect 467932 3136 467984 3188
rect 474004 3136 474056 3188
rect 496544 3204 496596 3256
rect 546500 3204 546552 3256
rect 478144 3136 478196 3188
rect 503628 3136 503680 3188
rect 550088 3136 550140 3188
rect 107568 3068 107620 3120
rect 189264 3068 189316 3120
rect 206284 3068 206336 3120
rect 231124 3068 231176 3120
rect 232504 3068 232556 3120
rect 235356 3068 235408 3120
rect 258632 3068 258684 3120
rect 259368 3068 259420 3120
rect 264612 3068 264664 3120
rect 268384 3068 268436 3120
rect 372528 3068 372580 3120
rect 460848 3068 460900 3120
rect 469864 3068 469916 3120
rect 489368 3068 489420 3120
rect 114744 3000 114796 3052
rect 191840 3000 191892 3052
rect 193220 3000 193272 3052
rect 194508 3000 194560 3052
rect 202880 3000 202932 3052
rect 211068 3000 211120 3052
rect 217324 3000 217376 3052
rect 220544 3000 220596 3052
rect 232412 3000 232464 3052
rect 252652 3000 252704 3052
rect 254584 3000 254636 3052
rect 377404 3000 377456 3052
rect 453672 3000 453724 3052
rect 475384 3000 475436 3052
rect 489184 3000 489236 3052
rect 539324 3068 539376 3120
rect 532240 3000 532292 3052
rect 124220 2932 124272 2984
rect 125508 2932 125560 2984
rect 125416 2864 125468 2916
rect 197360 2932 197412 2984
rect 203892 2932 203944 2984
rect 220820 2932 220872 2984
rect 221740 2932 221792 2984
rect 228364 2932 228416 2984
rect 308404 2932 308456 2984
rect 313372 2932 313424 2984
rect 376024 2932 376076 2984
rect 414480 2932 414532 2984
rect 416044 2932 416096 2984
rect 418160 2932 418212 2984
rect 150440 2864 150492 2916
rect 192484 2864 192536 2916
rect 92112 2796 92164 2848
rect 92388 2796 92440 2848
rect 146852 2796 146904 2848
rect 185584 2796 185636 2848
rect 205088 2796 205140 2848
rect 208216 2796 208268 2848
rect 216956 2864 217008 2916
rect 223764 2864 223816 2916
rect 368940 2864 368992 2916
rect 428740 2864 428792 2916
rect 429844 2864 429896 2916
rect 482376 2932 482428 2984
rect 480904 2864 480956 2916
rect 485780 2864 485832 2916
rect 213184 2796 213236 2848
rect 340788 2796 340840 2848
rect 400220 2796 400272 2848
rect 402244 2796 402296 2848
rect 446588 2796 446640 2848
rect 525064 2864 525116 2916
rect 517888 2796 517940 2848
rect 194416 1300 194468 1352
rect 23112 552 23164 604
rect 23388 552 23440 604
rect 67180 595 67232 604
rect 67180 561 67189 595
rect 67189 561 67223 595
rect 67223 561 67232 595
rect 67180 552 67232 561
rect 178960 552 179012 604
rect 179328 552 179380 604
rect 230112 552 230164 604
rect 230388 552 230440 604
rect 238392 552 238444 604
rect 238668 552 238720 604
rect 272892 552 272944 604
rect 273168 552 273220 604
rect 290096 552 290148 604
rect 290740 552 290792 604
rect 291384 552 291436 604
rect 291936 552 291988 604
rect 318984 552 319036 604
rect 319260 552 319312 604
rect 326436 595 326488 604
rect 326436 561 326445 595
rect 326445 561 326479 595
rect 326479 561 326488 595
rect 326436 552 326488 561
rect 332876 552 332928 604
rect 333612 552 333664 604
rect 336924 552 336976 604
rect 337108 552 337160 604
rect 343916 552 343968 604
rect 344284 552 344336 604
rect 456800 552 456852 604
rect 457260 552 457312 604
rect 470600 552 470652 604
rect 471520 552 471572 604
rect 473360 552 473412 604
rect 473912 552 473964 604
<< metal2 >>
rect 8086 703520 8198 704960
rect 24278 703520 24390 704960
rect 40470 703520 40582 704960
rect 56754 703520 56866 704960
rect 72946 703520 73058 704960
rect 89138 703520 89250 704960
rect 105422 703520 105534 704960
rect 121614 703520 121726 704960
rect 137806 703520 137918 704960
rect 154090 703520 154202 704960
rect 170282 703520 170394 704960
rect 186474 703520 186586 704960
rect 202758 703520 202870 704960
rect 218950 703520 219062 704960
rect 235142 703520 235254 704960
rect 251426 703520 251538 704960
rect 267618 703520 267730 704960
rect 283810 703520 283922 704960
rect 300094 703520 300206 704960
rect 316286 703520 316398 704960
rect 332478 703520 332590 704960
rect 348762 703520 348874 704960
rect 364954 703520 365066 704960
rect 381146 703520 381258 704960
rect 397430 703520 397542 704960
rect 413622 703520 413734 704960
rect 429814 703520 429926 704960
rect 446098 703520 446210 704960
rect 462290 703520 462402 704960
rect 478482 703520 478594 704960
rect 494766 703520 494878 704960
rect 510958 703520 511070 704960
rect 527150 703520 527262 704960
rect 543434 703520 543546 704960
rect 559626 703520 559738 704960
rect 575818 703520 575930 704960
rect 8128 700398 8156 703520
rect 8116 700392 8168 700398
rect 8116 700334 8168 700340
rect 13084 700392 13136 700398
rect 13084 700334 13136 700340
rect 3514 682272 3570 682281
rect 3514 682207 3570 682216
rect 3528 681766 3556 682207
rect 3516 681760 3568 681766
rect 3516 681702 3568 681708
rect 3422 667992 3478 668001
rect 3422 667927 3424 667936
rect 3476 667927 3478 667936
rect 3424 667898 3476 667904
rect 4802 653576 4858 653585
rect 4802 653511 4858 653520
rect 3422 624880 3478 624889
rect 3422 624815 3478 624824
rect 3436 623830 3464 624815
rect 3424 623824 3476 623830
rect 3424 623766 3476 623772
rect 3422 610464 3478 610473
rect 3422 610399 3478 610408
rect 3436 610026 3464 610399
rect 3424 610020 3476 610026
rect 3424 609962 3476 609968
rect 4066 596048 4122 596057
rect 4066 595983 4122 595992
rect 4080 594862 4108 595983
rect 4068 594856 4120 594862
rect 4068 594798 4120 594804
rect 3422 567352 3478 567361
rect 3422 567287 3478 567296
rect 3146 553072 3202 553081
rect 3146 553007 3202 553016
rect 3160 552090 3188 553007
rect 3148 552084 3200 552090
rect 3148 552026 3200 552032
rect 3330 495544 3386 495553
rect 3330 495479 3332 495488
rect 3384 495479 3386 495488
rect 3332 495450 3384 495456
rect 3054 452432 3110 452441
rect 3054 452367 3110 452376
rect 3068 451382 3096 452367
rect 3056 451376 3108 451382
rect 3056 451318 3108 451324
rect 2778 366208 2834 366217
rect 2778 366143 2834 366152
rect 2792 365770 2820 366143
rect 2780 365764 2832 365770
rect 2780 365706 2832 365712
rect 2962 337512 3018 337521
rect 2962 337447 3018 337456
rect 2976 336802 3004 337447
rect 2964 336796 3016 336802
rect 2964 336738 3016 336744
rect 3330 294400 3386 294409
rect 3330 294335 3386 294344
rect 3344 294030 3372 294335
rect 3332 294024 3384 294030
rect 3332 293966 3384 293972
rect 2778 265704 2834 265713
rect 2778 265639 2834 265648
rect 2792 264994 2820 265639
rect 2780 264988 2832 264994
rect 2780 264930 2832 264936
rect 3330 251288 3386 251297
rect 3330 251223 3332 251232
rect 3384 251223 3386 251232
rect 3332 251194 3384 251200
rect 3330 237008 3386 237017
rect 3330 236943 3386 236952
rect 2962 222592 3018 222601
rect 2962 222527 3018 222536
rect 2976 222222 3004 222527
rect 2964 222216 3016 222222
rect 2964 222158 3016 222164
rect 2962 208176 3018 208185
rect 2962 208111 3018 208120
rect 2976 207058 3004 208111
rect 2964 207052 3016 207058
rect 2964 206994 3016 207000
rect 3240 200184 3292 200190
rect 3240 200126 3292 200132
rect 2872 180804 2924 180810
rect 2872 180746 2924 180752
rect 2884 179489 2912 180746
rect 2870 179480 2926 179489
rect 2870 179415 2926 179424
rect 3252 165073 3280 200126
rect 3238 165064 3294 165073
rect 3238 164999 3294 165008
rect 3240 156052 3292 156058
rect 3240 155994 3292 156000
rect 3252 150793 3280 155994
rect 3344 154358 3372 236943
rect 3436 201006 3464 567287
rect 3514 538656 3570 538665
rect 3514 538591 3570 538600
rect 3424 201000 3476 201006
rect 3424 200942 3476 200948
rect 3424 197396 3476 197402
rect 3424 197338 3476 197344
rect 3332 154352 3384 154358
rect 3332 154294 3384 154300
rect 3238 150784 3294 150793
rect 3238 150719 3294 150728
rect 3332 136604 3384 136610
rect 3332 136546 3384 136552
rect 3344 136377 3372 136546
rect 3330 136368 3386 136377
rect 3330 136303 3386 136312
rect 3054 122088 3110 122097
rect 3054 122023 3110 122032
rect 3068 121038 3096 122023
rect 3056 121032 3108 121038
rect 3056 120974 3108 120980
rect 2780 93356 2832 93362
rect 2780 93298 2832 93304
rect 2792 93265 2820 93298
rect 2778 93256 2834 93265
rect 2778 93191 2834 93200
rect 3240 80028 3292 80034
rect 3240 79970 3292 79976
rect 3252 78985 3280 79970
rect 3238 78976 3294 78985
rect 3238 78911 3294 78920
rect 3332 64864 3384 64870
rect 3332 64806 3384 64812
rect 3344 64569 3372 64806
rect 3330 64560 3386 64569
rect 3330 64495 3386 64504
rect 3436 50153 3464 197338
rect 3528 189038 3556 538591
rect 3606 509960 3662 509969
rect 3606 509895 3662 509904
rect 3620 201074 3648 509895
rect 4066 481128 4122 481137
rect 4066 481063 4122 481072
rect 4080 480690 4108 481063
rect 4068 480684 4120 480690
rect 4068 480626 4120 480632
rect 3698 438016 3754 438025
rect 3698 437951 3754 437960
rect 3608 201068 3660 201074
rect 3608 201010 3660 201016
rect 3606 193896 3662 193905
rect 3606 193831 3662 193840
rect 3516 189032 3568 189038
rect 3516 188974 3568 188980
rect 3516 156120 3568 156126
rect 3516 156062 3568 156068
rect 3528 107681 3556 156062
rect 3620 155922 3648 193831
rect 3608 155916 3660 155922
rect 3608 155858 3660 155864
rect 3712 150414 3740 437951
rect 4066 423736 4122 423745
rect 4066 423671 4068 423680
rect 4120 423671 4122 423680
rect 4068 423642 4120 423648
rect 3882 395040 3938 395049
rect 3882 394975 3938 394984
rect 3790 380624 3846 380633
rect 3790 380559 3846 380568
rect 3804 151774 3832 380559
rect 3896 201142 3924 394975
rect 3974 323096 4030 323105
rect 3974 323031 4030 323040
rect 3884 201136 3936 201142
rect 3884 201078 3936 201084
rect 3988 152930 4016 323031
rect 4066 308816 4122 308825
rect 4066 308751 4122 308760
rect 4080 307834 4108 308751
rect 4068 307828 4120 307834
rect 4068 307770 4120 307776
rect 4066 280120 4122 280129
rect 4066 280055 4122 280064
rect 4080 153202 4108 280055
rect 4816 186318 4844 653511
rect 4896 594856 4948 594862
rect 4896 594798 4948 594804
rect 4908 187678 4936 594798
rect 4988 480684 5040 480690
rect 4988 480626 5040 480632
rect 5000 188970 5028 480626
rect 5080 423700 5132 423706
rect 5080 423642 5132 423648
rect 5092 190466 5120 423642
rect 5172 365764 5224 365770
rect 5172 365706 5224 365712
rect 5184 191826 5212 365706
rect 5264 307828 5316 307834
rect 5264 307770 5316 307776
rect 5276 193186 5304 307770
rect 5448 264988 5500 264994
rect 5448 264930 5500 264936
rect 5356 196308 5408 196314
rect 5356 196250 5408 196256
rect 5264 193180 5316 193186
rect 5264 193122 5316 193128
rect 5172 191820 5224 191826
rect 5172 191762 5224 191768
rect 5080 190460 5132 190466
rect 5080 190402 5132 190408
rect 4988 188964 5040 188970
rect 4988 188906 5040 188912
rect 4896 187672 4948 187678
rect 4896 187614 4948 187620
rect 4804 186312 4856 186318
rect 4804 186254 4856 186260
rect 4068 153196 4120 153202
rect 4068 153138 4120 153144
rect 3976 152924 4028 152930
rect 3976 152866 4028 152872
rect 3792 151768 3844 151774
rect 3792 151710 3844 151716
rect 3700 150408 3752 150414
rect 3700 150350 3752 150356
rect 3514 107672 3570 107681
rect 3514 107607 3570 107616
rect 5368 93362 5396 196250
rect 5460 193118 5488 264930
rect 5448 193112 5500 193118
rect 5448 193054 5500 193060
rect 13096 184890 13124 700334
rect 24320 699718 24348 703520
rect 40512 700330 40540 703520
rect 40500 700324 40552 700330
rect 40500 700266 40552 700272
rect 72988 699718 73016 703520
rect 89180 700398 89208 703520
rect 105464 700466 105492 703520
rect 133880 701004 133932 701010
rect 133880 700946 133932 700952
rect 133788 700936 133840 700942
rect 133788 700878 133840 700884
rect 132500 700868 132552 700874
rect 132500 700810 132552 700816
rect 131120 700732 131172 700738
rect 131120 700674 131172 700680
rect 105452 700460 105504 700466
rect 105452 700402 105504 700408
rect 89168 700392 89220 700398
rect 89168 700334 89220 700340
rect 126244 700392 126296 700398
rect 126244 700334 126296 700340
rect 24308 699712 24360 699718
rect 24308 699654 24360 699660
rect 24768 699712 24820 699718
rect 24768 699654 24820 699660
rect 72424 699712 72476 699718
rect 72424 699654 72476 699660
rect 72976 699712 73028 699718
rect 72976 699654 73028 699660
rect 19984 667956 20036 667962
rect 19984 667898 20036 667904
rect 14464 222216 14516 222222
rect 14464 222158 14516 222164
rect 14476 194546 14504 222158
rect 17224 196104 17276 196110
rect 17224 196046 17276 196052
rect 15844 194676 15896 194682
rect 15844 194618 15896 194624
rect 14464 194540 14516 194546
rect 14464 194482 14516 194488
rect 13084 184884 13136 184890
rect 13084 184826 13136 184832
rect 15856 180810 15884 194618
rect 15844 180804 15896 180810
rect 15844 180746 15896 180752
rect 17236 136610 17264 196046
rect 19996 146266 20024 667898
rect 21364 610020 21416 610026
rect 21364 609962 21416 609968
rect 21376 147626 21404 609962
rect 21364 147620 21416 147626
rect 21364 147562 21416 147568
rect 19984 146260 20036 146266
rect 19984 146202 20036 146208
rect 24780 144702 24808 699654
rect 28264 552084 28316 552090
rect 28264 552026 28316 552032
rect 28276 149054 28304 552026
rect 70124 524476 70176 524482
rect 70124 524418 70176 524424
rect 69848 500268 69900 500274
rect 69848 500210 69900 500216
rect 31024 495508 31076 495514
rect 31024 495450 31076 495456
rect 28264 149048 28316 149054
rect 28264 148990 28316 148996
rect 31036 148986 31064 495450
rect 69860 377913 69888 500210
rect 69940 396840 69992 396846
rect 69940 396782 69992 396788
rect 69952 385257 69980 396782
rect 70032 395684 70084 395690
rect 70032 395626 70084 395632
rect 69938 385248 69994 385257
rect 69938 385183 69994 385192
rect 69846 377904 69902 377913
rect 69846 377839 69902 377848
rect 70044 362953 70072 395626
rect 70030 362944 70086 362953
rect 70030 362879 70086 362888
rect 70030 355600 70086 355609
rect 70030 355535 70086 355544
rect 70044 341465 70072 355535
rect 70136 348265 70164 524418
rect 70216 407788 70268 407794
rect 70216 407730 70268 407736
rect 70228 370297 70256 407730
rect 70308 406564 70360 406570
rect 70308 406506 70360 406512
rect 70320 392601 70348 406506
rect 71688 398880 71740 398886
rect 71688 398822 71740 398828
rect 70306 392592 70362 392601
rect 70306 392527 70362 392536
rect 71594 392592 71650 392601
rect 71594 392527 71650 392536
rect 70306 377904 70362 377913
rect 70306 377839 70362 377848
rect 70214 370288 70270 370297
rect 70214 370223 70270 370232
rect 70122 348256 70178 348265
rect 70122 348191 70178 348200
rect 70030 341456 70086 341465
rect 70030 341391 70086 341400
rect 31024 148980 31076 148986
rect 31024 148922 31076 148928
rect 24768 144696 24820 144702
rect 24768 144638 24820 144644
rect 17224 136604 17276 136610
rect 17224 136546 17276 136552
rect 67548 119128 67600 119134
rect 67548 119070 67600 119076
rect 31668 118244 31720 118250
rect 31668 118186 31720 118192
rect 28908 118176 28960 118182
rect 28908 118118 28960 118124
rect 23388 118108 23440 118114
rect 23388 118050 23440 118056
rect 9588 117972 9640 117978
rect 9588 117914 9640 117920
rect 5356 93356 5408 93362
rect 5356 93298 5408 93304
rect 3422 50144 3478 50153
rect 3422 50079 3478 50088
rect 3424 35896 3476 35902
rect 3422 35864 3424 35873
rect 3476 35864 3478 35873
rect 3422 35799 3478 35808
rect 3148 22092 3200 22098
rect 3148 22034 3200 22040
rect 3160 21457 3188 22034
rect 3146 21448 3202 21457
rect 3146 21383 3202 21392
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 3424 8288 3476 8294
rect 3424 8230 3476 8236
rect 1676 7812 1728 7818
rect 1676 7754 1728 7760
rect 572 7608 624 7614
rect 572 7550 624 7556
rect 584 480 612 7550
rect 1688 480 1716 7754
rect 2872 7676 2924 7682
rect 2872 7618 2924 7624
rect 2884 480 2912 7618
rect 3436 7177 3464 8230
rect 5264 7744 5316 7750
rect 5264 7686 5316 7692
rect 3422 7168 3478 7177
rect 3422 7103 3478 7112
rect 4068 4820 4120 4826
rect 4068 4762 4120 4768
rect 4080 480 4108 4762
rect 5276 480 5304 7686
rect 6472 480 6500 8910
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7668 480 7696 7822
rect 9600 3534 9628 117914
rect 20720 8016 20772 8022
rect 20720 7958 20772 7964
rect 13636 7948 13688 7954
rect 13636 7890 13688 7896
rect 12440 4888 12492 4894
rect 12440 4830 12492 4836
rect 8852 3528 8904 3534
rect 8852 3470 8904 3476
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 10048 3528 10100 3534
rect 10048 3470 10100 3476
rect 8864 480 8892 3470
rect 10060 480 10088 3470
rect 11244 3460 11296 3466
rect 11244 3402 11296 3408
rect 11256 480 11284 3402
rect 12452 480 12480 4830
rect 13648 480 13676 7890
rect 18328 5092 18380 5098
rect 18328 5034 18380 5040
rect 17224 4956 17276 4962
rect 17224 4898 17276 4904
rect 14832 3664 14884 3670
rect 14832 3606 14884 3612
rect 14844 480 14872 3606
rect 16028 3596 16080 3602
rect 16028 3538 16080 3544
rect 16040 480 16068 3538
rect 17236 480 17264 4898
rect 18340 480 18368 5034
rect 19524 3732 19576 3738
rect 19524 3674 19576 3680
rect 19536 480 19564 3674
rect 20732 480 20760 7958
rect 21916 5024 21968 5030
rect 21916 4966 21968 4972
rect 21928 480 21956 4966
rect 23400 610 23428 118050
rect 26700 9036 26752 9042
rect 26700 8978 26752 8984
rect 25504 3868 25556 3874
rect 25504 3810 25556 3816
rect 24308 3800 24360 3806
rect 24308 3742 24360 3748
rect 23112 604 23164 610
rect 23112 546 23164 552
rect 23388 604 23440 610
rect 23388 546 23440 552
rect 23124 480 23152 546
rect 24320 480 24348 3742
rect 25516 480 25544 3810
rect 26712 480 26740 8978
rect 28920 3398 28948 118118
rect 29092 6180 29144 6186
rect 29092 6122 29144 6128
rect 27896 3392 27948 3398
rect 27896 3334 27948 3340
rect 28908 3392 28960 3398
rect 28908 3334 28960 3340
rect 27908 480 27936 3334
rect 29104 480 29132 6122
rect 30286 4856 30342 4865
rect 30286 4791 30342 4800
rect 30300 480 30328 4791
rect 31680 626 31708 118186
rect 60648 118040 60700 118046
rect 60648 117982 60700 117988
rect 55220 9376 55272 9382
rect 55220 9318 55272 9324
rect 54024 9240 54076 9246
rect 54024 9182 54076 9188
rect 46940 9172 46992 9178
rect 46940 9114 46992 9120
rect 40960 9104 41012 9110
rect 40960 9046 41012 9052
rect 34980 8220 35032 8226
rect 34980 8162 35032 8168
rect 33876 5160 33928 5166
rect 33876 5102 33928 5108
rect 32680 3936 32732 3942
rect 32680 3878 32732 3884
rect 31496 598 31708 626
rect 31496 480 31524 598
rect 32692 480 32720 3878
rect 33888 480 33916 5102
rect 34992 480 35020 8162
rect 36176 6248 36228 6254
rect 36176 6190 36228 6196
rect 36188 480 36216 6190
rect 37372 5228 37424 5234
rect 37372 5170 37424 5176
rect 37384 480 37412 5170
rect 39764 4004 39816 4010
rect 39764 3946 39816 3952
rect 38568 3256 38620 3262
rect 38568 3198 38620 3204
rect 38580 480 38608 3198
rect 39776 480 39804 3946
rect 40972 480 41000 9046
rect 44548 5296 44600 5302
rect 44548 5238 44600 5244
rect 42156 4140 42208 4146
rect 42156 4082 42208 4088
rect 42168 480 42196 4082
rect 43352 4072 43404 4078
rect 43352 4014 43404 4020
rect 43364 480 43392 4014
rect 44560 480 44588 5238
rect 45744 4412 45796 4418
rect 45744 4354 45796 4360
rect 45756 480 45784 4354
rect 46952 480 46980 9114
rect 51632 8152 51684 8158
rect 51632 8094 51684 8100
rect 48136 8084 48188 8090
rect 48136 8026 48188 8032
rect 48148 480 48176 8026
rect 49332 4480 49384 4486
rect 49332 4422 49384 4428
rect 49344 480 49372 4422
rect 50528 3392 50580 3398
rect 50528 3334 50580 3340
rect 50540 480 50568 3334
rect 51644 480 51672 8094
rect 52828 4344 52880 4350
rect 52828 4286 52880 4292
rect 52840 480 52868 4286
rect 54036 480 54064 9182
rect 55232 480 55260 9318
rect 58808 9308 58860 9314
rect 58808 9250 58860 9256
rect 57612 6316 57664 6322
rect 57612 6258 57664 6264
rect 56416 5840 56468 5846
rect 56416 5782 56468 5788
rect 56428 480 56456 5782
rect 57624 480 57652 6258
rect 58820 480 58848 9250
rect 60660 3330 60688 117982
rect 61200 9444 61252 9450
rect 61200 9386 61252 9392
rect 60004 3324 60056 3330
rect 60004 3266 60056 3272
rect 60648 3324 60700 3330
rect 60648 3266 60700 3272
rect 60016 480 60044 3266
rect 61212 480 61240 9386
rect 64788 6384 64840 6390
rect 64788 6326 64840 6332
rect 62396 5364 62448 5370
rect 62396 5306 62448 5312
rect 62408 480 62436 5306
rect 63592 4276 63644 4282
rect 63592 4218 63644 4224
rect 63604 480 63632 4218
rect 64800 480 64828 6326
rect 65984 5432 66036 5438
rect 65984 5374 66036 5380
rect 65996 480 66024 5374
rect 67560 4214 67588 119070
rect 70228 117978 70256 370223
rect 70320 119134 70348 377839
rect 71502 348256 71558 348265
rect 71502 348191 71558 348200
rect 70308 119128 70360 119134
rect 70308 119070 70360 119076
rect 71516 118386 71544 348191
rect 71504 118380 71556 118386
rect 71504 118322 71556 118328
rect 71608 118017 71636 392527
rect 71700 118318 71728 398822
rect 72436 183530 72464 699654
rect 119344 583364 119396 583370
rect 119344 583306 119396 583312
rect 85396 583296 85448 583302
rect 85396 583238 85448 583244
rect 84106 545864 84162 545873
rect 84106 545799 84162 545808
rect 84014 541512 84070 541521
rect 84014 541447 84070 541456
rect 83922 528728 83978 528737
rect 83922 528663 83978 528672
rect 82818 524920 82874 524929
rect 82818 524855 82874 524864
rect 82832 524482 82860 524855
rect 82820 524476 82872 524482
rect 82820 524418 82872 524424
rect 83936 497554 83964 528663
rect 83924 497548 83976 497554
rect 83924 497490 83976 497496
rect 75828 398132 75880 398138
rect 75828 398074 75880 398080
rect 75840 396250 75868 398074
rect 80796 397928 80848 397934
rect 80796 397870 80848 397876
rect 80808 396250 80836 397870
rect 75532 396222 75868 396250
rect 80500 396222 80836 396250
rect 84028 395894 84056 541447
rect 84016 395888 84068 395894
rect 84016 395830 84068 395836
rect 84120 395758 84148 545799
rect 85302 537160 85358 537169
rect 85302 537095 85358 537104
rect 85210 533080 85266 533089
rect 85210 533015 85266 533024
rect 85224 521286 85252 533015
rect 85212 521280 85264 521286
rect 85212 521222 85264 521228
rect 85316 520946 85344 537095
rect 85408 525609 85436 583238
rect 115388 578400 115440 578406
rect 115388 578342 115440 578348
rect 115204 578332 115256 578338
rect 115204 578274 115256 578280
rect 110328 575544 110380 575550
rect 110328 575486 110380 575492
rect 110340 554810 110368 575486
rect 109408 554804 109460 554810
rect 109408 554746 109460 554752
rect 110328 554804 110380 554810
rect 110328 554746 110380 554752
rect 92112 553988 92164 553994
rect 92112 553930 92164 553936
rect 89168 553920 89220 553926
rect 89168 553862 89220 553868
rect 89180 551820 89208 553862
rect 92124 551820 92152 553930
rect 95056 553784 95108 553790
rect 95056 553726 95108 553732
rect 95068 551820 95096 553726
rect 100760 553716 100812 553722
rect 100760 553658 100812 553664
rect 97816 553512 97868 553518
rect 97816 553454 97868 553460
rect 97828 551820 97856 553454
rect 100772 551820 100800 553658
rect 106464 553648 106516 553654
rect 106464 553590 106516 553596
rect 103704 553580 103756 553586
rect 103704 553522 103756 553528
rect 103716 551820 103744 553522
rect 106476 551820 106504 553590
rect 109420 551820 109448 554746
rect 115112 553852 115164 553858
rect 115112 553794 115164 553800
rect 112352 553444 112404 553450
rect 112352 553386 112404 553392
rect 112364 551820 112392 553386
rect 115124 551820 115152 553794
rect 86406 549944 86462 549953
rect 85488 549908 85540 549914
rect 86406 549879 86408 549888
rect 85488 549850 85540 549856
rect 86460 549879 86462 549888
rect 86408 549850 86460 549856
rect 85394 525600 85450 525609
rect 85394 525535 85450 525544
rect 85304 520940 85356 520946
rect 85304 520882 85356 520888
rect 85500 398886 85528 549850
rect 86604 518770 86632 520132
rect 89364 518906 89392 520132
rect 89352 518900 89404 518906
rect 89352 518842 89404 518848
rect 86592 518764 86644 518770
rect 86592 518706 86644 518712
rect 92308 518226 92336 520132
rect 92296 518220 92348 518226
rect 92296 518162 92348 518168
rect 95252 500274 95280 520132
rect 98012 518430 98040 520132
rect 98000 518424 98052 518430
rect 98000 518366 98052 518372
rect 100956 518294 100984 520132
rect 103532 520118 103914 520146
rect 100944 518288 100996 518294
rect 100944 518230 100996 518236
rect 96528 500948 96580 500954
rect 96528 500890 96580 500896
rect 96540 500274 96568 500890
rect 103532 500886 103560 520118
rect 106660 518362 106688 520132
rect 109604 518838 109632 520132
rect 111812 520118 112562 520146
rect 109592 518832 109644 518838
rect 109592 518774 109644 518780
rect 106648 518356 106700 518362
rect 106648 518298 106700 518304
rect 103520 500880 103572 500886
rect 103520 500822 103572 500828
rect 104808 500880 104860 500886
rect 104808 500822 104860 500828
rect 95240 500268 95292 500274
rect 95240 500210 95292 500216
rect 96528 500268 96580 500274
rect 96528 500210 96580 500216
rect 104820 407794 104848 500822
rect 111708 497684 111760 497690
rect 111708 497626 111760 497632
rect 108948 497616 109000 497622
rect 108948 497558 109000 497564
rect 104808 407788 104860 407794
rect 104808 407730 104860 407736
rect 85488 398880 85540 398886
rect 85488 398822 85540 398828
rect 85500 398750 85528 398822
rect 85488 398744 85540 398750
rect 85488 398686 85540 398692
rect 90272 398744 90324 398750
rect 90272 398686 90324 398692
rect 85948 397588 86000 397594
rect 85948 397530 86000 397536
rect 85960 396250 85988 397530
rect 85652 396222 85988 396250
rect 90284 396250 90312 398686
rect 100668 397860 100720 397866
rect 100668 397802 100720 397808
rect 95884 397656 95936 397662
rect 95884 397598 95936 397604
rect 95896 396250 95924 397598
rect 100680 396250 100708 397802
rect 106004 397724 106056 397730
rect 106004 397666 106056 397672
rect 106016 396250 106044 397666
rect 90284 396222 90620 396250
rect 95588 396222 95924 396250
rect 100556 396222 100708 396250
rect 105708 396222 106044 396250
rect 84108 395752 84160 395758
rect 84108 395694 84160 395700
rect 108960 395690 108988 497558
rect 111720 397798 111748 497626
rect 111812 497486 111840 520118
rect 115216 518838 115244 578274
rect 115296 553988 115348 553994
rect 115296 553930 115348 553936
rect 113180 518832 113232 518838
rect 113180 518774 113232 518780
rect 115204 518832 115256 518838
rect 115204 518774 115256 518780
rect 111800 497480 111852 497486
rect 111800 497422 111852 497428
rect 113192 397866 113220 518774
rect 115308 498137 115336 553930
rect 115400 549914 115428 578342
rect 115940 554804 115992 554810
rect 115940 554746 115992 554752
rect 115388 549908 115440 549914
rect 115388 549850 115440 549856
rect 115294 498128 115350 498137
rect 115294 498063 115350 498072
rect 115308 497690 115336 498063
rect 115296 497684 115348 497690
rect 115296 497626 115348 497632
rect 115952 398138 115980 554746
rect 116032 553444 116084 553450
rect 116032 553386 116084 553392
rect 116044 498098 116072 553386
rect 118054 546544 118110 546553
rect 118054 546479 118110 546488
rect 117778 537432 117834 537441
rect 117778 537367 117834 537376
rect 117792 536858 117820 537367
rect 117780 536852 117832 536858
rect 117780 536794 117832 536800
rect 117778 533352 117834 533361
rect 117778 533287 117834 533296
rect 117792 532778 117820 533287
rect 117780 532772 117832 532778
rect 117780 532714 117832 532720
rect 117964 529916 118016 529922
rect 117964 529858 118016 529864
rect 117976 529689 118004 529858
rect 117962 529680 118018 529689
rect 117962 529615 118018 529624
rect 117318 521112 117374 521121
rect 117318 521047 117374 521056
rect 117332 521014 117360 521047
rect 117320 521008 117372 521014
rect 117320 520950 117372 520956
rect 116032 498092 116084 498098
rect 116032 498034 116084 498040
rect 116044 497622 116072 498034
rect 116032 497616 116084 497622
rect 116032 497558 116084 497564
rect 115940 398132 115992 398138
rect 115940 398074 115992 398080
rect 113180 397860 113232 397866
rect 113180 397802 113232 397808
rect 114468 397860 114520 397866
rect 114468 397802 114520 397808
rect 110972 397792 111024 397798
rect 110972 397734 111024 397740
rect 111708 397792 111760 397798
rect 111708 397734 111760 397740
rect 110984 396250 111012 397734
rect 114480 396778 114508 397802
rect 115848 397520 115900 397526
rect 115848 397462 115900 397468
rect 114468 396772 114520 396778
rect 114468 396714 114520 396720
rect 115860 396250 115888 397462
rect 117976 396846 118004 529615
rect 118068 499526 118096 546479
rect 118606 542464 118662 542473
rect 118606 542399 118608 542408
rect 118660 542399 118662 542408
rect 118608 542370 118660 542376
rect 119356 529922 119384 583306
rect 124862 582584 124918 582593
rect 124862 582519 124918 582528
rect 122748 578468 122800 578474
rect 122748 578410 122800 578416
rect 120724 553784 120776 553790
rect 120724 553726 120776 553732
rect 119344 529916 119396 529922
rect 119344 529858 119396 529864
rect 118606 525192 118662 525201
rect 118606 525127 118662 525136
rect 118620 525094 118648 525127
rect 118608 525088 118660 525094
rect 118608 525030 118660 525036
rect 118056 499520 118108 499526
rect 118056 499462 118108 499468
rect 120736 498030 120764 553726
rect 122760 518770 122788 578410
rect 122748 518764 122800 518770
rect 122748 518706 122800 518712
rect 120724 498024 120776 498030
rect 120724 497966 120776 497972
rect 121368 498024 121420 498030
rect 121368 497966 121420 497972
rect 121380 399362 121408 497966
rect 120908 399356 120960 399362
rect 120908 399298 120960 399304
rect 121368 399356 121420 399362
rect 121368 399298 121420 399304
rect 117964 396840 118016 396846
rect 117964 396782 118016 396788
rect 120920 396250 120948 399298
rect 124876 397934 124904 582519
rect 125968 497480 126020 497486
rect 125968 497422 126020 497428
rect 125980 495553 126008 497422
rect 125966 495544 126022 495553
rect 125966 495479 126022 495488
rect 125874 492688 125930 492697
rect 125874 492623 125930 492632
rect 125888 486418 125916 492623
rect 125888 486390 126008 486418
rect 125980 481642 126008 486390
rect 125968 481636 126020 481642
rect 125968 481578 126020 481584
rect 126060 481636 126112 481642
rect 126060 481578 126112 481584
rect 126072 466290 126100 481578
rect 125980 466262 126100 466290
rect 125980 456890 126008 466262
rect 125968 456884 126020 456890
rect 125968 456826 126020 456832
rect 125968 456748 126020 456754
rect 125968 456690 126020 456696
rect 125980 454034 126008 456690
rect 125968 454028 126020 454034
rect 125968 453970 126020 453976
rect 126060 454028 126112 454034
rect 126060 453970 126112 453976
rect 126072 452606 126100 453970
rect 126060 452600 126112 452606
rect 126060 452542 126112 452548
rect 126060 443828 126112 443834
rect 126060 443770 126112 443776
rect 126072 437458 126100 443770
rect 125980 437430 126100 437458
rect 125980 434722 126008 437430
rect 125968 434716 126020 434722
rect 125968 434658 126020 434664
rect 125876 427780 125928 427786
rect 125876 427722 125928 427728
rect 125888 425082 125916 427722
rect 125888 425066 126008 425082
rect 125876 425060 126020 425066
rect 125928 425054 125968 425060
rect 125876 425002 125928 425008
rect 125968 425002 126020 425008
rect 125888 415449 125916 425002
rect 125980 424971 126008 425002
rect 125874 415440 125930 415449
rect 125874 415375 125930 415384
rect 126150 415440 126206 415449
rect 126150 415375 126152 415384
rect 126204 415375 126206 415384
rect 126152 415346 126204 415352
rect 126060 405748 126112 405754
rect 126060 405690 126112 405696
rect 125692 399356 125744 399362
rect 125692 399298 125744 399304
rect 124864 397928 124916 397934
rect 124864 397870 124916 397876
rect 124876 397458 124904 397870
rect 124864 397452 124916 397458
rect 124864 397394 124916 397400
rect 110676 396222 111012 396250
rect 115644 396222 115888 396250
rect 120612 396222 120948 396250
rect 125704 395808 125732 399298
rect 126072 398834 126100 405690
rect 125888 398806 126100 398834
rect 125888 395842 125916 398806
rect 126152 397452 126204 397458
rect 126152 397394 126204 397400
rect 125888 395814 126008 395842
rect 125704 395780 125824 395808
rect 125690 395720 125746 395729
rect 108948 395684 109000 395690
rect 125580 395678 125690 395706
rect 125690 395655 125746 395664
rect 108948 395626 109000 395632
rect 125796 394482 125824 395780
rect 125876 395684 125928 395690
rect 125876 395626 125928 395632
rect 125704 394454 125824 394482
rect 111708 340264 111760 340270
rect 111708 340206 111760 340212
rect 110328 340196 110380 340202
rect 110328 340138 110380 340144
rect 72588 340054 72924 340082
rect 77556 340054 77892 340082
rect 82524 340054 82768 340082
rect 87492 340054 87828 340082
rect 92460 340054 92796 340082
rect 97612 340054 97948 340082
rect 102580 340054 102916 340082
rect 107548 340054 107608 340082
rect 72896 337482 72924 340054
rect 72884 337476 72936 337482
rect 72884 337418 72936 337424
rect 77864 337414 77892 340054
rect 77852 337408 77904 337414
rect 77852 337350 77904 337356
rect 82740 336734 82768 340054
rect 87800 337958 87828 340054
rect 87788 337952 87840 337958
rect 87788 337894 87840 337900
rect 92768 336870 92796 340054
rect 97920 338026 97948 340054
rect 97908 338020 97960 338026
rect 97908 337962 97960 337968
rect 92756 336864 92808 336870
rect 92756 336806 92808 336812
rect 93768 336864 93820 336870
rect 93768 336806 93820 336812
rect 82728 336728 82780 336734
rect 82728 336670 82780 336676
rect 72424 183524 72476 183530
rect 72424 183466 72476 183472
rect 75920 118584 75972 118590
rect 75918 118552 75920 118561
rect 75972 118552 75974 118561
rect 82740 118522 82768 336670
rect 93780 202162 93808 336806
rect 93768 202156 93820 202162
rect 93768 202098 93820 202104
rect 97920 118590 97948 337962
rect 100668 337408 100720 337414
rect 100668 337350 100720 337356
rect 97908 118584 97960 118590
rect 85394 118552 85450 118561
rect 75918 118487 75974 118496
rect 82728 118516 82780 118522
rect 97908 118526 97960 118532
rect 85394 118487 85450 118496
rect 82728 118458 82780 118464
rect 85408 118402 85436 118487
rect 85488 118448 85540 118454
rect 85408 118396 85488 118402
rect 85408 118390 85540 118396
rect 85408 118374 85528 118390
rect 88340 118380 88392 118386
rect 88340 118322 88392 118328
rect 71688 118312 71740 118318
rect 71688 118254 71740 118260
rect 73896 118312 73948 118318
rect 73896 118254 73948 118260
rect 82636 118312 82688 118318
rect 82636 118254 82688 118260
rect 71594 118008 71650 118017
rect 70216 117972 70268 117978
rect 73908 117978 73936 118254
rect 76010 118008 76066 118017
rect 71594 117943 71650 117952
rect 73896 117972 73948 117978
rect 70216 117914 70268 117920
rect 76010 117943 76066 117952
rect 73896 117914 73948 117920
rect 70228 117473 70256 117914
rect 70214 117464 70270 117473
rect 70214 117399 70270 117408
rect 73908 115938 73936 117914
rect 73896 115932 73948 115938
rect 73896 115874 73948 115880
rect 73896 108996 73948 109002
rect 73896 108938 73948 108944
rect 73908 106298 73936 108938
rect 73908 106270 74028 106298
rect 74000 99414 74028 106270
rect 73804 99408 73856 99414
rect 73804 99350 73856 99356
rect 73988 99408 74040 99414
rect 73988 99350 74040 99356
rect 73816 89894 73844 99350
rect 73804 89888 73856 89894
rect 73804 89830 73856 89836
rect 73712 87032 73764 87038
rect 73712 86974 73764 86980
rect 73724 79914 73752 86974
rect 73724 79886 73844 79914
rect 73816 66298 73844 79886
rect 73804 66292 73856 66298
rect 73804 66234 73856 66240
rect 73896 66292 73948 66298
rect 73896 66234 73948 66240
rect 73908 58002 73936 66234
rect 73896 57996 73948 58002
rect 73896 57938 73948 57944
rect 73988 57860 74040 57866
rect 73988 57802 74040 57808
rect 74000 48521 74028 57802
rect 73986 48512 74042 48521
rect 73986 48447 74042 48456
rect 73618 48376 73674 48385
rect 73618 48311 73674 48320
rect 73632 48278 73660 48311
rect 73620 48272 73672 48278
rect 73620 48214 73672 48220
rect 73804 35352 73856 35358
rect 73804 35294 73856 35300
rect 73816 34513 73844 35294
rect 73618 34504 73674 34513
rect 73618 34439 73674 34448
rect 73802 34504 73858 34513
rect 73802 34439 73858 34448
rect 73632 24886 73660 34439
rect 73620 24880 73672 24886
rect 73620 24822 73672 24828
rect 73896 24880 73948 24886
rect 73896 24822 73948 24828
rect 73908 20058 73936 24822
rect 73896 20052 73948 20058
rect 73896 19994 73948 20000
rect 74264 12368 74316 12374
rect 74264 12310 74316 12316
rect 68284 9512 68336 9518
rect 68284 9454 68336 9460
rect 67548 4208 67600 4214
rect 67548 4150 67600 4156
rect 67180 604 67232 610
rect 67180 546 67232 552
rect 67192 480 67220 546
rect 68296 480 68324 9454
rect 71872 6452 71924 6458
rect 71872 6394 71924 6400
rect 69480 5500 69532 5506
rect 69480 5442 69532 5448
rect 69492 480 69520 5442
rect 70676 4208 70728 4214
rect 70676 4150 70728 4156
rect 70688 480 70716 4150
rect 71884 480 71912 6394
rect 73068 4752 73120 4758
rect 73068 4694 73120 4700
rect 73080 480 73108 4694
rect 74276 480 74304 12310
rect 75460 9580 75512 9586
rect 75460 9522 75512 9528
rect 75472 480 75500 9522
rect 76024 3194 76052 117943
rect 77852 7336 77904 7342
rect 77852 7278 77904 7284
rect 76656 4684 76708 4690
rect 76656 4626 76708 4632
rect 76012 3188 76064 3194
rect 76012 3130 76064 3136
rect 76668 480 76696 4626
rect 77864 480 77892 7278
rect 79048 6520 79100 6526
rect 79048 6462 79100 6468
rect 79060 480 79088 6462
rect 80244 4616 80296 4622
rect 80244 4558 80296 4564
rect 80256 480 80284 4558
rect 82648 3482 82676 118254
rect 88352 118046 88380 118322
rect 88340 118040 88392 118046
rect 88340 117982 88392 117988
rect 87328 9648 87380 9654
rect 87328 9590 87380 9596
rect 84936 7268 84988 7274
rect 84936 7210 84988 7216
rect 83832 4548 83884 4554
rect 83832 4490 83884 4496
rect 82556 3454 82676 3482
rect 82556 3330 82584 3454
rect 81440 3324 81492 3330
rect 81440 3266 81492 3272
rect 82544 3324 82596 3330
rect 82544 3266 82596 3272
rect 82636 3324 82688 3330
rect 82636 3266 82688 3272
rect 81452 480 81480 3266
rect 82648 480 82676 3266
rect 83844 480 83872 4490
rect 84948 480 84976 7210
rect 86132 6588 86184 6594
rect 86132 6530 86184 6536
rect 86144 480 86172 6530
rect 87340 480 87368 9590
rect 88352 4842 88380 117982
rect 97920 117366 97948 118526
rect 100680 117609 100708 337350
rect 102888 336870 102916 340054
rect 107580 338094 107608 340054
rect 107568 338088 107620 338094
rect 107568 338030 107620 338036
rect 103428 337476 103480 337482
rect 103428 337418 103480 337424
rect 102876 336864 102928 336870
rect 102876 336806 102928 336812
rect 103336 336864 103388 336870
rect 103336 336806 103388 336812
rect 103348 202230 103376 336806
rect 103336 202224 103388 202230
rect 103336 202166 103388 202172
rect 103440 118561 103468 337418
rect 103426 118552 103482 118561
rect 103426 118487 103482 118496
rect 100666 117600 100722 117609
rect 100666 117535 100722 117544
rect 92388 117360 92440 117366
rect 92388 117302 92440 117308
rect 97908 117360 97960 117366
rect 100680 117337 100708 117535
rect 103440 117337 103468 118487
rect 107580 118250 107608 338030
rect 107568 118244 107620 118250
rect 107568 118186 107620 118192
rect 108304 118244 108356 118250
rect 108304 118186 108356 118192
rect 107580 117978 107608 118186
rect 107568 117972 107620 117978
rect 107568 117914 107620 117920
rect 97908 117302 97960 117308
rect 100022 117328 100078 117337
rect 89720 6724 89772 6730
rect 89720 6666 89772 6672
rect 88352 4814 88564 4842
rect 88536 480 88564 4814
rect 89732 480 89760 6666
rect 90916 6656 90968 6662
rect 90916 6598 90968 6604
rect 90928 480 90956 6598
rect 92400 2854 92428 117302
rect 100022 117263 100078 117272
rect 100666 117328 100722 117337
rect 100666 117263 100722 117272
rect 102138 117328 102194 117337
rect 102138 117263 102194 117272
rect 103426 117328 103482 117337
rect 103426 117263 103482 117272
rect 95700 7200 95752 7206
rect 95700 7142 95752 7148
rect 94504 6792 94556 6798
rect 94504 6734 94556 6740
rect 93308 3256 93360 3262
rect 93308 3198 93360 3204
rect 92112 2848 92164 2854
rect 92112 2790 92164 2796
rect 92388 2848 92440 2854
rect 92388 2790 92440 2796
rect 92124 480 92152 2790
rect 93320 480 93348 3198
rect 94516 480 94544 6734
rect 95712 480 95740 7142
rect 96896 6860 96948 6866
rect 96896 6802 96948 6808
rect 96908 480 96936 6802
rect 98092 6112 98144 6118
rect 98092 6054 98144 6060
rect 98104 480 98132 6054
rect 100036 3194 100064 117263
rect 101588 6044 101640 6050
rect 101588 5986 101640 5992
rect 99288 3188 99340 3194
rect 99288 3130 99340 3136
rect 100024 3188 100076 3194
rect 100024 3130 100076 3136
rect 100484 3188 100536 3194
rect 100484 3130 100536 3136
rect 99300 480 99328 3130
rect 100496 480 100524 3130
rect 101600 480 101628 5986
rect 102152 3482 102180 117263
rect 106372 8900 106424 8906
rect 106372 8842 106424 8848
rect 103980 5976 104032 5982
rect 103980 5918 104032 5924
rect 102152 3454 102824 3482
rect 102796 480 102824 3454
rect 103992 480 104020 5918
rect 105176 5908 105228 5914
rect 105176 5850 105228 5856
rect 105188 480 105216 5850
rect 106384 480 106412 8842
rect 108316 5846 108344 118186
rect 110340 118114 110368 340138
rect 111720 118182 111748 340206
rect 112516 340190 113128 340218
rect 113100 337958 113128 340190
rect 117668 340054 118004 340082
rect 122636 340054 122788 340082
rect 113088 337952 113140 337958
rect 113088 337894 113140 337900
rect 113100 118454 113128 337894
rect 117228 337680 117280 337686
rect 117228 337622 117280 337628
rect 113088 118448 113140 118454
rect 117240 118425 117268 337622
rect 117976 337550 118004 340054
rect 122760 337890 122788 340054
rect 122748 337884 122800 337890
rect 122748 337826 122800 337832
rect 117964 337544 118016 337550
rect 117964 337486 118016 337492
rect 113088 118390 113140 118396
rect 117226 118416 117282 118425
rect 111708 118176 111760 118182
rect 111708 118118 111760 118124
rect 110328 118108 110380 118114
rect 110328 118050 110380 118056
rect 110340 117881 110368 118050
rect 110326 117872 110382 117881
rect 110326 117807 110382 117816
rect 111720 117434 111748 118118
rect 113100 118114 113128 118390
rect 117226 118351 117282 118360
rect 113088 118108 113140 118114
rect 113088 118050 113140 118056
rect 111708 117428 111760 117434
rect 111708 117370 111760 117376
rect 117240 117337 117268 118351
rect 122104 117904 122156 117910
rect 122104 117846 122156 117852
rect 122564 117904 122616 117910
rect 122760 117858 122788 337826
rect 125704 118114 125732 394454
rect 125784 394392 125836 394398
rect 125784 394334 125836 394340
rect 125796 118289 125824 394334
rect 125888 118318 125916 395626
rect 125980 336734 126008 395814
rect 126058 395720 126114 395729
rect 126058 395655 126114 395664
rect 126072 340134 126100 395655
rect 126164 394398 126192 397394
rect 126152 394392 126204 394398
rect 126152 394334 126204 394340
rect 126060 340128 126112 340134
rect 126060 340070 126112 340076
rect 125968 336728 126020 336734
rect 125968 336670 126020 336676
rect 126256 144430 126284 700334
rect 130384 583568 130436 583574
rect 130384 583510 130436 583516
rect 129004 583500 129056 583506
rect 129004 583442 129056 583448
rect 128360 553852 128412 553858
rect 128360 553794 128412 553800
rect 127716 518832 127768 518838
rect 127716 518774 127768 518780
rect 126336 518424 126388 518430
rect 126336 518366 126388 518372
rect 126348 497962 126376 518366
rect 126980 518220 127032 518226
rect 126980 518162 127032 518168
rect 126336 497956 126388 497962
rect 126336 497898 126388 497904
rect 126348 496874 126376 497898
rect 126336 496868 126388 496874
rect 126336 496810 126388 496816
rect 126888 496868 126940 496874
rect 126888 496810 126940 496816
rect 126426 417480 126482 417489
rect 126426 417415 126482 417424
rect 126336 397520 126388 397526
rect 126336 397462 126388 397468
rect 126348 201618 126376 397462
rect 126440 337686 126468 417415
rect 126520 396840 126572 396846
rect 126520 396782 126572 396788
rect 126532 358766 126560 396782
rect 126900 395729 126928 496810
rect 126886 395720 126942 395729
rect 126886 395655 126942 395664
rect 126520 358760 126572 358766
rect 126520 358702 126572 358708
rect 126888 340740 126940 340746
rect 126888 340682 126940 340688
rect 126900 340134 126928 340682
rect 126888 340128 126940 340134
rect 126888 340070 126940 340076
rect 126428 337680 126480 337686
rect 126428 337622 126480 337628
rect 126336 201612 126388 201618
rect 126336 201554 126388 201560
rect 126244 144424 126296 144430
rect 126244 144366 126296 144372
rect 126900 118402 126928 340070
rect 126992 338026 127020 518162
rect 127072 497548 127124 497554
rect 127072 497490 127124 497496
rect 126980 338020 127032 338026
rect 126980 337962 127032 337968
rect 127084 337958 127112 497490
rect 127256 398132 127308 398138
rect 127256 398074 127308 398080
rect 127164 397792 127216 397798
rect 127164 397734 127216 397740
rect 127176 340882 127204 397734
rect 127164 340876 127216 340882
rect 127164 340818 127216 340824
rect 127176 340270 127204 340818
rect 127268 340814 127296 398074
rect 127624 397724 127676 397730
rect 127624 397666 127676 397672
rect 127256 340808 127308 340814
rect 127256 340750 127308 340756
rect 127164 340264 127216 340270
rect 127164 340206 127216 340212
rect 127268 340202 127296 340750
rect 127256 340196 127308 340202
rect 127256 340138 127308 340144
rect 127072 337952 127124 337958
rect 127072 337894 127124 337900
rect 127636 201550 127664 397666
rect 127728 340610 127756 518774
rect 128268 396772 128320 396778
rect 128268 396714 128320 396720
rect 127716 340604 127768 340610
rect 127716 340546 127768 340552
rect 127728 337890 127756 340546
rect 127716 337884 127768 337890
rect 127716 337826 127768 337832
rect 127624 201544 127676 201550
rect 127624 201486 127676 201492
rect 128176 144764 128228 144770
rect 128176 144706 128228 144712
rect 128188 144537 128216 144706
rect 128174 144528 128230 144537
rect 128174 144463 128230 144472
rect 126900 118374 127020 118402
rect 125876 118312 125928 118318
rect 125782 118280 125838 118289
rect 125876 118254 125928 118260
rect 126888 118312 126940 118318
rect 126888 118254 126940 118260
rect 125782 118215 125838 118224
rect 126244 118244 126296 118250
rect 125692 118108 125744 118114
rect 125692 118050 125744 118056
rect 125796 117994 125824 118215
rect 126244 118186 126296 118192
rect 122616 117852 122788 117858
rect 122564 117846 122788 117852
rect 120724 117768 120776 117774
rect 120724 117710 120776 117716
rect 115938 117328 115994 117337
rect 115938 117263 115994 117272
rect 117226 117328 117282 117337
rect 117226 117263 117282 117272
rect 115952 7546 115980 117263
rect 119436 8832 119488 8838
rect 119436 8774 119488 8780
rect 115940 7540 115992 7546
rect 115940 7482 115992 7488
rect 117136 7540 117188 7546
rect 117136 7482 117188 7488
rect 118240 7540 118292 7546
rect 118240 7482 118292 7488
rect 109960 7132 110012 7138
rect 109960 7074 110012 7080
rect 108304 5840 108356 5846
rect 108304 5782 108356 5788
rect 108764 5840 108816 5846
rect 108764 5782 108816 5788
rect 107568 3120 107620 3126
rect 107568 3062 107620 3068
rect 107580 480 107608 3062
rect 108776 480 108804 5782
rect 109972 480 110000 7074
rect 113546 6216 113602 6225
rect 113546 6151 113602 6160
rect 112352 5772 112404 5778
rect 112352 5714 112404 5720
rect 111156 5704 111208 5710
rect 111156 5646 111208 5652
rect 111168 480 111196 5646
rect 112364 480 112392 5714
rect 113560 480 113588 6151
rect 115940 5636 115992 5642
rect 115940 5578 115992 5584
rect 114744 3052 114796 3058
rect 114744 2994 114796 3000
rect 114756 480 114784 2994
rect 115952 480 115980 5578
rect 117148 480 117176 7482
rect 118252 480 118280 7482
rect 119448 480 119476 8774
rect 120632 8764 120684 8770
rect 120632 8706 120684 8712
rect 120644 480 120672 8706
rect 120736 4214 120764 117710
rect 121828 7472 121880 7478
rect 121828 7414 121880 7420
rect 120724 4208 120776 4214
rect 120724 4150 120776 4156
rect 121840 480 121868 7414
rect 122116 4350 122144 117846
rect 122576 117830 122788 117846
rect 125520 117966 125824 117994
rect 123024 5568 123076 5574
rect 123024 5510 123076 5516
rect 122104 4344 122156 4350
rect 122104 4286 122156 4292
rect 123036 480 123064 5510
rect 125520 2990 125548 117966
rect 126256 4418 126284 118186
rect 126900 117774 126928 118254
rect 126992 118250 127020 118374
rect 126980 118244 127032 118250
rect 126980 118186 127032 118192
rect 126992 118114 127020 118186
rect 126980 118108 127032 118114
rect 126980 118050 127032 118056
rect 126888 117768 126940 117774
rect 128280 117745 128308 396714
rect 128372 358329 128400 553794
rect 128728 525088 128780 525094
rect 128728 525030 128780 525036
rect 128740 524822 128768 525030
rect 128728 524816 128780 524822
rect 128728 524758 128780 524764
rect 128452 521620 128504 521626
rect 128452 521562 128504 521568
rect 128464 521014 128492 521562
rect 128452 521008 128504 521014
rect 128452 520950 128504 520956
rect 128464 373289 128492 520950
rect 128740 509266 128768 524758
rect 129016 521626 129044 583442
rect 129280 583432 129332 583438
rect 129280 583374 129332 583380
rect 129188 578264 129240 578270
rect 129188 578206 129240 578212
rect 129096 553716 129148 553722
rect 129096 553658 129148 553664
rect 129004 521620 129056 521626
rect 129004 521562 129056 521568
rect 128648 509238 128768 509266
rect 128648 505102 128676 509238
rect 128636 505096 128688 505102
rect 128636 505038 128688 505044
rect 128820 505096 128872 505102
rect 128820 505038 128872 505044
rect 128832 495394 128860 505038
rect 129108 498166 129136 553658
rect 129200 524822 129228 578206
rect 129292 553858 129320 583374
rect 129648 563100 129700 563106
rect 129648 563042 129700 563048
rect 129280 553852 129332 553858
rect 129280 553794 129332 553800
rect 129188 524816 129240 524822
rect 129188 524758 129240 524764
rect 129554 500168 129610 500177
rect 129554 500103 129610 500112
rect 129096 498160 129148 498166
rect 129096 498102 129148 498108
rect 128740 495366 128860 495394
rect 128740 491298 128768 495366
rect 128636 491292 128688 491298
rect 128636 491234 128688 491240
rect 128728 491292 128780 491298
rect 128728 491234 128780 491240
rect 128648 481681 128676 491234
rect 128634 481672 128690 481681
rect 128634 481607 128690 481616
rect 128818 481672 128874 481681
rect 128818 481607 128874 481616
rect 128832 476082 128860 481607
rect 128740 476054 128860 476082
rect 128740 468466 128768 476054
rect 128556 468438 128768 468466
rect 128556 463729 128584 468438
rect 128542 463720 128598 463729
rect 128542 463655 128598 463664
rect 128818 463720 128874 463729
rect 128818 463655 128874 463664
rect 128832 456770 128860 463655
rect 128740 456742 128860 456770
rect 128740 449154 128768 456742
rect 128556 449126 128768 449154
rect 128556 444417 128584 449126
rect 128542 444408 128598 444417
rect 128542 444343 128598 444352
rect 128818 444408 128874 444417
rect 128818 444343 128874 444352
rect 128832 437458 128860 444343
rect 128740 437430 128860 437458
rect 128740 429842 128768 437430
rect 128556 429814 128768 429842
rect 128556 425105 128584 429814
rect 128542 425096 128598 425105
rect 128542 425031 128598 425040
rect 128818 425096 128874 425105
rect 128818 425031 128874 425040
rect 128832 418146 128860 425031
rect 128648 418118 128860 418146
rect 128648 415410 128676 418118
rect 128636 415404 128688 415410
rect 128636 415346 128688 415352
rect 128544 405748 128596 405754
rect 128544 405690 128596 405696
rect 128556 405618 128584 405690
rect 128544 405612 128596 405618
rect 128544 405554 128596 405560
rect 128636 398744 128688 398750
rect 128636 398686 128688 398692
rect 128648 388249 128676 398686
rect 128634 388240 128690 388249
rect 128634 388175 128690 388184
rect 128648 386442 128676 388175
rect 128636 386436 128688 386442
rect 128636 386378 128688 386384
rect 128912 386436 128964 386442
rect 128912 386378 128964 386384
rect 128924 376961 128952 386378
rect 129108 380633 129136 498102
rect 129464 398200 129516 398206
rect 129464 398142 129516 398148
rect 129476 397594 129504 398142
rect 129464 397588 129516 397594
rect 129464 397530 129516 397536
rect 129094 380624 129150 380633
rect 129094 380559 129150 380568
rect 128910 376952 128966 376961
rect 128910 376887 128966 376896
rect 128818 376816 128874 376825
rect 128818 376751 128874 376760
rect 128832 375358 128860 376751
rect 128820 375352 128872 375358
rect 128820 375294 128872 375300
rect 128450 373280 128506 373289
rect 128450 373215 128506 373224
rect 128820 365764 128872 365770
rect 128820 365706 128872 365712
rect 128358 358320 128414 358329
rect 128358 358255 128414 358264
rect 128832 347750 128860 365706
rect 128912 358760 128964 358766
rect 128912 358702 128964 358708
rect 128820 347744 128872 347750
rect 128820 347686 128872 347692
rect 128818 343632 128874 343641
rect 128818 343567 128874 343576
rect 128832 342514 128860 343567
rect 128820 342508 128872 342514
rect 128820 342450 128872 342456
rect 128924 342122 128952 358702
rect 129004 351008 129056 351014
rect 129002 350976 129004 350985
rect 129056 350976 129058 350985
rect 129002 350911 129058 350920
rect 128832 342094 128952 342122
rect 128832 340678 128860 342094
rect 128820 340672 128872 340678
rect 128820 340614 128872 340620
rect 128832 338042 128860 340614
rect 128912 340536 128964 340542
rect 128912 340478 128964 340484
rect 128740 338014 128860 338042
rect 128924 338026 128952 340478
rect 128912 338020 128964 338026
rect 128740 331294 128768 338014
rect 128912 337962 128964 337968
rect 129004 332376 129056 332382
rect 129004 332318 129056 332324
rect 128728 331288 128780 331294
rect 128728 331230 128780 331236
rect 128728 328500 128780 328506
rect 128728 328442 128780 328448
rect 128740 321586 128768 328442
rect 128648 321558 128768 321586
rect 128648 321450 128676 321558
rect 128648 321422 128768 321450
rect 128740 318782 128768 321422
rect 128636 318776 128688 318782
rect 128636 318718 128688 318724
rect 128728 318776 128780 318782
rect 128728 318718 128780 318724
rect 128648 317422 128676 318718
rect 128636 317416 128688 317422
rect 128636 317358 128688 317364
rect 128728 309188 128780 309194
rect 128728 309130 128780 309136
rect 128740 307766 128768 309130
rect 128728 307760 128780 307766
rect 128728 307702 128780 307708
rect 128728 302184 128780 302190
rect 128728 302126 128780 302132
rect 128740 298110 128768 302126
rect 128728 298104 128780 298110
rect 128728 298046 128780 298052
rect 128728 292460 128780 292466
rect 128728 292402 128780 292408
rect 128740 288402 128768 292402
rect 128648 288374 128768 288402
rect 128648 282946 128676 288374
rect 128636 282940 128688 282946
rect 128636 282882 128688 282888
rect 128636 278792 128688 278798
rect 128636 278734 128688 278740
rect 128648 273358 128676 278734
rect 128636 273352 128688 273358
rect 128636 273294 128688 273300
rect 128636 270496 128688 270502
rect 128636 270438 128688 270444
rect 128648 260794 128676 270438
rect 128648 260766 128768 260794
rect 128740 259418 128768 260766
rect 128728 259412 128780 259418
rect 128728 259354 128780 259360
rect 128636 241596 128688 241602
rect 128636 241538 128688 241544
rect 128648 240122 128676 241538
rect 128648 240094 128768 240122
rect 128740 234666 128768 240094
rect 128728 234660 128780 234666
rect 128728 234602 128780 234608
rect 128636 234592 128688 234598
rect 128636 234534 128688 234540
rect 128648 220810 128676 234534
rect 128556 220782 128676 220810
rect 128556 196042 128584 220782
rect 129016 215370 129044 332318
rect 128832 215342 129044 215370
rect 128832 215234 128860 215342
rect 128832 215206 128952 215234
rect 128924 205714 128952 215206
rect 128924 205686 129044 205714
rect 128544 196036 128596 196042
rect 128544 195978 128596 195984
rect 128636 195900 128688 195906
rect 128636 195842 128688 195848
rect 128648 191758 128676 195842
rect 129016 191758 129044 205686
rect 128636 191752 128688 191758
rect 128636 191694 128688 191700
rect 129004 191752 129056 191758
rect 129004 191694 129056 191700
rect 128636 186244 128688 186250
rect 128636 186186 128688 186192
rect 128648 182186 128676 186186
rect 129004 183932 129056 183938
rect 129004 183874 129056 183880
rect 129016 182209 129044 183874
rect 128818 182200 128874 182209
rect 128648 182158 128768 182186
rect 128740 182102 128768 182158
rect 128818 182135 128820 182144
rect 128872 182135 128874 182144
rect 129002 182200 129058 182209
rect 129002 182135 129058 182144
rect 128820 182106 128872 182112
rect 128728 182096 128780 182102
rect 128728 182038 128780 182044
rect 128912 182096 128964 182102
rect 128912 182038 128964 182044
rect 128636 172576 128688 172582
rect 128636 172518 128688 172524
rect 128648 166954 128676 172518
rect 128924 167074 128952 182038
rect 128912 167068 128964 167074
rect 128912 167010 128964 167016
rect 128648 166926 128768 166954
rect 128740 164218 128768 166926
rect 128912 166932 128964 166938
rect 128912 166874 128964 166880
rect 128636 164212 128688 164218
rect 128636 164154 128688 164160
rect 128728 164212 128780 164218
rect 128728 164154 128780 164160
rect 128648 162858 128676 164154
rect 128636 162852 128688 162858
rect 128636 162794 128688 162800
rect 128924 153377 128952 166874
rect 128910 153368 128966 153377
rect 128910 153303 128966 153312
rect 128636 153264 128688 153270
rect 128636 153206 128688 153212
rect 128818 153232 128874 153241
rect 128648 147762 128676 153206
rect 128874 153176 128952 153184
rect 128818 153167 128952 153176
rect 128832 153156 128952 153167
rect 128636 147756 128688 147762
rect 128636 147698 128688 147704
rect 128636 147552 128688 147558
rect 128636 147494 128688 147500
rect 128648 132870 128676 147494
rect 128924 144974 128952 153156
rect 128912 144968 128964 144974
rect 128912 144910 128964 144916
rect 128820 144900 128872 144906
rect 128820 144842 128872 144848
rect 128832 143562 128860 144842
rect 128832 143534 128952 143562
rect 128924 135425 128952 143534
rect 128910 135416 128966 135425
rect 128910 135351 128966 135360
rect 128818 135280 128874 135289
rect 128818 135215 128874 135224
rect 128832 135130 128860 135215
rect 128832 135102 128952 135130
rect 128636 132864 128688 132870
rect 128636 132806 128688 132812
rect 128820 132864 128872 132870
rect 128820 132806 128872 132812
rect 128728 118720 128780 118726
rect 128832 118697 128860 132806
rect 128924 118726 128952 135102
rect 128912 118720 128964 118726
rect 128728 118662 128780 118668
rect 128818 118688 128874 118697
rect 128740 118130 128768 118662
rect 128912 118662 128964 118668
rect 128818 118623 128874 118632
rect 128740 118102 128952 118130
rect 128924 117978 128952 118102
rect 128912 117972 128964 117978
rect 128912 117914 128964 117920
rect 126888 117710 126940 117716
rect 127622 117736 127678 117745
rect 127622 117671 127678 117680
rect 128266 117736 128322 117745
rect 128266 117671 128322 117680
rect 127636 8226 127664 117671
rect 128924 91746 128952 117914
rect 129108 117774 129136 380559
rect 129186 373280 129242 373289
rect 129186 373215 129242 373224
rect 129200 118250 129228 373215
rect 129370 365936 129426 365945
rect 129370 365871 129426 365880
rect 129384 365702 129412 365871
rect 129372 365696 129424 365702
rect 129372 365638 129424 365644
rect 129278 358320 129334 358329
rect 129278 358255 129334 358264
rect 129292 118318 129320 358255
rect 129280 118312 129332 118318
rect 129280 118254 129332 118260
rect 129188 118244 129240 118250
rect 129188 118186 129240 118192
rect 129096 117768 129148 117774
rect 129096 117710 129148 117716
rect 128740 91718 128952 91746
rect 128740 87009 128768 91718
rect 128726 87000 128782 87009
rect 128726 86935 128782 86944
rect 129002 87000 129058 87009
rect 129002 86935 129058 86944
rect 129016 77314 129044 86935
rect 128820 77308 128872 77314
rect 128820 77250 128872 77256
rect 129004 77308 129056 77314
rect 129004 77250 129056 77256
rect 128832 77194 128860 77250
rect 128740 77166 128860 77194
rect 128740 67726 128768 77166
rect 128728 67720 128780 67726
rect 128728 67662 128780 67668
rect 128912 67652 128964 67658
rect 128912 67594 128964 67600
rect 128924 66230 128952 67594
rect 128912 66224 128964 66230
rect 128912 66166 128964 66172
rect 129004 57860 129056 57866
rect 129004 57802 129056 57808
rect 129016 50946 129044 57802
rect 128924 50918 129044 50946
rect 128924 41426 128952 50918
rect 128924 41398 129044 41426
rect 129016 38622 129044 41398
rect 129004 38616 129056 38622
rect 129004 38558 129056 38564
rect 128912 29028 128964 29034
rect 128912 28970 128964 28976
rect 128924 22114 128952 28970
rect 128924 22086 129044 22114
rect 129016 12458 129044 22086
rect 128832 12430 129044 12458
rect 127624 8220 127676 8226
rect 127624 8162 127676 8168
rect 127808 8220 127860 8226
rect 127808 8162 127860 8168
rect 126612 7404 126664 7410
rect 126612 7346 126664 7352
rect 126244 4412 126296 4418
rect 126244 4354 126296 4360
rect 124220 2984 124272 2990
rect 124220 2926 124272 2932
rect 125508 2984 125560 2990
rect 125508 2926 125560 2932
rect 124232 480 124260 2926
rect 125416 2916 125468 2922
rect 125416 2858 125468 2864
rect 125428 480 125456 2858
rect 126624 480 126652 7346
rect 127820 480 127848 8162
rect 128832 4282 128860 12430
rect 129004 7336 129056 7342
rect 129004 7278 129056 7284
rect 128820 4276 128872 4282
rect 128820 4218 128872 4224
rect 129016 480 129044 7278
rect 129108 7274 129136 117710
rect 129096 7268 129148 7274
rect 129096 7210 129148 7216
rect 129200 7206 129228 118186
rect 129188 7200 129240 7206
rect 129188 7142 129240 7148
rect 129292 7070 129320 118254
rect 129384 117502 129412 365638
rect 129476 117570 129504 397530
rect 129568 118726 129596 500103
rect 129660 118862 129688 563042
rect 130396 518906 130424 583510
rect 131026 582448 131082 582457
rect 131026 582383 131082 582392
rect 130384 518900 130436 518906
rect 130384 518842 130436 518848
rect 130396 407182 130424 518842
rect 130934 500304 130990 500313
rect 130934 500239 130990 500248
rect 130384 407176 130436 407182
rect 130384 407118 130436 407124
rect 130396 351014 130424 407118
rect 130384 351008 130436 351014
rect 130384 350950 130436 350956
rect 129648 118856 129700 118862
rect 129648 118798 129700 118804
rect 129556 118720 129608 118726
rect 129556 118662 129608 118668
rect 129648 118108 129700 118114
rect 129648 118050 129700 118056
rect 129660 117978 129688 118050
rect 129648 117972 129700 117978
rect 129648 117914 129700 117920
rect 130396 117638 130424 350950
rect 130842 196208 130898 196217
rect 130842 196143 130898 196152
rect 130856 196110 130884 196143
rect 130844 196104 130896 196110
rect 130844 196046 130896 196052
rect 130842 194712 130898 194721
rect 130842 194647 130844 194656
rect 130896 194647 130898 194656
rect 130844 194618 130896 194624
rect 130844 194540 130896 194546
rect 130844 194482 130896 194488
rect 130856 194449 130884 194482
rect 130842 194440 130898 194449
rect 130842 194375 130898 194384
rect 130752 193180 130804 193186
rect 130752 193122 130804 193128
rect 130764 192545 130792 193122
rect 130844 193112 130896 193118
rect 130842 193080 130844 193089
rect 130896 193080 130898 193089
rect 130842 193015 130898 193024
rect 130750 192536 130806 192545
rect 130750 192471 130806 192480
rect 130844 191820 130896 191826
rect 130844 191762 130896 191768
rect 130856 191457 130884 191762
rect 130842 191448 130898 191457
rect 130842 191383 130898 191392
rect 130844 190460 130896 190466
rect 130844 190402 130896 190408
rect 130856 190369 130884 190402
rect 130842 190360 130898 190369
rect 130842 190295 130898 190304
rect 130752 189032 130804 189038
rect 130752 188974 130804 188980
rect 130842 189000 130898 189009
rect 130764 188329 130792 188974
rect 130842 188935 130844 188944
rect 130896 188935 130898 188944
rect 130844 188906 130896 188912
rect 130750 188320 130806 188329
rect 130750 188255 130806 188264
rect 130844 187672 130896 187678
rect 130844 187614 130896 187620
rect 130856 187241 130884 187614
rect 130842 187232 130898 187241
rect 130842 187167 130898 187176
rect 130948 118930 130976 500239
rect 130936 118924 130988 118930
rect 130936 118866 130988 118872
rect 131040 118794 131068 582383
rect 131132 156330 131160 700674
rect 131212 700596 131264 700602
rect 131212 700538 131264 700544
rect 131224 186318 131252 700538
rect 132316 700528 132368 700534
rect 132316 700470 132368 700476
rect 132132 498228 132184 498234
rect 132132 498170 132184 498176
rect 131948 341692 132000 341698
rect 131948 341634 132000 341640
rect 131672 341556 131724 341562
rect 131672 341498 131724 341504
rect 131580 263628 131632 263634
rect 131580 263570 131632 263576
rect 131304 227792 131356 227798
rect 131304 227734 131356 227740
rect 131212 186312 131264 186318
rect 131212 186254 131264 186260
rect 131212 186176 131264 186182
rect 131212 186118 131264 186124
rect 131224 185609 131252 186118
rect 131210 185600 131266 185609
rect 131210 185535 131266 185544
rect 131212 184884 131264 184890
rect 131212 184826 131264 184832
rect 131224 184521 131252 184826
rect 131210 184512 131266 184521
rect 131210 184447 131266 184456
rect 131210 183560 131266 183569
rect 131210 183495 131212 183504
rect 131264 183495 131266 183504
rect 131212 183466 131264 183472
rect 131212 183388 131264 183394
rect 131212 183330 131264 183336
rect 131224 178265 131252 183330
rect 131210 178256 131266 178265
rect 131210 178191 131266 178200
rect 131316 164529 131344 227734
rect 131488 216708 131540 216714
rect 131488 216650 131540 216656
rect 131396 200796 131448 200802
rect 131396 200738 131448 200744
rect 131408 198354 131436 200738
rect 131396 198348 131448 198354
rect 131396 198290 131448 198296
rect 131394 198248 131450 198257
rect 131394 198183 131450 198192
rect 131408 197402 131436 198183
rect 131396 197396 131448 197402
rect 131396 197338 131448 197344
rect 131394 197160 131450 197169
rect 131394 197095 131450 197104
rect 131408 196314 131436 197095
rect 131396 196308 131448 196314
rect 131396 196250 131448 196256
rect 131396 196036 131448 196042
rect 131396 195978 131448 195984
rect 131302 164520 131358 164529
rect 131302 164455 131358 164464
rect 131302 157176 131358 157185
rect 131302 157111 131358 157120
rect 131120 156324 131172 156330
rect 131120 156266 131172 156272
rect 131118 156224 131174 156233
rect 131118 156159 131174 156168
rect 131132 156058 131160 156159
rect 131316 156126 131344 157111
rect 131304 156120 131356 156126
rect 131304 156062 131356 156068
rect 131120 156052 131172 156058
rect 131120 155994 131172 156000
rect 131304 155984 131356 155990
rect 131304 155926 131356 155932
rect 131120 155916 131172 155922
rect 131120 155858 131172 155864
rect 131132 155145 131160 155858
rect 131118 155136 131174 155145
rect 131118 155071 131174 155080
rect 131212 155100 131264 155106
rect 131212 155042 131264 155048
rect 131120 154420 131172 154426
rect 131120 154362 131172 154368
rect 131132 154057 131160 154362
rect 131118 154048 131174 154057
rect 131118 153983 131174 153992
rect 131120 153196 131172 153202
rect 131120 153138 131172 153144
rect 131132 152969 131160 153138
rect 131118 152960 131174 152969
rect 131118 152895 131174 152904
rect 131120 151768 131172 151774
rect 131120 151710 131172 151716
rect 131132 150929 131160 151710
rect 131118 150920 131174 150929
rect 131118 150855 131174 150864
rect 131120 150408 131172 150414
rect 131120 150350 131172 150356
rect 131132 149841 131160 150350
rect 131118 149832 131174 149841
rect 131118 149767 131174 149776
rect 131120 148980 131172 148986
rect 131120 148922 131172 148928
rect 131132 148753 131160 148922
rect 131118 148744 131174 148753
rect 131118 148679 131174 148688
rect 131120 148640 131172 148646
rect 131120 148582 131172 148588
rect 131132 147801 131160 148582
rect 131118 147792 131174 147801
rect 131118 147727 131174 147736
rect 131224 147626 131252 155042
rect 131316 153134 131344 155926
rect 131304 153128 131356 153134
rect 131304 153070 131356 153076
rect 131304 152992 131356 152998
rect 131304 152934 131356 152940
rect 131316 152017 131344 152934
rect 131302 152008 131358 152017
rect 131302 151943 131358 151952
rect 131304 151904 131356 151910
rect 131304 151846 131356 151852
rect 131212 147620 131264 147626
rect 131212 147562 131264 147568
rect 131212 147484 131264 147490
rect 131212 147426 131264 147432
rect 131224 146713 131252 147426
rect 131210 146704 131266 146713
rect 131210 146639 131266 146648
rect 131120 146260 131172 146266
rect 131120 146202 131172 146208
rect 131132 145625 131160 146202
rect 131118 145616 131174 145625
rect 131118 145551 131174 145560
rect 131120 144424 131172 144430
rect 131120 144366 131172 144372
rect 131132 143585 131160 144366
rect 131118 143576 131174 143585
rect 131118 143511 131174 143520
rect 131316 139369 131344 151846
rect 131302 139360 131358 139369
rect 131302 139295 131358 139304
rect 131212 132524 131264 132530
rect 131212 132466 131264 132472
rect 131224 125662 131252 132466
rect 131408 132025 131436 195978
rect 131394 132016 131450 132025
rect 131394 131951 131450 131960
rect 131120 125656 131172 125662
rect 131120 125598 131172 125604
rect 131212 125656 131264 125662
rect 131212 125598 131264 125604
rect 131132 124166 131160 125598
rect 131500 124545 131528 216650
rect 131592 125633 131620 263570
rect 131684 167793 131712 341498
rect 131856 310548 131908 310554
rect 131856 310490 131908 310496
rect 131762 199336 131818 199345
rect 131762 199271 131818 199280
rect 131776 196110 131804 199271
rect 131764 196104 131816 196110
rect 131764 196046 131816 196052
rect 131764 195968 131816 195974
rect 131764 195910 131816 195916
rect 131670 167784 131726 167793
rect 131670 167719 131726 167728
rect 131670 158264 131726 158273
rect 131670 158199 131726 158208
rect 131578 125624 131634 125633
rect 131578 125559 131634 125568
rect 131486 124536 131542 124545
rect 131486 124471 131542 124480
rect 131120 124160 131172 124166
rect 131120 124102 131172 124108
rect 131028 118788 131080 118794
rect 131028 118730 131080 118736
rect 130384 117632 130436 117638
rect 130384 117574 130436 117580
rect 129464 117564 129516 117570
rect 129464 117506 129516 117512
rect 129372 117496 129424 117502
rect 129372 117438 129424 117444
rect 130200 7268 130252 7274
rect 130200 7210 130252 7216
rect 129280 7064 129332 7070
rect 129280 7006 129332 7012
rect 130212 480 130240 7210
rect 130396 4486 130424 117574
rect 131212 114572 131264 114578
rect 131212 114514 131264 114520
rect 131224 109018 131252 114514
rect 131224 108990 131344 109018
rect 131316 106282 131344 108990
rect 131304 106276 131356 106282
rect 131304 106218 131356 106224
rect 131304 99340 131356 99346
rect 131304 99282 131356 99288
rect 131316 96642 131344 99282
rect 131316 96614 131436 96642
rect 131408 88330 131436 96614
rect 131396 88324 131448 88330
rect 131396 88266 131448 88272
rect 131684 64870 131712 158199
rect 131672 64864 131724 64870
rect 131672 64806 131724 64812
rect 131776 8294 131804 195910
rect 131868 126721 131896 310490
rect 131960 128761 131988 341634
rect 132040 341624 132092 341630
rect 132040 341566 132092 341572
rect 131946 128752 132002 128761
rect 131946 128687 132002 128696
rect 132052 127809 132080 341566
rect 132144 130937 132172 498170
rect 132224 200864 132276 200870
rect 132224 200806 132276 200812
rect 132236 170921 132264 200806
rect 132222 170912 132278 170921
rect 132222 170847 132278 170856
rect 132222 159352 132278 159361
rect 132222 159287 132278 159296
rect 132130 130928 132186 130937
rect 132130 130863 132186 130872
rect 132038 127800 132094 127809
rect 132038 127735 132094 127744
rect 131854 126712 131910 126721
rect 131854 126647 131910 126656
rect 132130 121408 132186 121417
rect 132130 121343 132186 121352
rect 132144 77246 132172 121343
rect 132132 77240 132184 77246
rect 132132 77182 132184 77188
rect 132236 22098 132264 159287
rect 132328 138281 132356 700470
rect 132408 200932 132460 200938
rect 132408 200874 132460 200880
rect 132420 172009 132448 200874
rect 132512 179353 132540 700810
rect 133696 700800 133748 700806
rect 133696 700742 133748 700748
rect 132592 700392 132644 700398
rect 132592 700334 132644 700340
rect 132498 179344 132554 179353
rect 132498 179279 132554 179288
rect 132604 177177 132632 700334
rect 133420 700256 133472 700262
rect 133420 700198 133472 700204
rect 133328 699712 133380 699718
rect 133328 699654 133380 699660
rect 133144 462392 133196 462398
rect 133144 462334 133196 462340
rect 133052 415472 133104 415478
rect 133052 415414 133104 415420
rect 132960 342916 133012 342922
rect 132960 342858 133012 342864
rect 132972 342514 133000 342858
rect 132960 342508 133012 342514
rect 132960 342450 133012 342456
rect 132684 337544 132736 337550
rect 132684 337486 132736 337492
rect 132696 308310 132724 337486
rect 132776 321632 132828 321638
rect 132776 321574 132828 321580
rect 132684 308304 132736 308310
rect 132684 308246 132736 308252
rect 132684 274712 132736 274718
rect 132684 274654 132736 274660
rect 132590 177168 132646 177177
rect 132590 177103 132646 177112
rect 132406 172000 132462 172009
rect 132406 171935 132462 171944
rect 132696 165617 132724 274654
rect 132788 166705 132816 321574
rect 132868 308304 132920 308310
rect 132868 308246 132920 308252
rect 132880 196110 132908 308246
rect 132868 196104 132920 196110
rect 132868 196046 132920 196052
rect 132868 195968 132920 195974
rect 132868 195910 132920 195916
rect 132880 181490 132908 195910
rect 132868 181484 132920 181490
rect 132868 181426 132920 181432
rect 132774 166696 132830 166705
rect 132774 166631 132830 166640
rect 132682 165608 132738 165617
rect 132682 165543 132738 165552
rect 132592 164756 132644 164762
rect 132592 164698 132644 164704
rect 132604 164218 132632 164698
rect 132592 164212 132644 164218
rect 132592 164154 132644 164160
rect 132776 164144 132828 164150
rect 132776 164086 132828 164092
rect 132406 162480 132462 162489
rect 132406 162415 132462 162424
rect 132314 138272 132370 138281
rect 132314 138207 132370 138216
rect 132420 121174 132448 162415
rect 132682 161392 132738 161401
rect 132682 161327 132738 161336
rect 132696 155106 132724 161327
rect 132684 155100 132736 155106
rect 132684 155042 132736 155048
rect 132788 154986 132816 164086
rect 132696 154958 132816 154986
rect 132696 142118 132724 154958
rect 132684 142112 132736 142118
rect 132684 142054 132736 142060
rect 132776 135244 132828 135250
rect 132776 135186 132828 135192
rect 132788 132462 132816 135186
rect 132776 132456 132828 132462
rect 132776 132398 132828 132404
rect 132408 121168 132460 121174
rect 132408 121110 132460 121116
rect 132406 120456 132462 120465
rect 132406 120391 132462 120400
rect 132420 30326 132448 120391
rect 132972 117298 133000 342450
rect 133064 168745 133092 415414
rect 133156 169833 133184 462334
rect 133236 451308 133288 451314
rect 133236 451250 133288 451256
rect 133142 169824 133198 169833
rect 133142 169759 133198 169768
rect 133050 168736 133106 168745
rect 133050 168671 133106 168680
rect 133248 129849 133276 451250
rect 133340 182481 133368 699654
rect 133326 182472 133382 182481
rect 133326 182407 133382 182416
rect 133328 181484 133380 181490
rect 133328 181426 133380 181432
rect 133340 164762 133368 181426
rect 133432 181393 133460 700198
rect 133512 201204 133564 201210
rect 133512 201146 133564 201152
rect 133418 181384 133474 181393
rect 133418 181319 133474 181328
rect 133328 164756 133380 164762
rect 133328 164698 133380 164704
rect 133524 142497 133552 201146
rect 133604 199844 133656 199850
rect 133604 199786 133656 199792
rect 133616 163577 133644 199786
rect 133602 163568 133658 163577
rect 133602 163503 133658 163512
rect 133602 160440 133658 160449
rect 133602 160375 133658 160384
rect 133510 142488 133566 142497
rect 133510 142423 133566 142432
rect 133234 129840 133290 129849
rect 133234 129775 133290 129784
rect 132960 117292 133012 117298
rect 132960 117234 133012 117240
rect 133052 115932 133104 115938
rect 133052 115874 133104 115880
rect 133064 106457 133092 115874
rect 133050 106448 133106 106457
rect 133050 106383 133106 106392
rect 133510 106312 133566 106321
rect 133432 106270 133510 106298
rect 133432 104854 133460 106270
rect 133510 106247 133566 106256
rect 133420 104848 133472 104854
rect 133420 104790 133472 104796
rect 133144 95260 133196 95266
rect 133144 95202 133196 95208
rect 133156 91746 133184 95202
rect 133156 91718 133276 91746
rect 133248 70258 133276 91718
rect 133156 70230 133276 70258
rect 133156 60738 133184 70230
rect 133156 60710 133276 60738
rect 133248 57934 133276 60710
rect 133236 57928 133288 57934
rect 133236 57870 133288 57876
rect 133144 48340 133196 48346
rect 133144 48282 133196 48288
rect 133156 41426 133184 48282
rect 133156 41398 133276 41426
rect 133616 41410 133644 160375
rect 133708 141409 133736 700742
rect 133694 141400 133750 141409
rect 133694 141335 133750 141344
rect 133800 140457 133828 700878
rect 133892 180441 133920 700946
rect 137848 699718 137876 703520
rect 154132 703474 154160 703520
rect 154132 703446 154252 703474
rect 137836 699712 137888 699718
rect 137836 699654 137888 699660
rect 154224 698290 154252 703446
rect 170324 700670 170352 703520
rect 170312 700664 170364 700670
rect 170312 700606 170364 700612
rect 202800 700262 202828 703520
rect 218992 700806 219020 703520
rect 235184 700806 235212 703520
rect 267660 701010 267688 703520
rect 267648 701004 267700 701010
rect 267648 700946 267700 700952
rect 283852 700942 283880 703520
rect 300136 700942 300164 703520
rect 283840 700936 283892 700942
rect 283840 700878 283892 700884
rect 300124 700936 300176 700942
rect 300124 700878 300176 700884
rect 332520 700874 332548 703520
rect 332508 700868 332560 700874
rect 332508 700810 332560 700816
rect 218980 700800 219032 700806
rect 218980 700742 219032 700748
rect 235172 700800 235224 700806
rect 235172 700742 235224 700748
rect 348804 700738 348832 703520
rect 364996 700738 365024 703520
rect 348792 700732 348844 700738
rect 348792 700674 348844 700680
rect 364984 700732 365036 700738
rect 364984 700674 365036 700680
rect 397472 700602 397500 703520
rect 397460 700596 397512 700602
rect 397460 700538 397512 700544
rect 413664 700534 413692 703520
rect 413652 700528 413704 700534
rect 413652 700470 413704 700476
rect 202788 700256 202840 700262
rect 202788 700198 202840 700204
rect 429856 699718 429884 703520
rect 434076 700936 434128 700942
rect 434076 700878 434128 700884
rect 433984 700732 434036 700738
rect 433984 700674 434036 700680
rect 429844 699712 429896 699718
rect 429844 699654 429896 699660
rect 433892 699712 433944 699718
rect 433892 699654 433944 699660
rect 153568 698284 153620 698290
rect 153568 698226 153620 698232
rect 154212 698284 154264 698290
rect 154212 698226 154264 698232
rect 147588 697128 147640 697134
rect 147586 697096 147588 697105
rect 147640 697096 147642 697105
rect 147586 697031 147642 697040
rect 153580 688786 153608 698226
rect 154486 697232 154542 697241
rect 154486 697167 154542 697176
rect 173806 697232 173862 697241
rect 173806 697167 173862 697176
rect 193126 697232 193182 697241
rect 193126 697167 193182 697176
rect 212446 697232 212502 697241
rect 212446 697167 212502 697176
rect 231766 697232 231822 697241
rect 231766 697167 231822 697176
rect 251086 697232 251142 697241
rect 251086 697167 251142 697176
rect 270406 697232 270462 697241
rect 270406 697167 270462 697176
rect 289726 697232 289782 697241
rect 289726 697167 289782 697176
rect 309046 697232 309102 697241
rect 309046 697167 309102 697176
rect 328366 697232 328422 697241
rect 328366 697167 328422 697176
rect 154500 697134 154528 697167
rect 173820 697134 173848 697167
rect 193140 697134 193168 697167
rect 212460 697134 212488 697167
rect 231780 697134 231808 697167
rect 251100 697134 251128 697167
rect 270420 697134 270448 697167
rect 289740 697134 289768 697167
rect 309060 697134 309088 697167
rect 328380 697134 328408 697167
rect 154488 697128 154540 697134
rect 166908 697128 166960 697134
rect 154488 697070 154540 697076
rect 166906 697096 166908 697105
rect 173808 697128 173860 697134
rect 166960 697096 166962 697105
rect 186228 697128 186280 697134
rect 173808 697070 173860 697076
rect 186226 697096 186228 697105
rect 193128 697128 193180 697134
rect 186280 697096 186282 697105
rect 166906 697031 166962 697040
rect 205548 697128 205600 697134
rect 193128 697070 193180 697076
rect 205546 697096 205548 697105
rect 212448 697128 212500 697134
rect 205600 697096 205602 697105
rect 186226 697031 186282 697040
rect 224868 697128 224920 697134
rect 212448 697070 212500 697076
rect 224866 697096 224868 697105
rect 231768 697128 231820 697134
rect 224920 697096 224922 697105
rect 205546 697031 205602 697040
rect 244188 697128 244240 697134
rect 231768 697070 231820 697076
rect 244186 697096 244188 697105
rect 251088 697128 251140 697134
rect 244240 697096 244242 697105
rect 224866 697031 224922 697040
rect 263508 697128 263560 697134
rect 251088 697070 251140 697076
rect 263506 697096 263508 697105
rect 270408 697128 270460 697134
rect 263560 697096 263562 697105
rect 244186 697031 244242 697040
rect 282828 697128 282880 697134
rect 270408 697070 270460 697076
rect 282826 697096 282828 697105
rect 289728 697128 289780 697134
rect 282880 697096 282882 697105
rect 263506 697031 263562 697040
rect 302148 697128 302200 697134
rect 289728 697070 289780 697076
rect 302146 697096 302148 697105
rect 309048 697128 309100 697134
rect 302200 697096 302202 697105
rect 282826 697031 282882 697040
rect 321468 697128 321520 697134
rect 309048 697070 309100 697076
rect 321466 697096 321468 697105
rect 328368 697128 328420 697134
rect 321520 697096 321522 697105
rect 302146 697031 302202 697040
rect 328368 697070 328420 697076
rect 321466 697031 321522 697040
rect 153580 688758 153700 688786
rect 147770 686352 147826 686361
rect 147600 686310 147770 686338
rect 135258 686216 135314 686225
rect 135258 686151 135260 686160
rect 135312 686151 135314 686160
rect 142896 686180 142948 686186
rect 135260 686122 135312 686128
rect 142896 686122 142948 686128
rect 142908 685953 142936 686122
rect 147600 686089 147628 686310
rect 147770 686287 147826 686296
rect 147586 686080 147642 686089
rect 147586 686015 147642 686024
rect 153672 685982 153700 688758
rect 169022 686488 169078 686497
rect 169022 686423 169078 686432
rect 154578 686352 154634 686361
rect 154578 686287 154580 686296
rect 154632 686287 154634 686296
rect 159456 686316 159508 686322
rect 154580 686258 154632 686264
rect 159456 686258 159508 686264
rect 159468 686225 159496 686258
rect 169036 686225 169064 686423
rect 159454 686216 159510 686225
rect 159454 686151 159510 686160
rect 169022 686216 169078 686225
rect 169022 686151 169078 686160
rect 153292 685976 153344 685982
rect 142894 685944 142950 685953
rect 153292 685918 153344 685924
rect 153660 685976 153712 685982
rect 153660 685918 153712 685924
rect 142894 685879 142950 685888
rect 153304 684486 153332 685918
rect 153292 684480 153344 684486
rect 153292 684422 153344 684428
rect 153660 666596 153712 666602
rect 153660 666538 153712 666544
rect 153672 659682 153700 666538
rect 153488 659654 153700 659682
rect 153488 656878 153516 659654
rect 153476 656872 153528 656878
rect 153476 656814 153528 656820
rect 169022 650584 169078 650593
rect 169022 650519 169078 650528
rect 147770 650448 147826 650457
rect 147600 650406 147770 650434
rect 135258 650312 135314 650321
rect 135258 650247 135260 650256
rect 135312 650247 135314 650256
rect 142896 650276 142948 650282
rect 135260 650218 135312 650224
rect 142896 650218 142948 650224
rect 142908 650049 142936 650218
rect 147600 650185 147628 650406
rect 147770 650383 147826 650392
rect 154578 650448 154634 650457
rect 154578 650383 154580 650392
rect 154632 650383 154634 650392
rect 159456 650412 159508 650418
rect 154580 650354 154632 650360
rect 159456 650354 159508 650360
rect 159468 650321 159496 650354
rect 169036 650321 169064 650519
rect 159454 650312 159510 650321
rect 159454 650247 159510 650256
rect 169022 650312 169078 650321
rect 169022 650247 169078 650256
rect 147586 650176 147642 650185
rect 147586 650111 147642 650120
rect 142894 650040 142950 650049
rect 142894 649975 142950 649984
rect 153568 647284 153620 647290
rect 153568 647226 153620 647232
rect 153580 645862 153608 647226
rect 153568 645856 153620 645862
rect 153568 645798 153620 645804
rect 157062 639296 157118 639305
rect 157246 639296 157302 639305
rect 157118 639254 157246 639282
rect 157062 639231 157118 639240
rect 157246 639231 157302 639240
rect 171046 639296 171102 639305
rect 171046 639231 171102 639240
rect 171060 638897 171088 639231
rect 171046 638888 171102 638897
rect 171046 638823 171102 638832
rect 153292 636268 153344 636274
rect 153292 636210 153344 636216
rect 153304 630562 153332 636210
rect 153292 630556 153344 630562
rect 153292 630498 153344 630504
rect 153568 630556 153620 630562
rect 153568 630498 153620 630504
rect 153580 621110 153608 630498
rect 153568 621104 153620 621110
rect 153568 621046 153620 621052
rect 153476 620968 153528 620974
rect 153476 620910 153528 620916
rect 153488 611266 153516 620910
rect 153396 611238 153516 611266
rect 153396 601746 153424 611238
rect 157062 603392 157118 603401
rect 157246 603392 157302 603401
rect 157118 603350 157246 603378
rect 157062 603327 157118 603336
rect 157246 603327 157302 603336
rect 171046 603392 171102 603401
rect 171046 603327 171102 603336
rect 171060 602993 171088 603327
rect 171046 602984 171102 602993
rect 171046 602919 171102 602928
rect 153304 601718 153424 601746
rect 153304 598942 153332 601718
rect 153292 598936 153344 598942
rect 153292 598878 153344 598884
rect 169022 592648 169078 592657
rect 169022 592583 169078 592592
rect 147770 592512 147826 592521
rect 147600 592470 147770 592498
rect 135258 592376 135314 592385
rect 135258 592311 135260 592320
rect 135312 592311 135314 592320
rect 142896 592340 142948 592346
rect 135260 592282 135312 592288
rect 142896 592282 142948 592288
rect 142908 592113 142936 592282
rect 147600 592249 147628 592470
rect 147770 592447 147826 592456
rect 154578 592512 154634 592521
rect 154578 592447 154580 592456
rect 154632 592447 154634 592456
rect 159456 592476 159508 592482
rect 154580 592418 154632 592424
rect 159456 592418 159508 592424
rect 159468 592385 159496 592418
rect 169036 592385 169064 592583
rect 159454 592376 159510 592385
rect 159454 592311 159510 592320
rect 169022 592376 169078 592385
rect 169022 592311 169078 592320
rect 147586 592240 147642 592249
rect 147586 592175 147642 592184
rect 142894 592104 142950 592113
rect 142894 592039 142950 592048
rect 153476 589348 153528 589354
rect 153476 589290 153528 589296
rect 153488 579698 153516 589290
rect 270408 583704 270460 583710
rect 270408 583646 270460 583652
rect 307024 583704 307076 583710
rect 307024 583646 307076 583652
rect 191102 582992 191158 583001
rect 191102 582927 191158 582936
rect 153384 579692 153436 579698
rect 153384 579634 153436 579640
rect 153476 579692 153528 579698
rect 153476 579634 153528 579640
rect 153396 560318 153424 579634
rect 153292 560312 153344 560318
rect 153292 560254 153344 560260
rect 153384 560312 153436 560318
rect 153384 560254 153436 560260
rect 140044 553648 140096 553654
rect 140044 553590 140096 553596
rect 134156 398132 134208 398138
rect 134156 398074 134208 398080
rect 134168 397662 134196 398074
rect 134156 397656 134208 397662
rect 134156 397598 134208 397604
rect 134168 396030 134196 397598
rect 134156 396024 134208 396030
rect 134156 395966 134208 395972
rect 133972 386436 134024 386442
rect 133972 386378 134024 386384
rect 133984 386306 134012 386378
rect 133972 386300 134024 386306
rect 133972 386242 134024 386248
rect 134156 376780 134208 376786
rect 134156 376722 134208 376728
rect 134168 369866 134196 376722
rect 133984 369838 134196 369866
rect 133984 362250 134012 369838
rect 133984 362222 134288 362250
rect 134260 357406 134288 362222
rect 134248 357400 134300 357406
rect 134248 357342 134300 357348
rect 134248 347812 134300 347818
rect 134248 347754 134300 347760
rect 133970 341456 134026 341465
rect 133970 341391 134026 341400
rect 133878 180432 133934 180441
rect 133984 180402 134012 341391
rect 134260 331158 134288 347754
rect 134248 331152 134300 331158
rect 134248 331094 134300 331100
rect 134248 331016 134300 331022
rect 134248 330958 134300 330964
rect 134260 318782 134288 330958
rect 134248 318776 134300 318782
rect 134248 318718 134300 318724
rect 134156 309188 134208 309194
rect 134156 309130 134208 309136
rect 134168 302190 134196 309130
rect 134156 302184 134208 302190
rect 134156 302126 134208 302132
rect 134340 302184 134392 302190
rect 134340 302126 134392 302132
rect 134352 298110 134380 302126
rect 134340 298104 134392 298110
rect 134340 298046 134392 298052
rect 134248 288448 134300 288454
rect 134248 288390 134300 288396
rect 134260 278866 134288 288390
rect 134156 278860 134208 278866
rect 134156 278802 134208 278808
rect 134248 278860 134300 278866
rect 134248 278802 134300 278808
rect 134168 278746 134196 278802
rect 134168 278730 134288 278746
rect 134168 278724 134300 278730
rect 134168 278718 134248 278724
rect 134248 278666 134300 278672
rect 134248 269136 134300 269142
rect 134248 269078 134300 269084
rect 134260 265690 134288 269078
rect 134260 265662 134380 265690
rect 134352 260846 134380 265662
rect 134340 260840 134392 260846
rect 134340 260782 134392 260788
rect 134248 250640 134300 250646
rect 134248 250582 134300 250588
rect 134260 249801 134288 250582
rect 134062 249792 134118 249801
rect 134062 249727 134118 249736
rect 134246 249792 134302 249801
rect 134246 249727 134302 249736
rect 134076 240174 134104 249727
rect 134064 240168 134116 240174
rect 134064 240110 134116 240116
rect 134340 240168 134392 240174
rect 134340 240110 134392 240116
rect 134352 235346 134380 240110
rect 134340 235340 134392 235346
rect 134340 235282 134392 235288
rect 134248 222216 134300 222222
rect 134248 222158 134300 222164
rect 134260 215370 134288 222158
rect 134168 215342 134288 215370
rect 134168 205714 134196 215342
rect 134168 205686 134288 205714
rect 134156 201612 134208 201618
rect 134156 201554 134208 201560
rect 134168 200002 134196 201554
rect 134260 200122 134288 205686
rect 140056 202366 140084 553590
rect 146944 553580 146996 553586
rect 146944 553522 146996 553528
rect 144184 536852 144236 536858
rect 144184 536794 144236 536800
rect 140044 202360 140096 202366
rect 140044 202302 140096 202308
rect 142528 202224 142580 202230
rect 142528 202166 142580 202172
rect 134708 202156 134760 202162
rect 134708 202098 134760 202104
rect 134340 201544 134392 201550
rect 134340 201486 134392 201492
rect 134248 200116 134300 200122
rect 134248 200058 134300 200064
rect 134352 200002 134380 201486
rect 134720 200002 134748 202098
rect 142540 200002 142568 202166
rect 144196 202162 144224 536794
rect 146956 202230 146984 553522
rect 153304 553330 153332 560254
rect 160744 553920 160796 553926
rect 160744 553862 160796 553868
rect 153844 553512 153896 553518
rect 153844 553454 153896 553460
rect 153304 553302 153424 553330
rect 153396 543810 153424 553302
rect 153396 543782 153516 543810
rect 152464 542428 152516 542434
rect 152464 542370 152516 542376
rect 151084 518356 151136 518362
rect 151084 518298 151136 518304
rect 151096 202298 151124 518298
rect 152476 497894 152504 542370
rect 153488 531350 153516 543782
rect 153384 531344 153436 531350
rect 153384 531286 153436 531292
rect 153476 531344 153528 531350
rect 153476 531286 153528 531292
rect 153396 524482 153424 531286
rect 153384 524476 153436 524482
rect 153384 524418 153436 524424
rect 153476 524408 153528 524414
rect 153476 524350 153528 524356
rect 153488 521665 153516 524350
rect 153290 521656 153346 521665
rect 153290 521591 153346 521600
rect 153474 521656 153530 521665
rect 153474 521591 153530 521600
rect 153304 512038 153332 521591
rect 153292 512032 153344 512038
rect 153292 511974 153344 511980
rect 153568 512032 153620 512038
rect 153568 511974 153620 511980
rect 153580 505238 153608 511974
rect 153568 505232 153620 505238
rect 153568 505174 153620 505180
rect 153384 505096 153436 505102
rect 153384 505038 153436 505044
rect 152464 497888 152516 497894
rect 152464 497830 152516 497836
rect 153108 497888 153160 497894
rect 153108 497830 153160 497836
rect 153120 406502 153148 497830
rect 153396 495446 153424 505038
rect 153384 495440 153436 495446
rect 153384 495382 153436 495388
rect 153568 495440 153620 495446
rect 153568 495382 153620 495388
rect 153580 492658 153608 495382
rect 153292 492652 153344 492658
rect 153292 492594 153344 492600
rect 153568 492652 153620 492658
rect 153568 492594 153620 492600
rect 153304 483041 153332 492594
rect 153290 483032 153346 483041
rect 153290 482967 153346 482976
rect 153474 483032 153530 483041
rect 153474 482967 153530 482976
rect 153488 476134 153516 482967
rect 153292 476128 153344 476134
rect 153476 476128 153528 476134
rect 153344 476076 153424 476082
rect 153292 476070 153424 476076
rect 153476 476070 153528 476076
rect 153304 476054 153424 476070
rect 153396 473346 153424 476054
rect 153384 473340 153436 473346
rect 153384 473282 153436 473288
rect 153384 466404 153436 466410
rect 153384 466346 153436 466352
rect 153396 463706 153424 466346
rect 153396 463678 153516 463706
rect 153488 456770 153516 463678
rect 153396 456742 153516 456770
rect 153396 447273 153424 456742
rect 153382 447264 153438 447273
rect 153382 447199 153438 447208
rect 153382 444408 153438 444417
rect 153382 444343 153384 444352
rect 153436 444343 153438 444352
rect 153384 444314 153436 444320
rect 153384 437436 153436 437442
rect 153384 437378 153436 437384
rect 153396 434738 153424 437378
rect 153396 434710 153516 434738
rect 153488 425241 153516 434710
rect 153474 425232 153530 425241
rect 153474 425167 153530 425176
rect 153198 425096 153254 425105
rect 153254 425054 153332 425082
rect 153198 425031 153254 425040
rect 153304 418266 153332 425054
rect 153292 418260 153344 418266
rect 153292 418202 153344 418208
rect 153200 418124 153252 418130
rect 153200 418066 153252 418072
rect 153212 415410 153240 418066
rect 153200 415404 153252 415410
rect 153200 415346 153252 415352
rect 153476 415404 153528 415410
rect 153476 415346 153528 415352
rect 153488 408354 153516 415346
rect 153396 408326 153516 408354
rect 153108 406496 153160 406502
rect 153108 406438 153160 406444
rect 153120 406026 153148 406438
rect 152464 406020 152516 406026
rect 152464 405962 152516 405968
rect 153108 406020 153160 406026
rect 153108 405962 153160 405968
rect 152476 398206 152504 405962
rect 153396 398954 153424 408326
rect 153384 398948 153436 398954
rect 153384 398890 153436 398896
rect 152464 398200 152516 398206
rect 152464 398142 152516 398148
rect 153384 396092 153436 396098
rect 153384 396034 153436 396040
rect 153396 395962 153424 396034
rect 153384 395956 153436 395962
rect 153384 395898 153436 395904
rect 153292 389156 153344 389162
rect 153292 389098 153344 389104
rect 153304 379506 153332 389098
rect 153292 379500 153344 379506
rect 153292 379442 153344 379448
rect 153476 379500 153528 379506
rect 153476 379442 153528 379448
rect 153488 371906 153516 379442
rect 153488 371878 153608 371906
rect 153580 367062 153608 371878
rect 153568 367056 153620 367062
rect 153568 366998 153620 367004
rect 153660 357468 153712 357474
rect 153660 357410 153712 357416
rect 153672 350690 153700 357410
rect 153580 350662 153700 350690
rect 153580 347818 153608 350662
rect 153476 347812 153528 347818
rect 153476 347754 153528 347760
rect 153568 347812 153620 347818
rect 153568 347754 153620 347760
rect 153488 347698 153516 347754
rect 153488 347670 153608 347698
rect 153580 338162 153608 347670
rect 153384 338156 153436 338162
rect 153384 338098 153436 338104
rect 153568 338156 153620 338162
rect 153568 338098 153620 338104
rect 153396 331242 153424 338098
rect 153396 331214 153516 331242
rect 153488 318850 153516 331214
rect 153384 318844 153436 318850
rect 153384 318786 153436 318792
rect 153476 318844 153528 318850
rect 153476 318786 153528 318792
rect 153396 311982 153424 318786
rect 153384 311976 153436 311982
rect 153384 311918 153436 311924
rect 153476 311976 153528 311982
rect 153476 311918 153528 311924
rect 153488 302258 153516 311918
rect 153292 302252 153344 302258
rect 153292 302194 153344 302200
rect 153476 302252 153528 302258
rect 153476 302194 153528 302200
rect 153304 302138 153332 302194
rect 153304 302110 153424 302138
rect 153396 292618 153424 302110
rect 153396 292590 153516 292618
rect 153488 282946 153516 292590
rect 153292 282940 153344 282946
rect 153292 282882 153344 282888
rect 153476 282940 153528 282946
rect 153476 282882 153528 282888
rect 153304 282826 153332 282882
rect 153304 282798 153424 282826
rect 153396 280158 153424 282798
rect 153384 280152 153436 280158
rect 153384 280094 153436 280100
rect 153568 273284 153620 273290
rect 153568 273226 153620 273232
rect 153580 270502 153608 273226
rect 153568 270496 153620 270502
rect 153568 270438 153620 270444
rect 153660 260908 153712 260914
rect 153660 260850 153712 260856
rect 153672 254046 153700 260850
rect 153660 254040 153712 254046
rect 153660 253982 153712 253988
rect 153568 253904 153620 253910
rect 153568 253846 153620 253852
rect 153580 244202 153608 253846
rect 153396 244174 153608 244202
rect 153396 241482 153424 244174
rect 153304 241454 153424 241482
rect 153304 234734 153332 241454
rect 153292 234728 153344 234734
rect 153292 234670 153344 234676
rect 153292 234592 153344 234598
rect 153292 234534 153344 234540
rect 153304 231826 153332 234534
rect 153212 231798 153332 231826
rect 153212 225010 153240 231798
rect 153200 225004 153252 225010
rect 153200 224946 153252 224952
rect 153200 222216 153252 222222
rect 153200 222158 153252 222164
rect 153212 215354 153240 222158
rect 153200 215348 153252 215354
rect 153200 215290 153252 215296
rect 153292 215212 153344 215218
rect 153292 215154 153344 215160
rect 153304 212498 153332 215154
rect 153292 212492 153344 212498
rect 153292 212434 153344 212440
rect 153384 202904 153436 202910
rect 153384 202846 153436 202852
rect 151084 202292 151136 202298
rect 151084 202234 151136 202240
rect 146944 202224 146996 202230
rect 146944 202166 146996 202172
rect 144184 202156 144236 202162
rect 144184 202098 144236 202104
rect 153396 201210 153424 202846
rect 153856 202434 153884 553454
rect 159364 532772 159416 532778
rect 159364 532714 159416 532720
rect 157984 518288 158036 518294
rect 157984 518230 158036 518236
rect 157996 202570 158024 518230
rect 157984 202564 158036 202570
rect 157984 202506 158036 202512
rect 159376 202502 159404 532714
rect 160756 202638 160784 553862
rect 188344 407856 188396 407862
rect 188344 407798 188396 407804
rect 168656 395616 168708 395622
rect 168656 395558 168708 395564
rect 160744 202632 160796 202638
rect 160744 202574 160796 202580
rect 159364 202496 159416 202502
rect 159364 202438 159416 202444
rect 153844 202428 153896 202434
rect 153844 202370 153896 202376
rect 168380 202360 168432 202366
rect 168380 202302 168432 202308
rect 153384 201204 153436 201210
rect 153384 201146 153436 201152
rect 168392 200002 168420 202302
rect 168668 200002 168696 395558
rect 179512 395548 179564 395554
rect 179512 395490 179564 395496
rect 169116 202632 169168 202638
rect 169116 202574 169168 202580
rect 169128 200002 169156 202574
rect 176936 202564 176988 202570
rect 176936 202506 176988 202512
rect 176948 200002 176976 202506
rect 178040 202496 178092 202502
rect 178040 202438 178092 202444
rect 178052 200002 178080 202438
rect 178684 202156 178736 202162
rect 178684 202098 178736 202104
rect 178696 200002 178724 202098
rect 179524 200002 179552 395490
rect 188356 356046 188384 407798
rect 191116 398138 191144 582927
rect 195888 562012 195940 562018
rect 195888 561954 195940 561960
rect 192484 506524 192536 506530
rect 192484 506466 192536 506472
rect 191104 398132 191156 398138
rect 191104 398074 191156 398080
rect 185584 356040 185636 356046
rect 185584 355982 185636 355988
rect 188344 356040 188396 356046
rect 188344 355982 188396 355988
rect 185596 341465 185624 355982
rect 192496 342922 192524 506466
rect 195612 409488 195664 409494
rect 195612 409430 195664 409436
rect 195520 409148 195572 409154
rect 195520 409090 195572 409096
rect 192484 342916 192536 342922
rect 192484 342858 192536 342864
rect 185582 341456 185638 341465
rect 185582 341391 185638 341400
rect 195532 205018 195560 409090
rect 195624 205154 195652 409430
rect 195796 409420 195848 409426
rect 195796 409362 195848 409368
rect 195704 409216 195756 409222
rect 195704 409158 195756 409164
rect 195612 205148 195664 205154
rect 195612 205090 195664 205096
rect 195520 205012 195572 205018
rect 195520 204954 195572 204960
rect 195716 204950 195744 409158
rect 195808 205086 195836 409362
rect 195900 205222 195928 561954
rect 197084 561944 197136 561950
rect 197084 561886 197136 561892
rect 208676 561944 208728 561950
rect 208676 561886 208728 561892
rect 217876 561944 217928 561950
rect 217876 561886 217928 561892
rect 196992 561808 197044 561814
rect 196992 561750 197044 561756
rect 196900 410168 196952 410174
rect 196900 410110 196952 410116
rect 196808 409556 196860 409562
rect 196808 409498 196860 409504
rect 196716 409352 196768 409358
rect 196716 409294 196768 409300
rect 196624 409284 196676 409290
rect 196624 409226 196676 409232
rect 196636 205290 196664 409226
rect 196728 205358 196756 409294
rect 196716 205352 196768 205358
rect 196716 205294 196768 205300
rect 196624 205284 196676 205290
rect 196624 205226 196676 205232
rect 195888 205216 195940 205222
rect 195888 205158 195940 205164
rect 195796 205080 195848 205086
rect 195796 205022 195848 205028
rect 195704 204944 195756 204950
rect 195704 204886 195756 204892
rect 182180 202428 182232 202434
rect 182180 202370 182232 202376
rect 181260 202292 181312 202298
rect 181260 202234 181312 202240
rect 180340 202224 180392 202230
rect 180340 202166 180392 202172
rect 180352 200002 180380 202166
rect 181272 200002 181300 202234
rect 182192 200002 182220 202370
rect 196820 201822 196848 409498
rect 196912 202774 196940 410110
rect 196900 202768 196952 202774
rect 196900 202710 196952 202716
rect 197004 202201 197032 561750
rect 197096 202881 197124 561886
rect 197268 561876 197320 561882
rect 197268 561818 197320 561824
rect 197176 561740 197228 561746
rect 197176 561682 197228 561688
rect 197082 202872 197138 202881
rect 197082 202807 197138 202816
rect 197188 202745 197216 561682
rect 197174 202736 197230 202745
rect 197174 202671 197230 202680
rect 197280 202473 197308 561818
rect 202420 561808 202472 561814
rect 202420 561750 202472 561756
rect 202432 559980 202460 561750
rect 205548 561740 205600 561746
rect 205548 561682 205600 561688
rect 205560 559980 205588 561682
rect 208688 559980 208716 561886
rect 214748 561876 214800 561882
rect 214748 561818 214800 561824
rect 211618 561776 211674 561785
rect 211618 561711 211674 561720
rect 211632 559980 211660 561711
rect 214760 559980 214788 561818
rect 217888 559980 217916 561886
rect 222198 556200 222254 556209
rect 222198 556135 222254 556144
rect 198646 534168 198702 534177
rect 198646 534103 198702 534112
rect 198554 524648 198610 524657
rect 198554 524583 198610 524592
rect 198188 521076 198240 521082
rect 198188 521018 198240 521024
rect 198096 518288 198148 518294
rect 198096 518230 198148 518236
rect 198004 407244 198056 407250
rect 198004 407186 198056 407192
rect 197728 406632 197780 406638
rect 197728 406574 197780 406580
rect 197740 365702 197768 406574
rect 198016 396778 198044 407186
rect 198004 396772 198056 396778
rect 198004 396714 198056 396720
rect 198002 378720 198058 378729
rect 198002 378655 198058 378664
rect 197910 374368 197966 374377
rect 197910 374303 197966 374312
rect 197818 370288 197874 370297
rect 197818 370223 197874 370232
rect 197728 365696 197780 365702
rect 197728 365638 197780 365644
rect 197726 361856 197782 361865
rect 197726 361791 197782 361800
rect 197542 357504 197598 357513
rect 197542 357439 197598 357448
rect 197450 353424 197506 353433
rect 197450 353359 197506 353368
rect 197358 349072 197414 349081
rect 197358 349007 197414 349016
rect 197372 202502 197400 349007
rect 197464 203726 197492 353359
rect 197452 203720 197504 203726
rect 197452 203662 197504 203668
rect 197556 202570 197584 357439
rect 197634 344992 197690 345001
rect 197634 344927 197690 344936
rect 197648 202638 197676 344927
rect 197740 203930 197768 361791
rect 197728 203924 197780 203930
rect 197728 203866 197780 203872
rect 197832 203658 197860 370223
rect 197820 203652 197872 203658
rect 197820 203594 197872 203600
rect 197636 202632 197688 202638
rect 197636 202574 197688 202580
rect 197544 202564 197596 202570
rect 197544 202506 197596 202512
rect 197360 202496 197412 202502
rect 197266 202464 197322 202473
rect 197360 202438 197412 202444
rect 197266 202399 197322 202408
rect 196990 202192 197046 202201
rect 197924 202162 197952 374303
rect 198016 203862 198044 378655
rect 198108 339046 198136 518230
rect 198096 339040 198148 339046
rect 198096 338982 198148 338988
rect 198200 338842 198228 521018
rect 198280 521008 198332 521014
rect 198280 520950 198332 520956
rect 198188 338836 198240 338842
rect 198188 338778 198240 338784
rect 198292 338774 198320 520950
rect 198462 399664 198518 399673
rect 198462 399599 198518 399608
rect 198370 387152 198426 387161
rect 198370 387087 198426 387096
rect 198280 338768 198332 338774
rect 198280 338710 198332 338716
rect 198004 203856 198056 203862
rect 198004 203798 198056 203804
rect 198384 203590 198412 387087
rect 198476 203794 198504 399599
rect 198464 203788 198516 203794
rect 198464 203730 198516 203736
rect 198372 203584 198424 203590
rect 198372 203526 198424 203532
rect 196990 202127 197046 202136
rect 197912 202156 197964 202162
rect 197912 202098 197964 202104
rect 196808 201816 196860 201822
rect 196808 201758 196860 201764
rect 198568 201550 198596 524583
rect 198660 201958 198688 534103
rect 198738 529272 198794 529281
rect 198738 529207 198794 529216
rect 198648 201952 198700 201958
rect 198648 201894 198700 201900
rect 198752 201890 198780 529207
rect 199384 521212 199436 521218
rect 199384 521154 199436 521160
rect 198830 403744 198886 403753
rect 198830 403679 198886 403688
rect 198844 202230 198872 403679
rect 198922 395312 198978 395321
rect 198922 395247 198978 395256
rect 198936 202298 198964 395247
rect 199014 391232 199070 391241
rect 199014 391167 199070 391176
rect 199028 203998 199056 391167
rect 199106 382800 199162 382809
rect 199106 382735 199162 382744
rect 199016 203992 199068 203998
rect 199016 203934 199068 203940
rect 199120 202366 199148 382735
rect 199198 365936 199254 365945
rect 199198 365871 199254 365880
rect 199212 202434 199240 365871
rect 199292 342916 199344 342922
rect 199292 342858 199344 342864
rect 199200 202428 199252 202434
rect 199200 202370 199252 202376
rect 199108 202360 199160 202366
rect 199108 202302 199160 202308
rect 198924 202292 198976 202298
rect 198924 202234 198976 202240
rect 198832 202224 198884 202230
rect 198832 202166 198884 202172
rect 198740 201884 198792 201890
rect 198740 201826 198792 201832
rect 199304 201754 199332 342858
rect 199396 338910 199424 521154
rect 199476 521144 199528 521150
rect 199476 521086 199528 521092
rect 199488 338978 199516 521086
rect 200224 520118 200606 520146
rect 202892 520118 203550 520146
rect 199752 410100 199804 410106
rect 199752 410042 199804 410048
rect 199568 409692 199620 409698
rect 199568 409634 199620 409640
rect 199476 338972 199528 338978
rect 199476 338914 199528 338920
rect 199384 338904 199436 338910
rect 199384 338846 199436 338852
rect 199292 201748 199344 201754
rect 199292 201690 199344 201696
rect 199580 201686 199608 409634
rect 199660 409624 199712 409630
rect 199660 409566 199712 409572
rect 199568 201680 199620 201686
rect 199568 201622 199620 201628
rect 199672 201618 199700 409566
rect 199764 202450 199792 410042
rect 199844 410032 199896 410038
rect 199844 409974 199896 409980
rect 199856 202586 199884 409974
rect 199936 409964 199988 409970
rect 199936 409906 199988 409912
rect 199948 202842 199976 409906
rect 200028 409896 200080 409902
rect 200028 409838 200080 409844
rect 199936 202836 199988 202842
rect 199936 202778 199988 202784
rect 200040 202706 200068 409838
rect 200224 342922 200252 520118
rect 200580 410168 200632 410174
rect 200580 410110 200632 410116
rect 200592 408748 200620 410110
rect 202892 409698 202920 520118
rect 206664 517546 206692 520132
rect 205640 517540 205692 517546
rect 205640 517482 205692 517488
rect 206652 517540 206704 517546
rect 206652 517482 206704 517488
rect 203338 410408 203394 410417
rect 203338 410343 203394 410352
rect 202880 409692 202932 409698
rect 202880 409634 202932 409640
rect 203352 408748 203380 410343
rect 205652 409630 205680 517482
rect 206284 410508 206336 410514
rect 206284 410450 206336 410456
rect 205640 409624 205692 409630
rect 205640 409566 205692 409572
rect 206296 408748 206324 410450
rect 209044 409896 209096 409902
rect 209044 409838 209096 409844
rect 209056 408748 209084 409838
rect 209792 409562 209820 520132
rect 212552 520118 212934 520146
rect 215312 520118 216062 520146
rect 211988 410576 212040 410582
rect 211988 410518 212040 410524
rect 209780 409556 209832 409562
rect 209780 409498 209832 409504
rect 212000 408748 212028 410518
rect 212552 409494 212580 520118
rect 214748 409964 214800 409970
rect 214748 409906 214800 409912
rect 212540 409488 212592 409494
rect 212540 409430 212592 409436
rect 214760 408748 214788 409906
rect 215312 409426 215340 520118
rect 218992 518294 219020 520132
rect 218980 518288 219032 518294
rect 218980 518230 219032 518236
rect 217692 410100 217744 410106
rect 217692 410042 217744 410048
rect 215300 409420 215352 409426
rect 215300 409362 215352 409368
rect 217704 408748 217732 410042
rect 220452 410032 220504 410038
rect 220452 409974 220504 409980
rect 220464 408748 220492 409974
rect 222212 409222 222240 556135
rect 222290 552120 222346 552129
rect 222290 552055 222346 552064
rect 222200 409216 222252 409222
rect 222200 409158 222252 409164
rect 222304 409154 222332 552055
rect 222566 546952 222622 546961
rect 222566 546887 222622 546896
rect 222474 542600 222530 542609
rect 222474 542535 222530 542544
rect 222382 538384 222438 538393
rect 222382 538319 222438 538328
rect 222396 521218 222424 538319
rect 222384 521212 222436 521218
rect 222384 521154 222436 521160
rect 222488 521014 222516 542535
rect 222580 521150 222608 546887
rect 222658 533352 222714 533361
rect 222658 533287 222714 533296
rect 222568 521144 222620 521150
rect 222568 521086 222620 521092
rect 222672 521082 222700 533287
rect 222750 529000 222806 529009
rect 222750 528935 222806 528944
rect 222660 521076 222712 521082
rect 222660 521018 222712 521024
rect 222476 521008 222528 521014
rect 222476 520950 222528 520956
rect 222764 409358 222792 528935
rect 222842 524512 222898 524521
rect 222842 524447 222898 524456
rect 222752 409352 222804 409358
rect 222752 409294 222804 409300
rect 222856 409290 222884 524447
rect 267280 451376 267332 451382
rect 267280 451318 267332 451324
rect 251732 410848 251784 410854
rect 251732 410790 251784 410796
rect 266360 410848 266412 410854
rect 266360 410790 266412 410796
rect 246028 410780 246080 410786
rect 246028 410722 246080 410728
rect 228916 410712 228968 410718
rect 228916 410654 228968 410660
rect 223396 410644 223448 410650
rect 223396 410586 223448 410592
rect 222844 409284 222896 409290
rect 222844 409226 222896 409232
rect 222292 409148 222344 409154
rect 222292 409090 222344 409096
rect 223408 408748 223436 410586
rect 226154 410136 226210 410145
rect 226154 410071 226210 410080
rect 226168 408748 226196 410071
rect 228928 408748 228956 410654
rect 243268 410372 243320 410378
rect 243268 410314 243320 410320
rect 240324 410304 240376 410310
rect 231858 410272 231914 410281
rect 240324 410246 240376 410252
rect 231858 410207 231914 410216
rect 237564 410236 237616 410242
rect 231872 408748 231900 410207
rect 237564 410178 237616 410184
rect 234620 410168 234672 410174
rect 234620 410110 234672 410116
rect 234632 408748 234660 410110
rect 237576 408748 237604 410178
rect 240336 408748 240364 410246
rect 243280 408748 243308 410314
rect 246040 408748 246068 410722
rect 248972 410440 249024 410446
rect 248972 410382 249024 410388
rect 248984 408748 249012 410382
rect 251744 408748 251772 410790
rect 257436 410100 257488 410106
rect 257436 410042 257488 410048
rect 254676 410032 254728 410038
rect 254676 409974 254728 409980
rect 254688 408748 254716 409974
rect 257448 408748 257476 410042
rect 263138 410000 263194 410009
rect 260380 409964 260432 409970
rect 263138 409935 263194 409944
rect 260380 409906 260432 409912
rect 260392 408748 260420 409906
rect 263152 408748 263180 409935
rect 265900 409896 265952 409902
rect 265900 409838 265952 409844
rect 265912 408748 265940 409838
rect 200212 342916 200264 342922
rect 200212 342858 200264 342864
rect 200592 337754 200620 340068
rect 203352 337822 203380 340068
rect 203340 337816 203392 337822
rect 203340 337758 203392 337764
rect 200580 337748 200632 337754
rect 200580 337690 200632 337696
rect 206112 337618 206140 340068
rect 209056 337890 209084 340068
rect 211830 340054 212488 340082
rect 209964 339040 210016 339046
rect 209964 338982 210016 338988
rect 209044 337884 209096 337890
rect 209044 337826 209096 337832
rect 206100 337612 206152 337618
rect 206100 337554 206152 337560
rect 209976 328506 210004 338982
rect 209780 328500 209832 328506
rect 209780 328442 209832 328448
rect 209964 328500 210016 328506
rect 209964 328442 210016 328448
rect 209792 318782 209820 328442
rect 209780 318776 209832 318782
rect 209780 318718 209832 318724
rect 209780 309188 209832 309194
rect 209780 309130 209832 309136
rect 209792 299470 209820 309130
rect 209780 299464 209832 299470
rect 209780 299406 209832 299412
rect 209780 289876 209832 289882
rect 209780 289818 209832 289824
rect 209792 280158 209820 289818
rect 209780 280152 209832 280158
rect 209780 280094 209832 280100
rect 209780 270564 209832 270570
rect 209780 270506 209832 270512
rect 209792 260846 209820 270506
rect 209780 260840 209832 260846
rect 209780 260782 209832 260788
rect 209780 251320 209832 251326
rect 209780 251262 209832 251268
rect 209792 241505 209820 251262
rect 209778 241496 209834 241505
rect 209778 241431 209834 241440
rect 209962 241496 210018 241505
rect 209962 241431 210018 241440
rect 209976 231878 210004 241431
rect 209780 231872 209832 231878
rect 209780 231814 209832 231820
rect 209964 231872 210016 231878
rect 209964 231814 210016 231820
rect 209792 222193 209820 231814
rect 209778 222184 209834 222193
rect 209778 222119 209834 222128
rect 209962 222184 210018 222193
rect 209962 222119 210018 222128
rect 209976 212566 210004 222119
rect 209780 212560 209832 212566
rect 209780 212502 209832 212508
rect 209964 212560 210016 212566
rect 209964 212502 210016 212508
rect 209792 202858 209820 212502
rect 209792 202830 209912 202858
rect 200028 202700 200080 202706
rect 200028 202642 200080 202648
rect 199856 202558 200068 202586
rect 199764 202422 199976 202450
rect 199948 202026 199976 202422
rect 200040 202094 200068 202558
rect 200028 202088 200080 202094
rect 200028 202030 200080 202036
rect 199936 202020 199988 202026
rect 199936 201962 199988 201968
rect 199660 201612 199712 201618
rect 199660 201554 199712 201560
rect 198556 201544 198608 201550
rect 198556 201486 198608 201492
rect 202880 201544 202932 201550
rect 202880 201486 202932 201492
rect 202892 200002 202920 201486
rect 209884 200258 209912 202830
rect 211712 201884 211764 201890
rect 211712 201826 211764 201832
rect 211158 201648 211214 201657
rect 211158 201583 211214 201592
rect 209872 200252 209924 200258
rect 209872 200194 209924 200200
rect 210286 200252 210338 200258
rect 210286 200194 210338 200200
rect 134168 199974 134228 200002
rect 134352 199974 134596 200002
rect 134720 199974 135056 200002
rect 142540 199974 142876 200002
rect 168392 199974 168544 200002
rect 168668 199974 169004 200002
rect 169128 199974 169372 200002
rect 176948 199974 177192 200002
rect 178052 199974 178112 200002
rect 178696 199974 178940 200002
rect 179524 199974 179860 200002
rect 180352 199974 180688 200002
rect 181272 199974 181608 200002
rect 182192 199974 182436 200002
rect 202860 199974 202920 200002
rect 210298 199988 210326 200194
rect 211172 200002 211200 201583
rect 211140 199974 211200 200002
rect 211724 200002 211752 201826
rect 212460 201550 212488 340054
rect 214104 338972 214156 338978
rect 214104 338914 214156 338920
rect 214116 338042 214144 338914
rect 214024 338014 214144 338042
rect 214024 331362 214052 338014
rect 214760 337686 214788 340068
rect 215300 338904 215352 338910
rect 215300 338846 215352 338852
rect 214748 337680 214800 337686
rect 214748 337622 214800 337628
rect 214012 331356 214064 331362
rect 214012 331298 214064 331304
rect 213920 328500 213972 328506
rect 213920 328442 213972 328448
rect 212538 201920 212594 201929
rect 212538 201855 212594 201864
rect 212448 201544 212500 201550
rect 212448 201486 212500 201492
rect 212552 200002 212580 201855
rect 213458 201784 213514 201793
rect 213458 201719 213514 201728
rect 213472 200002 213500 201719
rect 213932 200258 213960 328442
rect 213920 200252 213972 200258
rect 213920 200194 213972 200200
rect 214610 200252 214662 200258
rect 214610 200194 214662 200200
rect 211724 199974 211968 200002
rect 212552 199974 212888 200002
rect 213472 199974 213716 200002
rect 214622 199988 214650 200194
rect 215312 200002 215340 338846
rect 217520 337822 217548 340068
rect 220464 337958 220492 340068
rect 220820 338836 220872 338842
rect 220820 338778 220872 338784
rect 220452 337952 220504 337958
rect 220452 337894 220504 337900
rect 220084 337884 220136 337890
rect 220084 337826 220136 337832
rect 215944 337816 215996 337822
rect 215944 337758 215996 337764
rect 217508 337816 217560 337822
rect 217508 337758 217560 337764
rect 215956 201890 215984 337758
rect 218058 202056 218114 202065
rect 218058 201991 218114 202000
rect 216036 201952 216088 201958
rect 216036 201894 216088 201900
rect 215944 201884 215996 201890
rect 215944 201826 215996 201832
rect 216048 200002 216076 201894
rect 216864 201612 216916 201618
rect 216864 201554 216916 201560
rect 216876 200002 216904 201554
rect 218072 200002 218100 201991
rect 219532 201748 219584 201754
rect 219532 201690 219584 201696
rect 218612 201680 218664 201686
rect 218612 201622 218664 201628
rect 218624 200002 218652 201622
rect 219544 200002 219572 201690
rect 220096 201550 220124 337826
rect 220358 202872 220414 202881
rect 220358 202807 220414 202816
rect 220084 201544 220136 201550
rect 220084 201486 220136 201492
rect 220372 200002 220400 202807
rect 220832 201822 220860 338778
rect 222200 338768 222252 338774
rect 222200 338710 222252 338716
rect 220820 201816 220872 201822
rect 220820 201758 220872 201764
rect 221280 201816 221332 201822
rect 221280 201758 221332 201764
rect 221292 200002 221320 201758
rect 222212 200002 222240 338710
rect 223224 336870 223252 340068
rect 226168 337890 226196 340068
rect 226156 337884 226208 337890
rect 226156 337826 226208 337832
rect 228928 337346 228956 340068
rect 231872 338026 231900 340068
rect 231860 338020 231912 338026
rect 231860 337962 231912 337968
rect 228916 337340 228968 337346
rect 228916 337282 228968 337288
rect 232504 337340 232556 337346
rect 232504 337282 232556 337288
rect 223212 336864 223264 336870
rect 223212 336806 223264 336812
rect 229744 336864 229796 336870
rect 229744 336806 229796 336812
rect 226892 205352 226944 205358
rect 226892 205294 226944 205300
rect 223854 202736 223910 202745
rect 223854 202671 223910 202680
rect 223028 201748 223080 201754
rect 223028 201690 223080 201696
rect 223040 200002 223068 201690
rect 223868 200002 223896 202671
rect 225142 202600 225198 202609
rect 225142 202535 225198 202544
rect 225156 200002 225184 202535
rect 226338 202464 226394 202473
rect 226338 202399 226394 202408
rect 226352 200002 226380 202399
rect 215312 199974 215464 200002
rect 216048 199974 216384 200002
rect 216876 199974 217212 200002
rect 218072 199974 218132 200002
rect 218624 199974 218960 200002
rect 219544 199974 219880 200002
rect 220372 199974 220708 200002
rect 221292 199974 221536 200002
rect 222212 199974 222456 200002
rect 223040 199974 223284 200002
rect 223868 199974 224204 200002
rect 225156 199974 225492 200002
rect 226320 199974 226380 200002
rect 226904 200002 226932 205294
rect 227904 205284 227956 205290
rect 227904 205226 227956 205232
rect 227916 200002 227944 205226
rect 228640 205216 228692 205222
rect 228640 205158 228692 205164
rect 228652 200002 228680 205158
rect 229560 205148 229612 205154
rect 229560 205090 229612 205096
rect 229572 200002 229600 205090
rect 229756 201822 229784 336806
rect 230480 205080 230532 205086
rect 230480 205022 230532 205028
rect 229744 201816 229796 201822
rect 229744 201758 229796 201764
rect 230492 200002 230520 205022
rect 231216 205012 231268 205018
rect 231216 204954 231268 204960
rect 231228 200002 231256 204954
rect 232134 202328 232190 202337
rect 232134 202263 232190 202272
rect 232148 200002 232176 202263
rect 232516 202026 232544 337282
rect 234632 337142 234660 340068
rect 237288 338768 237340 338774
rect 237194 338736 237250 338745
rect 237288 338710 237340 338716
rect 237194 338671 237250 338680
rect 234620 337136 234672 337142
rect 234620 337078 234672 337084
rect 233240 204944 233292 204950
rect 233240 204886 233292 204892
rect 232504 202020 232556 202026
rect 232504 201962 232556 201968
rect 233252 200002 233280 204886
rect 233422 202192 233478 202201
rect 233422 202127 233478 202136
rect 233436 200002 233464 202127
rect 236644 202088 236696 202094
rect 236644 202030 236696 202036
rect 236656 200002 236684 202030
rect 236736 202020 236788 202026
rect 236736 201962 236788 201968
rect 226904 199974 227240 200002
rect 227916 199974 228068 200002
rect 228652 199974 228988 200002
rect 229572 199974 229816 200002
rect 230492 199974 230736 200002
rect 231228 199974 231564 200002
rect 232148 199974 232484 200002
rect 233252 199974 233312 200002
rect 233436 199974 233772 200002
rect 236348 199974 236684 200002
rect 236748 200002 236776 201962
rect 237208 200002 237236 338671
rect 237300 202094 237328 338710
rect 237576 337278 237604 340068
rect 240152 340054 240350 340082
rect 238116 337952 238168 337958
rect 238116 337894 238168 337900
rect 238024 337748 238076 337754
rect 238024 337690 238076 337696
rect 237564 337272 237616 337278
rect 237564 337214 237616 337220
rect 237748 337136 237800 337142
rect 237748 337078 237800 337084
rect 237288 202088 237340 202094
rect 237288 202030 237340 202036
rect 237380 201816 237432 201822
rect 237380 201758 237432 201764
rect 237392 200002 237420 201758
rect 237760 200002 237788 337078
rect 238036 201822 238064 337690
rect 238128 202026 238156 337894
rect 240048 337748 240100 337754
rect 240048 337690 240100 337696
rect 238760 203992 238812 203998
rect 238760 203934 238812 203940
rect 238116 202020 238168 202026
rect 238116 201962 238168 201968
rect 238024 201816 238076 201822
rect 238024 201758 238076 201764
rect 238208 201612 238260 201618
rect 238208 201554 238260 201560
rect 238220 200002 238248 201554
rect 236748 199974 236808 200002
rect 237208 199974 237268 200002
rect 237392 199974 237636 200002
rect 237760 199974 238096 200002
rect 238220 199974 238556 200002
rect 238772 199918 238800 203934
rect 239680 202836 239732 202842
rect 239680 202778 239732 202784
rect 239220 202768 239272 202774
rect 239220 202710 239272 202716
rect 239232 200002 239260 202710
rect 239692 200002 239720 202778
rect 240060 202774 240088 337690
rect 240152 202842 240180 340054
rect 241428 337816 241480 337822
rect 241428 337758 241480 337764
rect 241440 202842 241468 337758
rect 243096 337754 243124 340068
rect 244188 338836 244240 338842
rect 244188 338778 244240 338784
rect 243084 337748 243136 337754
rect 243084 337690 243136 337696
rect 243084 337272 243136 337278
rect 243084 337214 243136 337220
rect 240140 202836 240192 202842
rect 240140 202778 240192 202784
rect 240508 202836 240560 202842
rect 240508 202778 240560 202784
rect 241428 202836 241480 202842
rect 241428 202778 241480 202784
rect 240048 202768 240100 202774
rect 240048 202710 240100 202716
rect 240520 200002 240548 202778
rect 242072 202768 242124 202774
rect 242072 202710 242124 202716
rect 241520 202700 241572 202706
rect 241520 202642 241572 202648
rect 240968 202088 241020 202094
rect 240968 202030 241020 202036
rect 240980 200002 241008 202030
rect 241060 201680 241112 201686
rect 241060 201622 241112 201628
rect 238924 199974 239260 200002
rect 239384 199974 239720 200002
rect 240304 199974 240548 200002
rect 240672 199974 241008 200002
rect 241072 200002 241100 201622
rect 241532 200002 241560 202642
rect 242084 200002 242112 202710
rect 242164 201884 242216 201890
rect 242164 201826 242216 201832
rect 241072 199974 241132 200002
rect 241532 199974 241592 200002
rect 242052 199974 242112 200002
rect 242176 200002 242204 201826
rect 242992 201748 243044 201754
rect 242992 201690 243044 201696
rect 243004 200002 243032 201690
rect 242176 199974 242420 200002
rect 242880 199974 243032 200002
rect 243096 199918 243124 337214
rect 244096 336864 244148 336870
rect 244096 336806 244148 336812
rect 244004 209772 244056 209778
rect 244004 209714 244056 209720
rect 243176 201680 243228 201686
rect 243176 201622 243228 201628
rect 243188 200002 243216 201622
rect 244016 200002 244044 209714
rect 244108 201754 244136 336806
rect 244200 209778 244228 338778
rect 246040 337822 246068 340068
rect 248696 338020 248748 338026
rect 248696 337962 248748 337968
rect 248512 337884 248564 337890
rect 248512 337826 248564 337832
rect 246028 337816 246080 337822
rect 246028 337758 246080 337764
rect 247684 337748 247736 337754
rect 247684 337690 247736 337696
rect 244924 337340 244976 337346
rect 244924 337282 244976 337288
rect 244188 209772 244240 209778
rect 244188 209714 244240 209720
rect 244648 202632 244700 202638
rect 244648 202574 244700 202580
rect 244096 201748 244148 201754
rect 244096 201690 244148 201696
rect 244660 200002 244688 202574
rect 244740 202564 244792 202570
rect 244740 202506 244792 202512
rect 243188 199974 243340 200002
rect 243708 199974 244044 200002
rect 244628 199974 244688 200002
rect 244752 200002 244780 202506
rect 244936 201754 244964 337282
rect 247592 203992 247644 203998
rect 247592 203934 247644 203940
rect 245200 202700 245252 202706
rect 245200 202642 245252 202648
rect 244924 201748 244976 201754
rect 244924 201690 244976 201696
rect 245212 200002 245240 202642
rect 247500 202564 247552 202570
rect 247500 202506 247552 202512
rect 246028 201748 246080 201754
rect 246028 201690 246080 201696
rect 245660 201612 245712 201618
rect 245660 201554 245712 201560
rect 245672 200002 245700 201554
rect 246040 200002 246068 201690
rect 246488 201544 246540 201550
rect 246488 201486 246540 201492
rect 246500 200002 246528 201486
rect 247512 200002 247540 202506
rect 244752 199974 245088 200002
rect 245212 199974 245456 200002
rect 245672 199974 245916 200002
rect 246040 199974 246376 200002
rect 246500 199974 246836 200002
rect 247204 199974 247540 200002
rect 247604 200002 247632 203934
rect 247696 202774 247724 337690
rect 247684 202768 247736 202774
rect 247684 202710 247736 202716
rect 247776 201952 247828 201958
rect 247776 201894 247828 201900
rect 247788 200002 247816 201894
rect 248524 200002 248552 337826
rect 248708 202042 248736 337962
rect 248800 336870 248828 340068
rect 250996 337884 251048 337890
rect 250996 337826 251048 337832
rect 248788 336864 248840 336870
rect 248788 336806 248840 336812
rect 250536 204060 250588 204066
rect 250536 204002 250588 204008
rect 248708 202014 249288 202042
rect 248972 201884 249024 201890
rect 248972 201826 249024 201832
rect 248984 200002 249012 201826
rect 247604 199974 247664 200002
rect 247788 199974 248124 200002
rect 248492 199974 248552 200002
rect 248952 199974 249012 200002
rect 249260 200002 249288 202014
rect 250076 201748 250128 201754
rect 250076 201690 250128 201696
rect 250088 200002 250116 201690
rect 250548 200002 250576 204002
rect 250904 202700 250956 202706
rect 250904 202642 250956 202648
rect 250916 200002 250944 202642
rect 251008 201754 251036 337826
rect 251744 337142 251772 340068
rect 253664 338904 253716 338910
rect 253664 338846 253716 338852
rect 251732 337136 251784 337142
rect 251732 337078 251784 337084
rect 252468 337136 252520 337142
rect 252468 337078 252520 337084
rect 252480 203674 252508 337078
rect 253572 204128 253624 204134
rect 253572 204070 253624 204076
rect 252388 203646 252508 203674
rect 251824 202768 251876 202774
rect 251824 202710 251876 202716
rect 251456 201952 251508 201958
rect 251456 201894 251508 201900
rect 250996 201748 251048 201754
rect 250996 201690 251048 201696
rect 251468 200002 251496 201894
rect 251836 200002 251864 202710
rect 251916 202496 251968 202502
rect 251916 202438 251968 202444
rect 249260 199974 249412 200002
rect 249872 199974 250116 200002
rect 250240 199974 250576 200002
rect 250700 199974 250944 200002
rect 251160 199974 251496 200002
rect 251620 199974 251864 200002
rect 251928 200002 251956 202438
rect 252388 201686 252416 203646
rect 252468 202496 252520 202502
rect 252468 202438 252520 202444
rect 252376 201680 252428 201686
rect 252376 201622 252428 201628
rect 252480 200002 252508 202438
rect 253112 201748 253164 201754
rect 253112 201690 253164 201696
rect 253124 200002 253152 201690
rect 253584 200002 253612 204070
rect 251928 199974 251988 200002
rect 252448 199974 252508 200002
rect 252908 199974 253152 200002
rect 253276 199974 253612 200002
rect 253676 200002 253704 338846
rect 253756 337816 253808 337822
rect 253756 337758 253808 337764
rect 253768 201754 253796 337758
rect 254504 336870 254532 340068
rect 257448 337754 257476 340068
rect 257712 338972 257764 338978
rect 257712 338914 257764 338920
rect 257436 337748 257488 337754
rect 257436 337690 257488 337696
rect 255320 337612 255372 337618
rect 255320 337554 255372 337560
rect 254492 336864 254544 336870
rect 254492 336806 254544 336812
rect 255332 204354 255360 337554
rect 257724 336734 257752 338914
rect 260208 337890 260236 340068
rect 262128 338428 262180 338434
rect 262128 338370 262180 338376
rect 260196 337884 260248 337890
rect 260196 337826 260248 337832
rect 258724 337680 258776 337686
rect 258724 337622 258776 337628
rect 258264 336864 258316 336870
rect 258264 336806 258316 336812
rect 257712 336728 257764 336734
rect 257712 336670 257764 336676
rect 257804 336728 257856 336734
rect 257804 336670 257856 336676
rect 257816 335306 257844 336670
rect 257804 335300 257856 335306
rect 257804 335242 257856 335248
rect 257712 317484 257764 317490
rect 257712 317426 257764 317432
rect 257724 317393 257752 317426
rect 257710 317384 257766 317393
rect 257710 317319 257766 317328
rect 257802 311808 257858 311817
rect 257802 311743 257858 311752
rect 257816 307766 257844 311743
rect 257804 307760 257856 307766
rect 257804 307702 257856 307708
rect 257896 298172 257948 298178
rect 257896 298114 257948 298120
rect 257908 288454 257936 298114
rect 257804 288448 257856 288454
rect 257804 288390 257856 288396
rect 257896 288448 257948 288454
rect 257896 288390 257948 288396
rect 257816 288318 257844 288390
rect 257804 288312 257856 288318
rect 257804 288254 257856 288260
rect 257896 278792 257948 278798
rect 257896 278734 257948 278740
rect 257908 273306 257936 278734
rect 257816 273278 257936 273306
rect 257816 270502 257844 273278
rect 257804 270496 257856 270502
rect 257804 270438 257856 270444
rect 257804 263560 257856 263566
rect 257804 263502 257856 263508
rect 257816 260846 257844 263502
rect 257804 260840 257856 260846
rect 257804 260782 257856 260788
rect 257804 253836 257856 253842
rect 257804 253778 257856 253784
rect 257816 251190 257844 253778
rect 257804 251184 257856 251190
rect 257804 251126 257856 251132
rect 257712 241528 257764 241534
rect 257712 241470 257764 241476
rect 257724 234666 257752 241470
rect 257712 234660 257764 234666
rect 257712 234602 257764 234608
rect 257804 234524 257856 234530
rect 257804 234466 257856 234472
rect 257816 231826 257844 234466
rect 257724 231798 257844 231826
rect 257724 225010 257752 231798
rect 257712 225004 257764 225010
rect 257712 224946 257764 224952
rect 257712 222216 257764 222222
rect 257712 222158 257764 222164
rect 257724 215354 257752 222158
rect 257712 215348 257764 215354
rect 257712 215290 257764 215296
rect 257804 215212 257856 215218
rect 257804 215154 257856 215160
rect 257816 212514 257844 215154
rect 257724 212486 257844 212514
rect 257724 205698 257752 212486
rect 257712 205692 257764 205698
rect 257712 205634 257764 205640
rect 255332 204326 256188 204354
rect 255780 204196 255832 204202
rect 255780 204138 255832 204144
rect 254032 202428 254084 202434
rect 254032 202370 254084 202376
rect 253756 201748 253808 201754
rect 253756 201690 253808 201696
rect 254044 200002 254072 202370
rect 255228 201816 255280 201822
rect 255228 201758 255280 201764
rect 254860 201544 254912 201550
rect 254860 201486 254912 201492
rect 254872 200002 254900 201486
rect 255240 200002 255268 201758
rect 255792 200002 255820 204138
rect 255964 202428 256016 202434
rect 255964 202370 256016 202376
rect 255976 200002 256004 202370
rect 253676 199974 253736 200002
rect 254044 199974 254196 200002
rect 254656 199974 254900 200002
rect 255024 199974 255268 200002
rect 255484 199974 255820 200002
rect 255944 199974 256004 200002
rect 256160 200002 256188 204326
rect 257160 203924 257212 203930
rect 257160 203866 257212 203872
rect 257066 202192 257122 202201
rect 257066 202127 257122 202136
rect 257080 200002 257108 202127
rect 256160 199974 256404 200002
rect 256772 199974 257108 200002
rect 257172 200002 257200 203866
rect 257712 202904 257764 202910
rect 257712 202846 257764 202852
rect 257724 200274 257752 202846
rect 258276 202450 258304 336806
rect 258736 202774 258764 337622
rect 260380 203856 260432 203862
rect 260380 203798 260432 203804
rect 258724 202768 258776 202774
rect 258724 202710 258776 202716
rect 258276 202422 258764 202450
rect 258448 202360 258500 202366
rect 258448 202302 258500 202308
rect 258356 202020 258408 202026
rect 258356 201962 258408 201968
rect 257678 200246 257752 200274
rect 257172 199974 257232 200002
rect 257678 199988 257706 200246
rect 258368 200002 258396 201962
rect 258060 199974 258396 200002
rect 258460 200002 258488 202302
rect 258736 200002 258764 202422
rect 260196 202224 260248 202230
rect 260196 202166 260248 202172
rect 259460 201748 259512 201754
rect 259460 201690 259512 201696
rect 259472 200002 259500 201690
rect 260104 201544 260156 201550
rect 260104 201486 260156 201492
rect 260116 200002 260144 201486
rect 258460 199974 258520 200002
rect 258736 199974 258980 200002
rect 259440 199974 259500 200002
rect 259808 199974 260144 200002
rect 260208 200002 260236 202166
rect 260392 200002 260420 203798
rect 262140 202450 262168 338370
rect 263152 337822 263180 340068
rect 265926 340054 266308 340082
rect 263140 337816 263192 337822
rect 263140 337758 263192 337764
rect 262772 203788 262824 203794
rect 262772 203730 262824 203736
rect 261772 202422 262168 202450
rect 260840 201612 260892 201618
rect 260840 201554 260892 201560
rect 260852 200002 260880 201554
rect 261772 200002 261800 202422
rect 261944 202360 261996 202366
rect 261944 202302 261996 202308
rect 260208 199974 260268 200002
rect 260392 199974 260728 200002
rect 260852 199974 261188 200002
rect 261556 199974 261800 200002
rect 261956 200002 261984 202302
rect 262678 201648 262734 201657
rect 262678 201583 262734 201592
rect 262692 200002 262720 201583
rect 261956 199974 262016 200002
rect 262476 199974 262720 200002
rect 262784 200002 262812 203730
rect 262956 203720 263008 203726
rect 262956 203662 263008 203668
rect 262968 200002 262996 203662
rect 265256 203652 265308 203658
rect 265256 203594 265308 203600
rect 263876 202768 263928 202774
rect 263876 202710 263928 202716
rect 263600 201680 263652 201686
rect 263600 201622 263652 201628
rect 263612 200002 263640 201622
rect 263888 200002 263916 202710
rect 265164 202360 265216 202366
rect 265164 202302 265216 202308
rect 264888 201816 264940 201822
rect 264888 201758 264940 201764
rect 264900 200002 264928 201758
rect 265176 200002 265204 202302
rect 262784 199974 262844 200002
rect 262968 199974 263304 200002
rect 263612 199974 263764 200002
rect 263888 199974 264224 200002
rect 264592 199974 264928 200002
rect 265052 199974 265204 200002
rect 265268 200002 265296 203594
rect 266174 202872 266230 202881
rect 266174 202807 266230 202816
rect 266188 200002 266216 202807
rect 266280 201890 266308 340054
rect 266372 204950 266400 410790
rect 267004 410712 267056 410718
rect 267004 410654 267056 410660
rect 266728 410644 266780 410650
rect 266728 410586 266780 410592
rect 266452 410508 266504 410514
rect 266452 410450 266504 410456
rect 266360 204944 266412 204950
rect 266360 204886 266412 204892
rect 266360 202768 266412 202774
rect 266360 202710 266412 202716
rect 266268 201884 266320 201890
rect 266268 201826 266320 201832
rect 266372 200002 266400 202710
rect 265268 199974 265512 200002
rect 265972 199974 266216 200002
rect 266340 199974 266400 200002
rect 266464 200002 266492 410450
rect 266544 410372 266596 410378
rect 266544 410314 266596 410320
rect 266556 201958 266584 410314
rect 266636 410304 266688 410310
rect 266636 410246 266688 410252
rect 266544 201952 266596 201958
rect 266544 201894 266596 201900
rect 266648 201754 266676 410246
rect 266636 201748 266688 201754
rect 266636 201690 266688 201696
rect 266740 201618 266768 410586
rect 266820 410168 266872 410174
rect 266820 410110 266872 410116
rect 266832 202298 266860 410110
rect 266910 399664 266966 399673
rect 266910 399599 266966 399608
rect 266924 202366 266952 399599
rect 266912 202360 266964 202366
rect 266912 202302 266964 202308
rect 266820 202292 266872 202298
rect 266820 202234 266872 202240
rect 267016 201618 267044 410654
rect 267096 410576 267148 410582
rect 267096 410518 267148 410524
rect 267108 201754 267136 410518
rect 267186 357504 267242 357513
rect 267186 357439 267242 357448
rect 267200 202774 267228 357439
rect 267292 355366 267320 451318
rect 267832 410780 267884 410786
rect 267832 410722 267884 410728
rect 267740 410440 267792 410446
rect 267740 410382 267792 410388
rect 267372 410236 267424 410242
rect 267372 410178 267424 410184
rect 267280 355360 267332 355366
rect 267280 355302 267332 355308
rect 267278 353424 267334 353433
rect 267278 353359 267334 353368
rect 267188 202768 267240 202774
rect 267188 202710 267240 202716
rect 267292 202094 267320 353359
rect 267384 338774 267412 410178
rect 267464 410100 267516 410106
rect 267464 410042 267516 410048
rect 267476 338842 267504 410042
rect 267556 409964 267608 409970
rect 267556 409906 267608 409912
rect 267568 338978 267596 409906
rect 267646 349072 267702 349081
rect 267646 349007 267702 349016
rect 267556 338972 267608 338978
rect 267556 338914 267608 338920
rect 267464 338836 267516 338842
rect 267464 338778 267516 338784
rect 267372 338768 267424 338774
rect 267372 338710 267424 338716
rect 267464 204944 267516 204950
rect 267464 204886 267516 204892
rect 267372 203584 267424 203590
rect 267372 203526 267424 203532
rect 267280 202088 267332 202094
rect 267280 202030 267332 202036
rect 267096 201748 267148 201754
rect 267096 201690 267148 201696
rect 266728 201612 266780 201618
rect 266728 201554 266780 201560
rect 267004 201612 267056 201618
rect 267004 201554 267056 201560
rect 267384 200002 267412 203526
rect 266464 199974 266800 200002
rect 267260 199974 267412 200002
rect 267476 200002 267504 204886
rect 267660 201550 267688 349007
rect 267752 201822 267780 410382
rect 267844 202570 267872 410722
rect 268844 410032 268896 410038
rect 268844 409974 268896 409980
rect 267922 403744 267978 403753
rect 267922 403679 267978 403688
rect 267936 202842 267964 403679
rect 268014 395312 268070 395321
rect 268014 395247 268070 395256
rect 268028 204066 268056 395247
rect 268106 391232 268162 391241
rect 268106 391167 268162 391176
rect 268016 204060 268068 204066
rect 268016 204002 268068 204008
rect 267924 202836 267976 202842
rect 267924 202778 267976 202784
rect 268120 202638 268148 391167
rect 268198 386880 268254 386889
rect 268198 386815 268254 386824
rect 268212 203998 268240 386815
rect 268290 382800 268346 382809
rect 268290 382735 268346 382744
rect 268304 204202 268332 382735
rect 268382 378448 268438 378457
rect 268382 378383 268438 378392
rect 268292 204196 268344 204202
rect 268292 204138 268344 204144
rect 268200 203992 268252 203998
rect 268200 203934 268252 203940
rect 268396 202706 268424 378383
rect 268474 374368 268530 374377
rect 268474 374303 268530 374312
rect 268384 202700 268436 202706
rect 268384 202642 268436 202648
rect 268108 202632 268160 202638
rect 268108 202574 268160 202580
rect 267832 202564 267884 202570
rect 267832 202506 267884 202512
rect 268488 202502 268516 374303
rect 268566 370016 268622 370025
rect 268566 369951 268622 369960
rect 268476 202496 268528 202502
rect 268476 202438 268528 202444
rect 268580 202434 268608 369951
rect 268658 365936 268714 365945
rect 268658 365871 268714 365880
rect 268568 202428 268620 202434
rect 268568 202370 268620 202376
rect 268672 202026 268700 365871
rect 268750 361584 268806 361593
rect 268750 361519 268806 361528
rect 268660 202020 268712 202026
rect 268660 201962 268712 201968
rect 267740 201816 267792 201822
rect 267740 201758 267792 201764
rect 268200 201748 268252 201754
rect 268200 201690 268252 201696
rect 267740 201612 267792 201618
rect 267740 201554 267792 201560
rect 267648 201544 267700 201550
rect 267648 201486 267700 201492
rect 267752 200002 267780 201554
rect 268212 200002 268240 201690
rect 268764 200002 268792 361519
rect 268856 338910 268884 409974
rect 268936 409896 268988 409902
rect 268936 409838 268988 409844
rect 268844 338904 268896 338910
rect 268844 338846 268896 338852
rect 268948 338434 268976 409838
rect 269026 344992 269082 345001
rect 269026 344927 269082 344936
rect 268936 338428 268988 338434
rect 268936 338370 268988 338376
rect 269040 204134 269068 344927
rect 269028 204128 269080 204134
rect 269028 204070 269080 204076
rect 269488 202156 269540 202162
rect 269488 202098 269540 202104
rect 269120 201884 269172 201890
rect 269120 201826 269172 201832
rect 269132 200002 269160 201826
rect 269500 200002 269528 202098
rect 270420 200002 270448 583646
rect 287704 583636 287756 583642
rect 287704 583578 287756 583584
rect 281448 583024 281500 583030
rect 281448 582966 281500 582972
rect 274546 582856 274602 582865
rect 274546 582791 274602 582800
rect 272524 569968 272576 569974
rect 272524 569910 272576 569916
rect 271788 393984 271840 393990
rect 271788 393926 271840 393932
rect 271800 202842 271828 393926
rect 270960 202836 271012 202842
rect 270960 202778 271012 202784
rect 271788 202836 271840 202842
rect 271788 202778 271840 202784
rect 272248 202836 272300 202842
rect 272248 202778 272300 202784
rect 270972 200002 271000 202778
rect 271420 202768 271472 202774
rect 271420 202710 271472 202716
rect 271432 200002 271460 202710
rect 271696 202156 271748 202162
rect 271696 202098 271748 202104
rect 271708 200002 271736 202098
rect 272260 200002 272288 202778
rect 272536 202774 272564 569910
rect 273168 556232 273220 556238
rect 273168 556174 273220 556180
rect 273180 202842 273208 556174
rect 274560 202842 274588 582791
rect 280068 521688 280120 521694
rect 280068 521630 280120 521636
rect 279424 518968 279476 518974
rect 279424 518910 279476 518916
rect 277308 497140 277360 497146
rect 277308 497082 277360 497088
rect 277216 392624 277268 392630
rect 277216 392566 277268 392572
rect 273168 202836 273220 202842
rect 273168 202778 273220 202784
rect 273996 202836 274048 202842
rect 273996 202778 274048 202784
rect 274548 202836 274600 202842
rect 274548 202778 274600 202784
rect 277032 202836 277084 202842
rect 277032 202778 277084 202784
rect 272524 202768 272576 202774
rect 272524 202710 272576 202716
rect 273628 201680 273680 201686
rect 273628 201622 273680 201628
rect 273640 200002 273668 201622
rect 274008 200002 274036 202778
rect 275284 202428 275336 202434
rect 275284 202370 275336 202376
rect 275296 200002 275324 202370
rect 275744 202224 275796 202230
rect 275744 202166 275796 202172
rect 275756 200002 275784 202166
rect 277044 200002 277072 202778
rect 277228 200002 277256 392566
rect 277320 202842 277348 497082
rect 279436 202842 279464 518910
rect 279516 497004 279568 497010
rect 279516 496946 279568 496952
rect 277308 202836 277360 202842
rect 277308 202778 277360 202784
rect 278688 202836 278740 202842
rect 278688 202778 278740 202784
rect 279424 202836 279476 202842
rect 279424 202778 279476 202784
rect 278700 200002 278728 202778
rect 279240 202768 279292 202774
rect 279240 202710 279292 202716
rect 279252 200002 279280 202710
rect 279528 201686 279556 496946
rect 280080 202774 280108 521630
rect 281356 392692 281408 392698
rect 281356 392634 281408 392640
rect 281368 202842 281396 392634
rect 280528 202836 280580 202842
rect 280528 202778 280580 202784
rect 281356 202836 281408 202842
rect 281356 202778 281408 202784
rect 280068 202768 280120 202774
rect 280068 202710 280120 202716
rect 279516 201680 279568 201686
rect 279516 201622 279568 201628
rect 280540 200002 280568 202778
rect 281460 202366 281488 582966
rect 286968 538280 287020 538286
rect 286968 538222 287020 538228
rect 284944 516180 284996 516186
rect 284944 516122 284996 516128
rect 284300 497752 284352 497758
rect 284300 497694 284352 497700
rect 284208 497616 284260 497622
rect 284208 497558 284260 497564
rect 284022 491328 284078 491337
rect 284022 491263 284024 491272
rect 284076 491263 284078 491272
rect 284024 491234 284076 491240
rect 284116 485784 284168 485790
rect 284116 485726 284168 485732
rect 284128 481642 284156 485726
rect 284116 481636 284168 481642
rect 284116 481578 284168 481584
rect 284116 463820 284168 463826
rect 284116 463762 284168 463768
rect 284128 463690 284156 463762
rect 283840 463684 283892 463690
rect 283840 463626 283892 463632
rect 284116 463684 284168 463690
rect 284116 463626 284168 463632
rect 283852 454073 283880 463626
rect 283838 454064 283894 454073
rect 283838 453999 283894 454008
rect 284022 454064 284078 454073
rect 284022 453999 284024 454008
rect 284076 453999 284078 454008
rect 284024 453970 284076 453976
rect 284116 444508 284168 444514
rect 284116 444450 284168 444456
rect 284128 444378 284156 444450
rect 283840 444372 283892 444378
rect 283840 444314 283892 444320
rect 284116 444372 284168 444378
rect 284116 444314 284168 444320
rect 283852 434761 283880 444314
rect 283838 434752 283894 434761
rect 283838 434687 283894 434696
rect 284022 434752 284078 434761
rect 284022 434687 284024 434696
rect 284076 434687 284078 434696
rect 284024 434658 284076 434664
rect 284116 425196 284168 425202
rect 284116 425138 284168 425144
rect 284128 425066 284156 425138
rect 283840 425060 283892 425066
rect 283840 425002 283892 425008
rect 284116 425060 284168 425066
rect 284116 425002 284168 425008
rect 283852 415449 283880 425002
rect 283838 415440 283894 415449
rect 283838 415375 283894 415384
rect 284022 415440 284078 415449
rect 284022 415375 284024 415384
rect 284076 415375 284078 415384
rect 284024 415346 284076 415352
rect 284024 405748 284076 405754
rect 284024 405690 284076 405696
rect 284036 394874 284064 405690
rect 284024 394868 284076 394874
rect 284024 394810 284076 394816
rect 284024 394732 284076 394738
rect 284024 394674 284076 394680
rect 284036 393310 284064 394674
rect 284024 393304 284076 393310
rect 284024 393246 284076 393252
rect 284116 383716 284168 383722
rect 284116 383658 284168 383664
rect 284128 380225 284156 383658
rect 284114 380216 284170 380225
rect 284114 380151 284170 380160
rect 284114 367160 284170 367169
rect 284114 367095 284170 367104
rect 284128 367062 284156 367095
rect 284116 367056 284168 367062
rect 284116 366998 284168 367004
rect 284024 357468 284076 357474
rect 284024 357410 284076 357416
rect 284036 357354 284064 357410
rect 283944 357326 284064 357354
rect 283944 347993 283972 357326
rect 283930 347984 283986 347993
rect 283930 347919 283986 347928
rect 284114 347848 284170 347857
rect 284114 347783 284170 347792
rect 284128 347750 284156 347783
rect 284116 347744 284168 347750
rect 284116 347686 284168 347692
rect 284024 338224 284076 338230
rect 284024 338166 284076 338172
rect 284036 338094 284064 338166
rect 284024 338088 284076 338094
rect 284024 338030 284076 338036
rect 284116 328568 284168 328574
rect 284116 328510 284168 328516
rect 284128 328438 284156 328510
rect 284116 328432 284168 328438
rect 284116 328374 284168 328380
rect 284024 318844 284076 318850
rect 284024 318786 284076 318792
rect 284036 318730 284064 318786
rect 283944 318702 284064 318730
rect 283944 309262 283972 318702
rect 283932 309256 283984 309262
rect 283932 309198 283984 309204
rect 284116 309256 284168 309262
rect 284116 309198 284168 309204
rect 284128 309126 284156 309198
rect 284116 309120 284168 309126
rect 284116 309062 284168 309068
rect 284024 299600 284076 299606
rect 284024 299542 284076 299548
rect 284036 299470 284064 299542
rect 284024 299464 284076 299470
rect 284024 299406 284076 299412
rect 284116 289944 284168 289950
rect 284116 289886 284168 289892
rect 284128 289814 284156 289886
rect 284116 289808 284168 289814
rect 284116 289750 284168 289756
rect 284024 280288 284076 280294
rect 284024 280230 284076 280236
rect 284036 280158 284064 280230
rect 284024 280152 284076 280158
rect 284024 280094 284076 280100
rect 284024 270564 284076 270570
rect 284024 270506 284076 270512
rect 284036 263702 284064 270506
rect 284024 263696 284076 263702
rect 284024 263638 284076 263644
rect 284024 260976 284076 260982
rect 284024 260918 284076 260924
rect 284036 260846 284064 260918
rect 284024 260840 284076 260846
rect 284024 260782 284076 260788
rect 284116 254652 284168 254658
rect 284116 254594 284168 254600
rect 284128 241505 284156 254594
rect 284220 251462 284248 497558
rect 284312 491337 284340 497694
rect 284298 491328 284354 491337
rect 284298 491263 284354 491272
rect 284300 260840 284352 260846
rect 284300 260782 284352 260788
rect 284312 254658 284340 260782
rect 284300 254652 284352 254658
rect 284300 254594 284352 254600
rect 284208 251456 284260 251462
rect 284208 251398 284260 251404
rect 284208 251252 284260 251258
rect 284208 251194 284260 251200
rect 284114 241496 284170 241505
rect 284114 241431 284170 241440
rect 284116 231872 284168 231878
rect 284116 231814 284168 231820
rect 284128 224890 284156 231814
rect 284036 224862 284156 224890
rect 284036 222170 284064 224862
rect 283944 222142 284064 222170
rect 283944 215422 283972 222142
rect 283932 215416 283984 215422
rect 283932 215358 283984 215364
rect 283932 215280 283984 215286
rect 283932 215222 283984 215228
rect 283944 212537 283972 215222
rect 283654 212528 283710 212537
rect 283654 212463 283710 212472
rect 283930 212528 283986 212537
rect 283930 212463 283986 212472
rect 283668 202910 283696 212463
rect 283656 202904 283708 202910
rect 283656 202846 283708 202852
rect 283748 202904 283800 202910
rect 283748 202846 283800 202852
rect 282276 202768 282328 202774
rect 282276 202710 282328 202716
rect 280988 202360 281040 202366
rect 280988 202302 281040 202308
rect 281448 202360 281500 202366
rect 281448 202302 281500 202308
rect 281000 200002 281028 202302
rect 282288 200002 282316 202710
rect 282736 202360 282788 202366
rect 282736 202302 282788 202308
rect 282748 200002 282776 202302
rect 283564 202292 283616 202298
rect 283564 202234 283616 202240
rect 283576 200002 283604 202234
rect 283760 200274 283788 202846
rect 267476 199974 267628 200002
rect 267752 199974 268088 200002
rect 268212 199974 268548 200002
rect 268764 199974 269008 200002
rect 269132 199974 269376 200002
rect 269500 199974 269836 200002
rect 270296 199974 270448 200002
rect 270664 199974 271000 200002
rect 271124 199974 271460 200002
rect 271584 199974 271736 200002
rect 272044 199974 272288 200002
rect 273332 199974 273668 200002
rect 273792 199974 274036 200002
rect 275080 199974 275324 200002
rect 275448 199974 275784 200002
rect 276828 199974 277072 200002
rect 277196 199974 277256 200002
rect 278576 199974 278728 200002
rect 278944 199974 279280 200002
rect 280232 199974 280568 200002
rect 280692 199974 281028 200002
rect 281980 199974 282316 200002
rect 282440 199974 282776 200002
rect 283360 199974 283604 200002
rect 283714 200246 283788 200274
rect 283714 199988 283742 200246
rect 284220 200002 284248 251194
rect 284298 241496 284354 241505
rect 284298 241431 284354 241440
rect 284312 231878 284340 241431
rect 284300 231872 284352 231878
rect 284300 231814 284352 231820
rect 284956 202774 284984 516122
rect 285588 497412 285640 497418
rect 285588 497354 285640 497360
rect 285036 496868 285088 496874
rect 285036 496810 285088 496816
rect 284944 202768 284996 202774
rect 284944 202710 284996 202716
rect 285048 202434 285076 496810
rect 285036 202428 285088 202434
rect 285036 202370 285088 202376
rect 285600 200002 285628 497354
rect 286876 392828 286928 392834
rect 286876 392770 286928 392776
rect 286888 202502 286916 392770
rect 286232 202496 286284 202502
rect 286232 202438 286284 202444
rect 286876 202496 286928 202502
rect 286876 202438 286928 202444
rect 286244 200002 286272 202438
rect 286980 200002 287008 538222
rect 287520 202496 287572 202502
rect 287520 202438 287572 202444
rect 287532 200002 287560 202438
rect 287716 202230 287744 583578
rect 298468 583228 298520 583234
rect 298468 583170 298520 583176
rect 298376 583160 298428 583166
rect 298376 583102 298428 583108
rect 293868 583092 293920 583098
rect 293868 583034 293920 583040
rect 291108 582820 291160 582826
rect 291108 582762 291160 582768
rect 289728 497820 289780 497826
rect 289728 497762 289780 497768
rect 288348 497072 288400 497078
rect 288348 497014 288400 497020
rect 288256 392760 288308 392766
rect 288256 392702 288308 392708
rect 288268 202502 288296 392702
rect 288256 202496 288308 202502
rect 288256 202438 288308 202444
rect 287704 202224 287756 202230
rect 287704 202166 287756 202172
rect 288360 200138 288388 497014
rect 289740 202502 289768 497762
rect 291016 497684 291068 497690
rect 291016 497626 291068 497632
rect 291028 202502 291056 497626
rect 289452 202496 289504 202502
rect 289452 202438 289504 202444
rect 289728 202496 289780 202502
rect 289728 202438 289780 202444
rect 290556 202496 290608 202502
rect 290556 202438 290608 202444
rect 291016 202496 291068 202502
rect 291016 202438 291068 202444
rect 289268 202428 289320 202434
rect 289268 202370 289320 202376
rect 288808 202224 288860 202230
rect 288808 202166 288860 202172
rect 287992 200110 288388 200138
rect 287992 200002 288020 200110
rect 288820 200002 288848 202166
rect 289280 200002 289308 202370
rect 289464 200002 289492 202438
rect 290568 200002 290596 202438
rect 291120 200138 291148 582762
rect 292488 497344 292540 497350
rect 292488 497286 292540 497292
rect 292396 392964 292448 392970
rect 292396 392906 292448 392912
rect 292304 392896 292356 392902
rect 292304 392838 292356 392844
rect 292212 202496 292264 202502
rect 292212 202438 292264 202444
rect 291384 202020 291436 202026
rect 291384 201962 291436 201968
rect 291028 200110 291148 200138
rect 291028 200002 291056 200110
rect 291396 200002 291424 201962
rect 292224 200002 292252 202438
rect 284188 199974 284248 200002
rect 285476 199974 285628 200002
rect 285936 199974 286272 200002
rect 286764 199974 287008 200002
rect 287224 199974 287560 200002
rect 287684 199974 288020 200002
rect 288512 199974 288848 200002
rect 288972 199974 289308 200002
rect 289432 199974 289492 200002
rect 290260 199974 290596 200002
rect 290720 199974 291056 200002
rect 291180 199974 291424 200002
rect 292008 199974 292252 200002
rect 292316 200002 292344 392838
rect 292408 202502 292436 392906
rect 292396 202496 292448 202502
rect 292396 202438 292448 202444
rect 292500 202026 292528 497286
rect 292488 202020 292540 202026
rect 292488 201962 292540 201968
rect 293776 201612 293828 201618
rect 293776 201554 293828 201560
rect 293040 201544 293092 201550
rect 293040 201486 293092 201492
rect 293052 200002 293080 201486
rect 293788 200002 293816 201554
rect 293880 201550 293908 583034
rect 298284 582956 298336 582962
rect 298284 582898 298336 582904
rect 298192 582684 298244 582690
rect 298192 582626 298244 582632
rect 294604 582616 294656 582622
rect 294604 582558 294656 582564
rect 294616 202366 294644 582558
rect 298006 575784 298062 575793
rect 298006 575719 298062 575728
rect 298020 575550 298048 575719
rect 298008 575544 298060 575550
rect 298008 575486 298060 575492
rect 297454 572792 297510 572801
rect 297454 572727 297510 572736
rect 296626 565856 296682 565865
rect 296626 565791 296682 565800
rect 296076 534064 296128 534070
rect 296076 534006 296128 534012
rect 296088 521626 296116 534006
rect 296534 531448 296590 531457
rect 296534 531383 296590 531392
rect 295340 521620 295392 521626
rect 295340 521562 295392 521568
rect 296076 521620 296128 521626
rect 296076 521562 296128 521568
rect 295352 521286 295380 521562
rect 295340 521280 295392 521286
rect 295340 521222 295392 521228
rect 294696 509312 294748 509318
rect 294696 509254 294748 509260
rect 294604 202360 294656 202366
rect 294604 202302 294656 202308
rect 294708 201618 294736 509254
rect 295248 497208 295300 497214
rect 295248 497150 295300 497156
rect 295156 393032 295208 393038
rect 295156 392974 295208 392980
rect 294696 201612 294748 201618
rect 294696 201554 294748 201560
rect 293868 201544 293920 201550
rect 293868 201486 293920 201492
rect 294420 201544 294472 201550
rect 294420 201486 294472 201492
rect 294432 200002 294460 201486
rect 295168 200138 295196 392974
rect 295260 201550 295288 497150
rect 295352 406638 295380 521222
rect 295984 520940 296036 520946
rect 295984 520882 296036 520888
rect 295340 406632 295392 406638
rect 295340 406574 295392 406580
rect 295352 405754 295380 406574
rect 295996 406570 296024 520882
rect 295984 406564 296036 406570
rect 295984 406506 296036 406512
rect 295996 406434 296024 406506
rect 295984 406428 296036 406434
rect 295984 406370 296036 406376
rect 295340 405748 295392 405754
rect 295340 405690 295392 405696
rect 296076 405748 296128 405754
rect 296076 405690 296128 405696
rect 296088 395350 296116 405690
rect 296076 395344 296128 395350
rect 296076 395286 296128 395292
rect 296168 202020 296220 202026
rect 296168 201962 296220 201968
rect 295248 201544 295300 201550
rect 295248 201486 295300 201492
rect 295800 201544 295852 201550
rect 295800 201486 295852 201492
rect 294892 200110 295196 200138
rect 294892 200002 294920 200110
rect 295812 200002 295840 201486
rect 296180 200002 296208 201962
rect 296548 200002 296576 531383
rect 296640 201550 296668 565791
rect 296902 563408 296958 563417
rect 296902 563343 296958 563352
rect 296916 563106 296944 563343
rect 296904 563100 296956 563106
rect 296904 563042 296956 563048
rect 297270 556880 297326 556889
rect 297270 556815 297326 556824
rect 297284 556238 297312 556815
rect 297272 556232 297324 556238
rect 297272 556174 297324 556180
rect 297362 541104 297418 541113
rect 297362 541039 297418 541048
rect 297178 522200 297234 522209
rect 297178 522135 297234 522144
rect 297192 521694 297220 522135
rect 297180 521688 297232 521694
rect 297180 521630 297232 521636
rect 297270 519208 297326 519217
rect 297270 519143 297326 519152
rect 297284 518974 297312 519143
rect 297272 518968 297324 518974
rect 297272 518910 297324 518916
rect 297376 337550 297404 541039
rect 297468 534070 297496 572727
rect 298006 570072 298062 570081
rect 298006 570007 298062 570016
rect 298020 569974 298048 570007
rect 298008 569968 298060 569974
rect 298008 569910 298060 569916
rect 298006 544096 298062 544105
rect 298006 544031 298062 544040
rect 297638 538384 297694 538393
rect 297638 538319 297694 538328
rect 297652 538286 297680 538319
rect 297640 538280 297692 538286
rect 297640 538222 297692 538228
rect 297914 534848 297970 534857
rect 297914 534783 297970 534792
rect 297456 534064 297508 534070
rect 297456 534006 297508 534012
rect 297454 528864 297510 528873
rect 297454 528799 297510 528808
rect 297468 518226 297496 528799
rect 297456 518220 297508 518226
rect 297456 518162 297508 518168
rect 297822 516216 297878 516225
rect 297822 516151 297824 516160
rect 297876 516151 297878 516160
rect 297824 516122 297876 516128
rect 297822 513496 297878 513505
rect 297822 513431 297878 513440
rect 297730 509688 297786 509697
rect 297730 509623 297786 509632
rect 297744 509318 297772 509623
rect 297732 509312 297784 509318
rect 297732 509254 297784 509260
rect 297730 506696 297786 506705
rect 297730 506631 297786 506640
rect 297744 506530 297772 506631
rect 297732 506524 297784 506530
rect 297732 506466 297784 506472
rect 297730 503840 297786 503849
rect 297730 503775 297786 503784
rect 297456 386436 297508 386442
rect 297456 386378 297508 386384
rect 297468 383518 297496 386378
rect 297456 383512 297508 383518
rect 297456 383454 297508 383460
rect 297640 375420 297692 375426
rect 297640 375362 297692 375368
rect 297652 375306 297680 375362
rect 297560 375278 297680 375306
rect 297560 370530 297588 375278
rect 297548 370524 297600 370530
rect 297548 370466 297600 370472
rect 297744 357746 297772 503775
rect 297732 357740 297784 357746
rect 297732 357682 297784 357688
rect 297640 357468 297692 357474
rect 297640 357410 297692 357416
rect 297732 357468 297784 357474
rect 297732 357410 297784 357416
rect 297652 356046 297680 357410
rect 297640 356040 297692 356046
rect 297640 355982 297692 355988
rect 297548 346452 297600 346458
rect 297548 346394 297600 346400
rect 297560 340762 297588 346394
rect 297560 340734 297680 340762
rect 297364 337544 297416 337550
rect 297364 337486 297416 337492
rect 297652 323678 297680 340734
rect 297640 323672 297692 323678
rect 297640 323614 297692 323620
rect 297640 318912 297692 318918
rect 297560 318860 297640 318866
rect 297560 318854 297692 318860
rect 297560 318838 297680 318854
rect 297560 311982 297588 318838
rect 297548 311976 297600 311982
rect 297548 311918 297600 311924
rect 297640 311840 297692 311846
rect 297640 311782 297692 311788
rect 297652 307766 297680 311782
rect 297640 307760 297692 307766
rect 297640 307702 297692 307708
rect 297548 298172 297600 298178
rect 297548 298114 297600 298120
rect 297560 298058 297588 298114
rect 297638 298072 297694 298081
rect 297560 298030 297638 298058
rect 297638 298007 297694 298016
rect 297638 288552 297694 288561
rect 297638 288487 297694 288496
rect 297652 288386 297680 288487
rect 297640 288380 297692 288386
rect 297640 288322 297692 288328
rect 297640 270564 297692 270570
rect 297640 270506 297692 270512
rect 297652 270450 297680 270506
rect 297560 270422 297680 270450
rect 297560 263702 297588 270422
rect 297548 263696 297600 263702
rect 297548 263638 297600 263644
rect 297548 260908 297600 260914
rect 297548 260850 297600 260856
rect 297560 260817 297588 260850
rect 297362 260808 297418 260817
rect 297362 260743 297418 260752
rect 297546 260808 297602 260817
rect 297546 260743 297602 260752
rect 297376 251326 297404 260743
rect 297364 251320 297416 251326
rect 297364 251262 297416 251268
rect 297640 251320 297692 251326
rect 297640 251262 297692 251268
rect 297652 244390 297680 251262
rect 297640 244384 297692 244390
rect 297640 244326 297692 244332
rect 297640 244248 297692 244254
rect 297640 244190 297692 244196
rect 297652 241618 297680 244190
rect 297560 241590 297680 241618
rect 297560 240145 297588 241590
rect 297362 240136 297418 240145
rect 297362 240071 297418 240080
rect 297546 240136 297602 240145
rect 297546 240071 297602 240080
rect 297376 230518 297404 240071
rect 297364 230512 297416 230518
rect 297364 230454 297416 230460
rect 297456 230512 297508 230518
rect 297456 230454 297508 230460
rect 297468 222222 297496 230454
rect 297364 222216 297416 222222
rect 297364 222158 297416 222164
rect 297456 222216 297508 222222
rect 297456 222158 297508 222164
rect 297376 212566 297404 222158
rect 297364 212560 297416 212566
rect 297364 212502 297416 212508
rect 297640 212560 297692 212566
rect 297640 212502 297692 212508
rect 297548 210316 297600 210322
rect 297548 210258 297600 210264
rect 297456 202904 297508 202910
rect 297456 202846 297508 202852
rect 296628 201544 296680 201550
rect 297468 201532 297496 202846
rect 297560 201686 297588 210258
rect 297652 202910 297680 212502
rect 297640 202904 297692 202910
rect 297640 202846 297692 202852
rect 297744 201890 297772 357410
rect 297836 308106 297864 513431
rect 297824 308100 297876 308106
rect 297824 308042 297876 308048
rect 297824 307828 297876 307834
rect 297824 307770 297876 307776
rect 297732 201884 297784 201890
rect 297732 201826 297784 201832
rect 297836 201754 297864 307770
rect 297928 210202 297956 534783
rect 298020 210322 298048 544031
rect 298204 520946 298232 582626
rect 298192 520940 298244 520946
rect 298192 520882 298244 520888
rect 298296 499050 298324 582898
rect 298388 499118 298416 583102
rect 298376 499112 298428 499118
rect 298376 499054 298428 499060
rect 298284 499044 298336 499050
rect 298284 498986 298336 498992
rect 298480 498914 298508 583170
rect 302790 582992 302846 583001
rect 302790 582927 302846 582936
rect 298560 582888 298612 582894
rect 298560 582830 298612 582836
rect 298572 498982 298600 582830
rect 300492 582752 300544 582758
rect 298834 582720 298890 582729
rect 300492 582694 300544 582700
rect 298834 582655 298890 582664
rect 298652 582548 298704 582554
rect 298652 582490 298704 582496
rect 298560 498976 298612 498982
rect 298560 498918 298612 498924
rect 298468 498908 298520 498914
rect 298468 498850 298520 498856
rect 298664 498846 298692 582490
rect 298744 582480 298796 582486
rect 298744 582422 298796 582428
rect 298652 498840 298704 498846
rect 298652 498782 298704 498788
rect 298652 393168 298704 393174
rect 298652 393110 298704 393116
rect 298560 210452 298612 210458
rect 298560 210394 298612 210400
rect 298008 210316 298060 210322
rect 298008 210258 298060 210264
rect 297928 210174 298048 210202
rect 297916 202768 297968 202774
rect 297916 202710 297968 202716
rect 297824 201748 297876 201754
rect 297824 201690 297876 201696
rect 297548 201680 297600 201686
rect 297548 201622 297600 201628
rect 297468 201504 297588 201532
rect 296628 201486 296680 201492
rect 297560 200002 297588 201504
rect 297928 200002 297956 202710
rect 298020 202434 298048 210174
rect 298008 202428 298060 202434
rect 298008 202370 298060 202376
rect 298572 202366 298600 210394
rect 298664 202842 298692 393110
rect 298652 202836 298704 202842
rect 298652 202778 298704 202784
rect 298756 202502 298784 582422
rect 298848 202774 298876 582655
rect 300400 582412 300452 582418
rect 300400 582354 300452 582360
rect 299388 579692 299440 579698
rect 299388 579634 299440 579640
rect 299294 560416 299350 560425
rect 299294 560351 299350 560360
rect 299202 553616 299258 553625
rect 299202 553551 299258 553560
rect 299110 550760 299166 550769
rect 299110 550695 299166 550704
rect 299018 547904 299074 547913
rect 299018 547839 299074 547848
rect 298926 525872 298982 525881
rect 298926 525807 298982 525816
rect 298836 202768 298888 202774
rect 298836 202710 298888 202716
rect 298940 202570 298968 525807
rect 299032 210458 299060 547839
rect 299020 210452 299072 210458
rect 299020 210394 299072 210400
rect 299124 210338 299152 550695
rect 299032 210310 299152 210338
rect 298928 202564 298980 202570
rect 298928 202506 298980 202512
rect 298744 202496 298796 202502
rect 298744 202438 298796 202444
rect 298560 202360 298612 202366
rect 298560 202302 298612 202308
rect 299032 202094 299060 210310
rect 299112 202836 299164 202842
rect 299112 202778 299164 202784
rect 299020 202088 299072 202094
rect 299020 202030 299072 202036
rect 298376 201952 298428 201958
rect 298376 201894 298428 201900
rect 298388 200002 298416 201894
rect 298652 201816 298704 201822
rect 298652 201758 298704 201764
rect 292316 199974 292468 200002
rect 292928 199974 293080 200002
rect 293756 199974 293816 200002
rect 294216 199974 294460 200002
rect 294584 199974 294920 200002
rect 295504 199974 295840 200002
rect 295964 199974 296208 200002
rect 296332 199974 296576 200002
rect 297252 199974 297588 200002
rect 297712 199974 297956 200002
rect 298080 199974 298416 200002
rect 298664 200002 298692 201758
rect 299124 200002 299152 202778
rect 299216 202706 299244 553551
rect 299204 202700 299256 202706
rect 299204 202642 299256 202648
rect 299308 202502 299336 560351
rect 299400 202638 299428 579634
rect 299480 579352 299532 579358
rect 299480 579294 299532 579300
rect 299492 202774 299520 579294
rect 300412 498642 300440 582354
rect 300504 499186 300532 582694
rect 302804 579972 302832 582927
rect 307036 579972 307064 583646
rect 319720 583636 319772 583642
rect 319720 583578 319772 583584
rect 311256 583568 311308 583574
rect 311256 583510 311308 583516
rect 309232 582412 309284 582418
rect 309232 582354 309284 582360
rect 309244 579972 309272 582354
rect 311268 579972 311296 583510
rect 313464 582616 313516 582622
rect 313464 582558 313516 582564
rect 313476 579972 313504 582558
rect 319732 579972 319760 583578
rect 330392 583500 330444 583506
rect 330392 583442 330444 583448
rect 326160 583024 326212 583030
rect 326160 582966 326212 582972
rect 324134 582584 324190 582593
rect 321928 582548 321980 582554
rect 324134 582519 324190 582528
rect 321928 582490 321980 582496
rect 321940 579972 321968 582490
rect 324148 579972 324176 582519
rect 326172 579972 326200 582966
rect 328368 582480 328420 582486
rect 328368 582422 328420 582428
rect 328380 579972 328408 582422
rect 330404 579972 330432 583442
rect 347504 583432 347556 583438
rect 347504 583374 347556 583380
rect 336832 583364 336884 583370
rect 336832 583306 336884 583312
rect 334624 583296 334676 583302
rect 334624 583238 334676 583244
rect 332600 583228 332652 583234
rect 332600 583170 332652 583176
rect 332612 579972 332640 583170
rect 334636 579972 334664 583238
rect 336844 579972 336872 583306
rect 341064 583160 341116 583166
rect 341064 583102 341116 583108
rect 338856 583092 338908 583098
rect 338856 583034 338908 583040
rect 338868 579972 338896 583034
rect 341076 579972 341104 583102
rect 345296 582684 345348 582690
rect 345296 582626 345348 582632
rect 345308 579972 345336 582626
rect 347516 579972 347544 583374
rect 353760 582956 353812 582962
rect 353760 582898 353812 582904
rect 351736 582820 351788 582826
rect 351736 582762 351788 582768
rect 349526 582448 349582 582457
rect 349526 582383 349582 582392
rect 349540 579972 349568 582383
rect 351748 579972 351776 582762
rect 353772 579972 353800 582898
rect 355968 582888 356020 582894
rect 355968 582830 356020 582836
rect 368662 582856 368718 582865
rect 355980 579972 356008 582830
rect 368662 582791 368718 582800
rect 362408 582752 362460 582758
rect 360198 582720 360254 582729
rect 362408 582694 362460 582700
rect 360198 582655 360254 582664
rect 357992 582616 358044 582622
rect 357992 582558 358044 582564
rect 358004 579972 358032 582558
rect 360212 579972 360240 582655
rect 362420 579972 362448 582694
rect 366640 582684 366692 582690
rect 366640 582626 366692 582632
rect 366652 579972 366680 582626
rect 368676 579972 368704 582791
rect 378232 582684 378284 582690
rect 378232 582626 378284 582632
rect 370872 582548 370924 582554
rect 370872 582490 370924 582496
rect 370884 579972 370912 582490
rect 372896 582412 372948 582418
rect 372896 582354 372948 582360
rect 372908 579972 372936 582354
rect 304828 579698 305026 579714
rect 304816 579692 305026 579698
rect 304868 579686 305026 579692
rect 304816 579634 304868 579640
rect 300676 579352 300728 579358
rect 300610 579300 300676 579306
rect 300610 579294 300728 579300
rect 315212 579352 315264 579358
rect 317420 579352 317472 579358
rect 315264 579300 315514 579306
rect 315212 579294 315514 579300
rect 342996 579352 343048 579358
rect 317472 579300 317722 579306
rect 317420 579294 317722 579300
rect 364248 579352 364300 579358
rect 343048 579300 343298 579306
rect 342996 579294 343298 579300
rect 375380 579352 375432 579358
rect 364300 579300 364458 579306
rect 364248 579294 364458 579300
rect 300610 579278 300716 579294
rect 315224 579278 315514 579294
rect 317432 579278 317722 579294
rect 343008 579278 343298 579294
rect 364260 579278 364458 579294
rect 375130 579300 375380 579306
rect 375130 579294 375432 579300
rect 375130 579278 375420 579294
rect 377154 579278 377260 579306
rect 300610 500126 300716 500154
rect 302634 500126 302924 500154
rect 304842 500126 304948 500154
rect 300492 499180 300544 499186
rect 300492 499122 300544 499128
rect 300400 498636 300452 498642
rect 300400 498578 300452 498584
rect 300688 495394 300716 500126
rect 302896 499526 302924 500126
rect 302884 499520 302936 499526
rect 302884 499462 302936 499468
rect 302240 498636 302292 498642
rect 302240 498578 302292 498584
rect 301504 497276 301556 497282
rect 301504 497218 301556 497224
rect 300596 495366 300716 495394
rect 300596 485858 300624 495366
rect 299756 485852 299808 485858
rect 299756 485794 299808 485800
rect 300584 485852 300636 485858
rect 300584 485794 300636 485800
rect 299768 476134 299796 485794
rect 299572 476128 299624 476134
rect 299756 476128 299808 476134
rect 299624 476076 299704 476082
rect 299572 476070 299704 476076
rect 299756 476070 299808 476076
rect 299584 476054 299704 476070
rect 299676 473346 299704 476054
rect 299664 473340 299716 473346
rect 299664 473282 299716 473288
rect 299664 466404 299716 466410
rect 299664 466346 299716 466352
rect 299676 463706 299704 466346
rect 299676 463678 299796 463706
rect 299768 456822 299796 463678
rect 299572 456816 299624 456822
rect 299756 456816 299808 456822
rect 299624 456764 299704 456770
rect 299572 456758 299704 456764
rect 299756 456758 299808 456764
rect 299584 456742 299704 456758
rect 299676 454034 299704 456742
rect 299664 454028 299716 454034
rect 299664 453970 299716 453976
rect 299664 447092 299716 447098
rect 299664 447034 299716 447040
rect 299676 444394 299704 447034
rect 299676 444366 299796 444394
rect 299768 437510 299796 444366
rect 299572 437504 299624 437510
rect 299756 437504 299808 437510
rect 299624 437452 299704 437458
rect 299572 437446 299704 437452
rect 299756 437446 299808 437452
rect 299584 437430 299704 437446
rect 299676 434722 299704 437430
rect 299664 434716 299716 434722
rect 299664 434658 299716 434664
rect 299664 427780 299716 427786
rect 299664 427722 299716 427728
rect 299676 425082 299704 427722
rect 299676 425054 299796 425082
rect 299768 418198 299796 425054
rect 299572 418192 299624 418198
rect 299756 418192 299808 418198
rect 299624 418140 299704 418146
rect 299572 418134 299704 418140
rect 299756 418134 299808 418140
rect 299584 418118 299704 418134
rect 299676 415410 299704 418118
rect 299664 415404 299716 415410
rect 299664 415346 299716 415352
rect 299756 405748 299808 405754
rect 299756 405690 299808 405696
rect 299768 398834 299796 405690
rect 299584 398806 299796 398834
rect 299584 396030 299612 398806
rect 299572 396024 299624 396030
rect 299572 395966 299624 395972
rect 300768 393236 300820 393242
rect 300768 393178 300820 393184
rect 300676 392488 300728 392494
rect 300676 392430 300728 392436
rect 299664 386436 299716 386442
rect 299664 386378 299716 386384
rect 299676 379522 299704 386378
rect 299584 379494 299704 379522
rect 299584 379386 299612 379494
rect 299584 379358 299704 379386
rect 299676 362302 299704 379358
rect 299664 362296 299716 362302
rect 299664 362238 299716 362244
rect 299756 357468 299808 357474
rect 299756 357410 299808 357416
rect 299768 337482 299796 357410
rect 299756 337476 299808 337482
rect 299756 337418 299808 337424
rect 300124 202836 300176 202842
rect 300124 202778 300176 202784
rect 299480 202768 299532 202774
rect 299480 202710 299532 202716
rect 299388 202632 299440 202638
rect 299388 202574 299440 202580
rect 299296 202496 299348 202502
rect 299296 202438 299348 202444
rect 300136 200002 300164 202778
rect 298664 199974 299000 200002
rect 299124 199974 299368 200002
rect 299828 199974 300164 200002
rect 300688 200002 300716 392430
rect 300780 202842 300808 393178
rect 300768 202836 300820 202842
rect 300768 202778 300820 202784
rect 301412 202836 301464 202842
rect 301412 202778 301464 202784
rect 301424 200002 301452 202778
rect 301516 202026 301544 497218
rect 302148 393304 302200 393310
rect 302148 393246 302200 393252
rect 302056 392556 302108 392562
rect 302056 392498 302108 392504
rect 301872 208548 301924 208554
rect 301872 208490 301924 208496
rect 301504 202020 301556 202026
rect 301504 201962 301556 201968
rect 301884 200002 301912 208490
rect 302068 202842 302096 392498
rect 302160 208554 302188 393246
rect 302148 208548 302200 208554
rect 302148 208490 302200 208496
rect 302056 202836 302108 202842
rect 302056 202778 302108 202784
rect 300688 199974 300748 200002
rect 301116 199974 301452 200002
rect 301576 199974 301912 200002
rect 302252 200002 302280 498578
rect 302896 391270 302924 499462
rect 304264 496936 304316 496942
rect 304264 496878 304316 496884
rect 302884 391264 302936 391270
rect 302884 391206 302936 391212
rect 302896 338094 302924 391206
rect 302884 338088 302936 338094
rect 302884 338030 302936 338036
rect 303080 202694 303292 202722
rect 303080 202570 303108 202694
rect 303068 202564 303120 202570
rect 303068 202506 303120 202512
rect 303160 202564 303212 202570
rect 303160 202506 303212 202512
rect 303172 200002 303200 202506
rect 302252 199974 302404 200002
rect 302864 199974 303200 200002
rect 303264 200002 303292 202694
rect 304276 202570 304304 496878
rect 304920 202706 304948 500126
rect 306472 498840 306524 498846
rect 306472 498782 306524 498788
rect 304356 202700 304408 202706
rect 304356 202642 304408 202648
rect 304908 202700 304960 202706
rect 304908 202642 304960 202648
rect 304264 202564 304316 202570
rect 304264 202506 304316 202512
rect 303896 201748 303948 201754
rect 303896 201690 303948 201696
rect 303908 200002 303936 201690
rect 304368 200002 304396 202642
rect 305000 202360 305052 202366
rect 305000 202302 305052 202308
rect 305012 200002 305040 202302
rect 306484 201754 306512 498782
rect 306852 496874 306880 500004
rect 308968 499990 309074 500018
rect 308968 496874 308996 499990
rect 310612 499112 310664 499118
rect 310612 499054 310664 499060
rect 309140 498908 309192 498914
rect 309140 498850 309192 498856
rect 310428 498908 310480 498914
rect 310428 498850 310480 498856
rect 309048 498840 309100 498846
rect 309048 498782 309100 498788
rect 306840 496868 306892 496874
rect 306840 496810 306892 496816
rect 308956 496868 309008 496874
rect 308956 496810 309008 496816
rect 307668 394052 307720 394058
rect 307668 393994 307720 394000
rect 307680 202570 307708 393994
rect 308956 392420 309008 392426
rect 308956 392362 309008 392368
rect 308864 215280 308916 215286
rect 308864 215222 308916 215228
rect 308876 205714 308904 215222
rect 308784 205686 308904 205714
rect 306656 202564 306708 202570
rect 306656 202506 306708 202512
rect 307668 202564 307720 202570
rect 307668 202506 307720 202512
rect 306472 201748 306524 201754
rect 306472 201690 306524 201696
rect 305644 201680 305696 201686
rect 305644 201622 305696 201628
rect 305656 200002 305684 201622
rect 306668 200002 306696 202506
rect 307300 201748 307352 201754
rect 307300 201690 307352 201696
rect 307024 201544 307076 201550
rect 307024 201486 307076 201492
rect 307036 200002 307064 201486
rect 303264 199974 303324 200002
rect 303908 199974 304152 200002
rect 304368 199974 304612 200002
rect 305012 199974 305072 200002
rect 305656 199974 305900 200002
rect 306360 199974 306696 200002
rect 306820 199974 307064 200002
rect 307312 200002 307340 201690
rect 308404 201612 308456 201618
rect 308404 201554 308456 201560
rect 308416 200002 308444 201554
rect 308784 200002 308812 205686
rect 308968 201618 308996 392362
rect 309060 215286 309088 498782
rect 309048 215280 309100 215286
rect 309048 215222 309100 215228
rect 309152 202842 309180 498850
rect 309140 202836 309192 202842
rect 309140 202778 309192 202784
rect 309600 202836 309652 202842
rect 309600 202778 309652 202784
rect 309140 202700 309192 202706
rect 309140 202642 309192 202648
rect 308956 201612 309008 201618
rect 308956 201554 309008 201560
rect 307312 199974 307648 200002
rect 308108 199974 308444 200002
rect 308568 199974 308812 200002
rect 309152 200002 309180 202642
rect 309612 200002 309640 202778
rect 310440 200002 310468 498850
rect 310624 202434 310652 499054
rect 311084 497010 311112 500004
rect 311900 499180 311952 499186
rect 311900 499122 311952 499128
rect 311072 497004 311124 497010
rect 311072 496946 311124 496952
rect 311912 202842 311940 499122
rect 313292 498137 313320 500004
rect 314672 499990 315330 500018
rect 313278 498128 313334 498137
rect 313278 498063 313334 498072
rect 314568 392352 314620 392358
rect 314568 392294 314620 392300
rect 314580 202842 314608 392294
rect 311900 202836 311952 202842
rect 311900 202778 311952 202784
rect 312544 202836 312596 202842
rect 312544 202778 312596 202784
rect 313556 202836 313608 202842
rect 313556 202778 313608 202784
rect 314568 202836 314620 202842
rect 314568 202778 314620 202784
rect 311164 202700 311216 202706
rect 311164 202642 311216 202648
rect 310612 202428 310664 202434
rect 310612 202370 310664 202376
rect 311176 200002 311204 202642
rect 311256 202428 311308 202434
rect 311256 202370 311308 202376
rect 309152 199974 309396 200002
rect 309612 199974 309856 200002
rect 310316 199974 310468 200002
rect 311144 199974 311204 200002
rect 311268 200002 311296 202370
rect 311992 202088 312044 202094
rect 311992 202030 312044 202036
rect 312004 200002 312032 202030
rect 311268 199974 311604 200002
rect 311972 199974 312032 200002
rect 312556 200002 312584 202778
rect 313568 200002 313596 202778
rect 313648 202768 313700 202774
rect 313648 202710 313700 202716
rect 312556 199974 312892 200002
rect 313352 199974 313596 200002
rect 313660 200002 313688 202710
rect 314672 201618 314700 499990
rect 314752 499044 314804 499050
rect 314752 498986 314804 498992
rect 314764 202842 314792 498986
rect 316040 498976 316092 498982
rect 316040 498918 316092 498924
rect 317328 498976 317380 498982
rect 317328 498918 317380 498924
rect 315948 394120 316000 394126
rect 315948 394062 316000 394068
rect 314752 202836 314804 202842
rect 314752 202778 314804 202784
rect 315580 202836 315632 202842
rect 315580 202778 315632 202784
rect 315304 202088 315356 202094
rect 315304 202030 315356 202036
rect 314936 201816 314988 201822
rect 314936 201758 314988 201764
rect 314660 201612 314712 201618
rect 314660 201554 314712 201560
rect 314948 200002 314976 201758
rect 315316 200002 315344 202030
rect 315396 202020 315448 202026
rect 315396 201962 315448 201968
rect 313660 199974 313720 200002
rect 314640 199974 314976 200002
rect 315100 199974 315344 200002
rect 315408 200002 315436 201962
rect 315592 200002 315620 202778
rect 315960 201822 315988 394062
rect 315948 201816 316000 201822
rect 315948 201758 316000 201764
rect 316052 201550 316080 498918
rect 316684 496868 316736 496874
rect 316684 496810 316736 496816
rect 316696 202842 316724 496810
rect 316684 202836 316736 202842
rect 316684 202778 316736 202784
rect 317340 201634 317368 498918
rect 317524 497146 317552 500004
rect 319732 497894 319760 500004
rect 321468 499044 321520 499050
rect 321468 498986 321520 498992
rect 319720 497888 319772 497894
rect 319720 497830 319772 497836
rect 320088 497888 320140 497894
rect 320088 497830 320140 497836
rect 317512 497140 317564 497146
rect 317512 497082 317564 497088
rect 319444 497140 319496 497146
rect 319444 497082 319496 497088
rect 318616 202768 318668 202774
rect 318616 202710 318668 202716
rect 317064 201606 317368 201634
rect 316040 201544 316092 201550
rect 316040 201486 316092 201492
rect 317064 200002 317092 201606
rect 317144 201544 317196 201550
rect 317144 201486 317196 201492
rect 315408 199974 315468 200002
rect 315592 199974 315928 200002
rect 316756 199974 317092 200002
rect 317156 200002 317184 201486
rect 318628 200002 318656 202710
rect 319456 202094 319484 497082
rect 319444 202088 319496 202094
rect 319444 202030 319496 202036
rect 320100 201550 320128 497830
rect 320640 202632 320692 202638
rect 320640 202574 320692 202580
rect 319076 201544 319128 201550
rect 319076 201486 319128 201492
rect 320088 201544 320140 201550
rect 320088 201486 320140 201492
rect 320548 201544 320600 201550
rect 320548 201486 320600 201492
rect 319088 200002 319116 201486
rect 320560 200002 320588 201486
rect 317156 199974 317216 200002
rect 318504 199974 318656 200002
rect 318964 199974 319116 200002
rect 320252 199974 320588 200002
rect 320652 200002 320680 202574
rect 321480 201550 321508 498986
rect 321756 497078 321784 500004
rect 321744 497072 321796 497078
rect 321744 497014 321796 497020
rect 323964 496874 323992 500004
rect 325712 499990 326002 500018
rect 327092 499990 328210 500018
rect 329852 499990 330234 500018
rect 324228 499112 324280 499118
rect 324228 499054 324280 499060
rect 322204 496868 322256 496874
rect 322204 496810 322256 496816
rect 323952 496868 324004 496874
rect 323952 496810 324004 496816
rect 321652 202836 321704 202842
rect 321652 202778 321704 202784
rect 321468 201544 321520 201550
rect 321468 201486 321520 201492
rect 321664 200002 321692 202778
rect 322216 202230 322244 496810
rect 322848 392284 322900 392290
rect 322848 392226 322900 392232
rect 322204 202224 322256 202230
rect 322204 202166 322256 202172
rect 322860 200138 322888 392226
rect 324044 201544 324096 201550
rect 324044 201486 324096 201492
rect 322768 200110 322888 200138
rect 322768 200002 322796 200110
rect 324056 200002 324084 201486
rect 324240 200002 324268 499054
rect 325712 202570 325740 499990
rect 325700 202564 325752 202570
rect 325700 202506 325752 202512
rect 325148 202496 325200 202502
rect 325148 202438 325200 202444
rect 320652 199974 320712 200002
rect 321664 199974 322000 200002
rect 322460 199974 322796 200002
rect 323748 199974 324084 200002
rect 324208 199974 324268 200002
rect 325160 200002 325188 202438
rect 325700 202428 325752 202434
rect 325700 202370 325752 202376
rect 325712 200002 325740 202370
rect 327092 201550 327120 499990
rect 329852 337414 329880 499990
rect 332428 496942 332456 500004
rect 334452 497962 334480 500004
rect 334440 497956 334492 497962
rect 334440 497898 334492 497904
rect 334624 497072 334676 497078
rect 334624 497014 334676 497020
rect 333244 497004 333296 497010
rect 333244 496946 333296 496952
rect 332416 496936 332468 496942
rect 332416 496878 332468 496884
rect 330484 496868 330536 496874
rect 330484 496810 330536 496816
rect 329840 337408 329892 337414
rect 329840 337350 329892 337356
rect 330496 202706 330524 496810
rect 333256 202774 333284 496946
rect 333888 374060 333940 374066
rect 333888 374002 333940 374008
rect 333796 358080 333848 358086
rect 333796 358022 333848 358028
rect 333244 202768 333296 202774
rect 333244 202710 333296 202716
rect 330484 202700 330536 202706
rect 330484 202642 330536 202648
rect 333152 202428 333204 202434
rect 333152 202370 333204 202376
rect 332508 202224 332560 202230
rect 332508 202166 332560 202172
rect 327080 201544 327132 201550
rect 327080 201486 327132 201492
rect 332520 200002 332548 202166
rect 333164 200002 333192 202370
rect 333808 200138 333836 358022
rect 333900 202434 333928 374002
rect 333888 202428 333940 202434
rect 333888 202370 333940 202376
rect 334636 202366 334664 497014
rect 336660 496874 336688 500004
rect 338868 498030 338896 500004
rect 338856 498024 338908 498030
rect 338856 497966 338908 497972
rect 337476 497956 337528 497962
rect 337476 497898 337528 497904
rect 336648 496868 336700 496874
rect 336648 496810 336700 496816
rect 337384 496868 337436 496874
rect 337384 496810 337436 496816
rect 334624 202360 334676 202366
rect 334624 202302 334676 202308
rect 337396 202298 337424 496810
rect 337384 202292 337436 202298
rect 337384 202234 337436 202240
rect 337488 202162 337516 497898
rect 340892 497214 340920 500004
rect 340880 497208 340932 497214
rect 340880 497150 340932 497156
rect 343100 496874 343128 500004
rect 345124 497418 345152 500004
rect 347332 498098 347360 500004
rect 347320 498092 347372 498098
rect 347320 498034 347372 498040
rect 345112 497412 345164 497418
rect 345112 497354 345164 497360
rect 349356 497146 349384 500004
rect 351564 497350 351592 500004
rect 351552 497344 351604 497350
rect 351552 497286 351604 497292
rect 353588 497282 353616 500004
rect 353576 497276 353628 497282
rect 353576 497218 353628 497224
rect 349344 497140 349396 497146
rect 349344 497082 349396 497088
rect 355796 497010 355824 500004
rect 358004 497894 358032 500004
rect 357992 497888 358044 497894
rect 357992 497830 358044 497836
rect 360028 497554 360056 500004
rect 360016 497548 360068 497554
rect 360016 497490 360068 497496
rect 362236 497078 362264 500004
rect 364260 498166 364288 500004
rect 364248 498160 364300 498166
rect 364248 498102 364300 498108
rect 366468 497826 366496 500004
rect 366456 497820 366508 497826
rect 366456 497762 366508 497768
rect 368492 497758 368520 500004
rect 370700 497962 370728 500004
rect 370688 497956 370740 497962
rect 370688 497898 370740 497904
rect 368480 497752 368532 497758
rect 368480 497694 368532 497700
rect 372724 497486 372752 500004
rect 374932 497622 374960 500004
rect 377140 497690 377168 500004
rect 377128 497684 377180 497690
rect 377128 497626 377180 497632
rect 374920 497616 374972 497622
rect 374920 497558 374972 497564
rect 372712 497480 372764 497486
rect 372712 497422 372764 497428
rect 362224 497072 362276 497078
rect 362224 497014 362276 497020
rect 355784 497004 355836 497010
rect 355784 496946 355836 496952
rect 343088 496868 343140 496874
rect 343088 496810 343140 496816
rect 358084 407176 358136 407182
rect 358084 407118 358136 407124
rect 344284 406428 344336 406434
rect 344284 406370 344336 406376
rect 344296 395418 344324 406370
rect 349068 395480 349120 395486
rect 349068 395422 349120 395428
rect 344284 395412 344336 395418
rect 344284 395354 344336 395360
rect 344928 395276 344980 395282
rect 344928 395218 344980 395224
rect 343548 394868 343600 394874
rect 343548 394810 343600 394816
rect 342168 358216 342220 358222
rect 342168 358158 342220 358164
rect 342180 202842 342208 358158
rect 341340 202836 341392 202842
rect 341340 202778 341392 202784
rect 342168 202836 342220 202842
rect 342168 202778 342220 202784
rect 337476 202156 337528 202162
rect 337476 202098 337528 202104
rect 333532 200110 333836 200138
rect 333532 200002 333560 200110
rect 341352 200002 341380 202778
rect 342076 202156 342128 202162
rect 342076 202098 342128 202104
rect 342088 200002 342116 202098
rect 343560 200546 343588 394810
rect 344008 202292 344060 202298
rect 344008 202234 344060 202240
rect 343284 200518 343588 200546
rect 343284 200138 343312 200518
rect 343192 200110 343312 200138
rect 343192 200002 343220 200110
rect 344020 200002 344048 202234
rect 344940 200002 344968 395218
rect 347688 394936 347740 394942
rect 347688 394878 347740 394884
rect 346676 202564 346728 202570
rect 346676 202506 346728 202512
rect 345756 202360 345808 202366
rect 345756 202302 345808 202308
rect 345768 200002 345796 202302
rect 346688 200002 346716 202506
rect 347700 200138 347728 394878
rect 348332 202428 348384 202434
rect 348332 202370 348384 202376
rect 347516 200110 347728 200138
rect 347516 200002 347544 200110
rect 348344 200002 348372 202370
rect 349080 200002 349108 395422
rect 355968 395208 356020 395214
rect 355968 395150 356020 395156
rect 355876 395140 355928 395146
rect 355876 395082 355928 395088
rect 353208 395072 353260 395078
rect 353208 395014 353260 395020
rect 351828 387864 351880 387870
rect 351828 387806 351880 387812
rect 351184 380928 351236 380934
rect 351184 380870 351236 380876
rect 350448 358284 350500 358290
rect 350448 358226 350500 358232
rect 350460 200138 350488 358226
rect 351196 202570 351224 380870
rect 351184 202564 351236 202570
rect 351184 202506 351236 202512
rect 351736 202088 351788 202094
rect 351736 202030 351788 202036
rect 351000 201748 351052 201754
rect 351000 201690 351052 201696
rect 350092 200110 350488 200138
rect 350092 200002 350120 200110
rect 351012 200002 351040 201690
rect 351748 200002 351776 202030
rect 351840 201754 351868 387806
rect 353220 202502 353248 395014
rect 354588 358352 354640 358358
rect 354588 358294 354640 358300
rect 352748 202496 352800 202502
rect 352748 202438 352800 202444
rect 353208 202496 353260 202502
rect 353208 202438 353260 202444
rect 351828 201748 351880 201754
rect 351828 201690 351880 201696
rect 352760 200002 352788 202438
rect 353576 201680 353628 201686
rect 353576 201622 353628 201628
rect 353588 200002 353616 201622
rect 354600 200138 354628 358294
rect 355324 201748 355376 201754
rect 355324 201690 355376 201696
rect 354508 200110 354628 200138
rect 354508 200002 354536 200110
rect 355336 200002 355364 201690
rect 325160 199974 325496 200002
rect 325712 199974 325956 200002
rect 332488 199974 332548 200002
rect 332856 199974 333192 200002
rect 333316 199974 333560 200002
rect 341136 199974 341380 200002
rect 342056 199974 342116 200002
rect 342884 199974 343220 200002
rect 343712 199974 344048 200002
rect 344632 199974 344968 200002
rect 345460 199974 345796 200002
rect 346380 199974 346716 200002
rect 347208 199974 347544 200002
rect 348128 199974 348372 200002
rect 348956 199974 349108 200002
rect 349876 199974 350120 200002
rect 350704 199974 351040 200002
rect 351624 199974 351776 200002
rect 352452 199974 352788 200002
rect 353280 199974 353616 200002
rect 354200 199974 354536 200002
rect 355028 199974 355364 200002
rect 355888 200002 355916 395082
rect 355980 201754 356008 395150
rect 357438 391368 357494 391377
rect 357438 391303 357494 391312
rect 357452 391270 357480 391303
rect 357440 391264 357492 391270
rect 357440 391206 357492 391212
rect 357440 387864 357492 387870
rect 357438 387832 357440 387841
rect 357492 387832 357494 387841
rect 357438 387767 357494 387776
rect 357348 386572 357400 386578
rect 357348 386514 357400 386520
rect 357360 386374 357388 386514
rect 357348 386368 357400 386374
rect 357348 386310 357400 386316
rect 357438 381032 357494 381041
rect 357438 380967 357494 380976
rect 357452 380934 357480 380967
rect 357440 380928 357492 380934
rect 357440 380870 357492 380876
rect 358096 377777 358124 407118
rect 361856 395480 361908 395486
rect 361856 395422 361908 395428
rect 360016 394800 360068 394806
rect 360016 394742 360068 394748
rect 358542 384568 358598 384577
rect 358542 384503 358598 384512
rect 358082 377768 358138 377777
rect 358082 377703 358138 377712
rect 357164 376780 357216 376786
rect 357164 376722 357216 376728
rect 357176 376666 357204 376722
rect 357176 376650 357296 376666
rect 357176 376644 357308 376650
rect 357176 376638 357256 376644
rect 357256 376586 357308 376592
rect 357438 374232 357494 374241
rect 357438 374167 357494 374176
rect 357452 374066 357480 374167
rect 357440 374060 357492 374066
rect 357440 374002 357492 374008
rect 358082 370968 358138 370977
rect 358082 370903 358138 370912
rect 357348 367124 357400 367130
rect 357348 367066 357400 367072
rect 356702 364168 356758 364177
rect 356702 364103 356758 364112
rect 355968 201748 356020 201754
rect 355968 201690 356020 201696
rect 356716 201686 356744 364103
rect 357360 280294 357388 367066
rect 358096 340610 358124 370903
rect 358174 367432 358230 367441
rect 358174 367367 358230 367376
rect 358188 340746 358216 367367
rect 358556 364410 358584 384503
rect 358544 364404 358596 364410
rect 358544 364346 358596 364352
rect 358728 364404 358780 364410
rect 358728 364346 358780 364352
rect 358740 354634 358768 364346
rect 360028 360194 360056 394742
rect 360108 394732 360160 394738
rect 360108 394674 360160 394680
rect 360016 360188 360068 360194
rect 360016 360130 360068 360136
rect 360120 360126 360148 394674
rect 361868 393380 361896 395422
rect 364248 395344 364300 395350
rect 364248 395286 364300 395292
rect 364260 393380 364288 395286
rect 375656 395140 375708 395146
rect 375656 395082 375708 395088
rect 373448 394936 373500 394942
rect 373448 394878 373500 394884
rect 371056 394868 371108 394874
rect 371056 394810 371108 394816
rect 368848 394800 368900 394806
rect 368848 394742 368900 394748
rect 366456 394732 366508 394738
rect 366456 394674 366508 394680
rect 366468 393380 366496 394674
rect 368860 393380 368888 394742
rect 371068 393380 371096 394810
rect 373460 393380 373488 394878
rect 375668 393380 375696 395082
rect 377232 392834 377260 579278
rect 377402 575512 377458 575521
rect 377402 575447 377458 575456
rect 377310 565856 377366 565865
rect 377310 565791 377366 565800
rect 377036 392828 377088 392834
rect 377036 392770 377088 392776
rect 377220 392828 377272 392834
rect 377220 392770 377272 392776
rect 377048 392714 377076 392770
rect 377324 392714 377352 565791
rect 377416 407862 377444 575447
rect 378138 557220 378194 557229
rect 378138 557155 378194 557164
rect 377494 537568 377550 537577
rect 377494 537503 377550 537512
rect 377404 407856 377456 407862
rect 377404 407798 377456 407804
rect 377508 392970 377536 537503
rect 378048 395072 378100 395078
rect 378048 395014 378100 395020
rect 378060 393380 378088 395014
rect 377496 392964 377548 392970
rect 377496 392906 377548 392912
rect 378152 392902 378180 557155
rect 378244 498982 378272 582626
rect 378416 582616 378468 582622
rect 378416 582558 378468 582564
rect 378324 579352 378376 579358
rect 378324 579294 378376 579300
rect 378336 499050 378364 579294
rect 378428 499118 378456 582558
rect 378600 582548 378652 582554
rect 378600 582490 378652 582496
rect 378508 582412 378560 582418
rect 378508 582354 378560 582360
rect 378416 499112 378468 499118
rect 378416 499054 378468 499060
rect 378324 499044 378376 499050
rect 378324 498986 378376 498992
rect 378232 498976 378284 498982
rect 378232 498918 378284 498924
rect 378520 498846 378548 582354
rect 378612 498914 378640 582490
rect 380714 569120 380770 569129
rect 380714 569055 380770 569064
rect 379702 550760 379758 550769
rect 379702 550695 379758 550704
rect 379518 519208 379574 519217
rect 379518 519143 379574 519152
rect 379532 506682 379560 519143
rect 379440 506654 379560 506682
rect 379440 500886 379468 506654
rect 379518 506560 379574 506569
rect 379518 506495 379574 506504
rect 379532 500954 379560 506495
rect 379520 500948 379572 500954
rect 379520 500890 379572 500896
rect 379428 500880 379480 500886
rect 379428 500822 379480 500828
rect 378600 498908 378652 498914
rect 378600 498850 378652 498856
rect 378508 498840 378560 498846
rect 378508 498782 378560 498788
rect 379520 398676 379572 398682
rect 379520 398618 379572 398624
rect 379532 394754 379560 398618
rect 379440 394726 379560 394754
rect 379440 394058 379468 394726
rect 379518 394632 379574 394641
rect 379518 394567 379574 394576
rect 379428 394052 379480 394058
rect 379428 393994 379480 394000
rect 379428 393508 379480 393514
rect 379428 393450 379480 393456
rect 379440 392902 379468 393450
rect 379532 393038 379560 394567
rect 379610 394496 379666 394505
rect 379610 394431 379666 394440
rect 379520 393032 379572 393038
rect 379520 392974 379572 392980
rect 379624 392902 379652 394431
rect 379716 393514 379744 550695
rect 379794 547088 379850 547097
rect 379794 547023 379850 547032
rect 379704 393508 379756 393514
rect 379704 393450 379756 393456
rect 379704 393372 379756 393378
rect 379704 393314 379756 393320
rect 378140 392896 378192 392902
rect 378140 392838 378192 392844
rect 379428 392896 379480 392902
rect 379428 392838 379480 392844
rect 379612 392896 379664 392902
rect 379612 392838 379664 392844
rect 379716 392834 379744 393314
rect 379808 393242 379836 547023
rect 379886 543824 379942 543833
rect 379886 543759 379942 543768
rect 379796 393236 379848 393242
rect 379796 393178 379848 393184
rect 379900 392834 379928 543759
rect 379978 534576 380034 534585
rect 379978 534511 380034 534520
rect 379704 392828 379756 392834
rect 379704 392770 379756 392776
rect 379888 392828 379940 392834
rect 379888 392770 379940 392776
rect 379992 392766 380020 534511
rect 380070 531448 380126 531457
rect 380070 531383 380126 531392
rect 380084 397474 380112 531383
rect 380162 525056 380218 525065
rect 380162 524991 380218 525000
rect 380176 398410 380204 524991
rect 380254 521792 380310 521801
rect 380254 521727 380310 521736
rect 380164 398404 380216 398410
rect 380164 398346 380216 398352
rect 380084 397446 380204 397474
rect 380072 397384 380124 397390
rect 380072 397326 380124 397332
rect 380084 393106 380112 397326
rect 380176 393446 380204 397446
rect 380268 397390 380296 521727
rect 380346 515536 380402 515545
rect 380346 515471 380402 515480
rect 380256 397384 380308 397390
rect 380256 397326 380308 397332
rect 380256 395412 380308 395418
rect 380256 395354 380308 395360
rect 380164 393440 380216 393446
rect 380164 393382 380216 393388
rect 380268 393380 380296 395354
rect 380360 393310 380388 515471
rect 380438 512544 380494 512553
rect 380438 512479 380494 512488
rect 380452 398546 380480 512479
rect 380530 509552 380586 509561
rect 380530 509487 380586 509496
rect 380440 398540 380492 398546
rect 380440 398482 380492 398488
rect 380440 398404 380492 398410
rect 380440 398346 380492 398352
rect 380452 393990 380480 398346
rect 380440 393984 380492 393990
rect 380440 393926 380492 393932
rect 380348 393304 380400 393310
rect 380348 393246 380400 393252
rect 380544 393174 380572 509487
rect 380622 503024 380678 503033
rect 380622 502959 380678 502968
rect 380636 398682 380664 502959
rect 380624 398676 380676 398682
rect 380624 398618 380676 398624
rect 380624 398540 380676 398546
rect 380624 398482 380676 398488
rect 380636 394126 380664 398482
rect 380624 394120 380676 394126
rect 380624 394062 380676 394068
rect 380532 393168 380584 393174
rect 380532 393110 380584 393116
rect 380072 393100 380124 393106
rect 380072 393042 380124 393048
rect 380728 392766 380756 569055
rect 391204 556300 391256 556306
rect 391204 556242 391256 556248
rect 380806 553480 380862 553489
rect 380806 553415 380862 553424
rect 380820 392766 380848 553415
rect 386420 407244 386472 407250
rect 386420 407186 386472 407192
rect 386432 402966 386460 407186
rect 386420 402960 386472 402966
rect 386420 402902 386472 402908
rect 387248 402960 387300 402966
rect 387248 402902 387300 402908
rect 384856 395276 384908 395282
rect 384856 395218 384908 395224
rect 382648 395004 382700 395010
rect 382648 394946 382700 394952
rect 382660 393380 382688 394946
rect 384868 393380 384896 395218
rect 387260 393380 387288 402902
rect 389456 395208 389508 395214
rect 389456 395150 389508 395156
rect 389468 393380 389496 395150
rect 377048 392686 377352 392714
rect 379980 392760 380032 392766
rect 379980 392702 380032 392708
rect 380716 392760 380768 392766
rect 380716 392702 380768 392708
rect 380808 392760 380860 392766
rect 380808 392702 380860 392708
rect 390650 380216 390706 380225
rect 390572 380174 390650 380202
rect 390572 367062 390600 380174
rect 390650 380151 390706 380160
rect 390560 367056 390612 367062
rect 390560 366998 390612 367004
rect 390744 366988 390796 366994
rect 390744 366930 390796 366936
rect 390650 366888 390706 366897
rect 390650 366823 390706 366832
rect 364524 360188 364576 360194
rect 364524 360130 364576 360136
rect 360108 360120 360160 360126
rect 360108 360062 360160 360068
rect 360212 360046 360594 360074
rect 360108 358692 360160 358698
rect 360108 358634 360160 358640
rect 359464 358624 359516 358630
rect 359464 358566 359516 358572
rect 358556 354606 358768 354634
rect 358556 345098 358584 354606
rect 358544 345092 358596 345098
rect 358544 345034 358596 345040
rect 358728 345092 358780 345098
rect 358728 345034 358780 345040
rect 358176 340740 358228 340746
rect 358176 340682 358228 340688
rect 358084 340604 358136 340610
rect 358084 340546 358136 340552
rect 358740 335322 358768 345034
rect 358556 335294 358768 335322
rect 358556 325718 358584 335294
rect 358544 325712 358596 325718
rect 358544 325654 358596 325660
rect 358728 325712 358780 325718
rect 358728 325654 358780 325660
rect 358740 316010 358768 325654
rect 358556 315982 358768 316010
rect 358556 306406 358584 315982
rect 358544 306400 358596 306406
rect 358544 306342 358596 306348
rect 358728 306400 358780 306406
rect 358728 306342 358780 306348
rect 358740 296698 358768 306342
rect 358556 296670 358768 296698
rect 358556 287094 358584 296670
rect 358544 287088 358596 287094
rect 358544 287030 358596 287036
rect 358728 287088 358780 287094
rect 358728 287030 358780 287036
rect 357256 280288 357308 280294
rect 357256 280230 357308 280236
rect 357348 280288 357400 280294
rect 357348 280230 357400 280236
rect 357268 280158 357296 280230
rect 357256 280152 357308 280158
rect 357256 280094 357308 280100
rect 358740 277386 358768 287030
rect 358556 277358 358768 277386
rect 357348 270564 357400 270570
rect 357348 270506 357400 270512
rect 357360 263514 357388 270506
rect 358556 267782 358584 277358
rect 358544 267776 358596 267782
rect 358728 267776 358780 267782
rect 358544 267718 358596 267724
rect 358648 267724 358728 267730
rect 358648 267718 358780 267724
rect 358648 267702 358768 267718
rect 358648 263514 358676 267702
rect 357268 263486 357388 263514
rect 358556 263486 358676 263514
rect 357268 251274 357296 263486
rect 358556 251274 358584 263486
rect 357176 251246 357296 251274
rect 358464 251246 358584 251274
rect 357176 251190 357204 251246
rect 358464 251190 358492 251246
rect 357164 251184 357216 251190
rect 357164 251126 357216 251132
rect 357348 251184 357400 251190
rect 357348 251126 357400 251132
rect 358452 251184 358504 251190
rect 358452 251126 358504 251132
rect 358636 251184 358688 251190
rect 358636 251126 358688 251132
rect 357360 234530 357388 251126
rect 358648 234530 358676 251126
rect 357164 234524 357216 234530
rect 357164 234466 357216 234472
rect 357348 234524 357400 234530
rect 357348 234466 357400 234472
rect 358452 234524 358504 234530
rect 358452 234466 358504 234472
rect 358636 234524 358688 234530
rect 358636 234466 358688 234472
rect 357176 224890 357204 234466
rect 358464 224890 358492 234466
rect 357176 224862 357296 224890
rect 358464 224862 358584 224890
rect 357268 212566 357296 224862
rect 358556 215370 358584 224862
rect 358556 215342 358676 215370
rect 357164 212560 357216 212566
rect 357164 212502 357216 212508
rect 357256 212560 357308 212566
rect 357256 212502 357308 212508
rect 356704 201680 356756 201686
rect 356704 201622 356756 201628
rect 357176 200138 357204 212502
rect 358648 205714 358676 215342
rect 358648 205686 358768 205714
rect 358740 202706 358768 205686
rect 358728 202700 358780 202706
rect 358728 202642 358780 202648
rect 357900 202564 357952 202570
rect 357900 202506 357952 202512
rect 357084 200110 357204 200138
rect 357084 200002 357112 200110
rect 357912 200002 357940 202506
rect 359476 202502 359504 358566
rect 360120 202638 360148 358634
rect 360212 340678 360240 360046
rect 362224 358420 362276 358426
rect 362224 358362 362276 358368
rect 361488 358148 361540 358154
rect 361488 358090 361540 358096
rect 360200 340672 360252 340678
rect 360200 340614 360252 340620
rect 361396 202700 361448 202706
rect 361396 202642 361448 202648
rect 359648 202632 359700 202638
rect 359648 202574 359700 202580
rect 360108 202632 360160 202638
rect 360108 202574 360160 202580
rect 360568 202632 360620 202638
rect 360568 202574 360620 202580
rect 358728 202496 358780 202502
rect 358728 202438 358780 202444
rect 359464 202496 359516 202502
rect 359464 202438 359516 202444
rect 358740 200002 358768 202438
rect 359660 200002 359688 202574
rect 360580 200002 360608 202574
rect 361408 200002 361436 202642
rect 361500 202638 361528 358090
rect 362236 202706 362264 358362
rect 362788 357474 362816 360060
rect 363696 358556 363748 358562
rect 363696 358498 363748 358504
rect 362868 358488 362920 358494
rect 362868 358430 362920 358436
rect 362776 357468 362828 357474
rect 362776 357410 362828 357416
rect 362224 202700 362276 202706
rect 362224 202642 362276 202648
rect 362880 202638 362908 358430
rect 363604 357468 363656 357474
rect 363604 357410 363656 357416
rect 363420 202836 363472 202842
rect 363420 202778 363472 202784
rect 361488 202632 361540 202638
rect 361488 202574 361540 202580
rect 362316 202632 362368 202638
rect 362316 202574 362368 202580
rect 362868 202632 362920 202638
rect 362868 202574 362920 202580
rect 362328 200002 362356 202574
rect 362868 202088 362920 202094
rect 362868 202030 362920 202036
rect 362880 200002 362908 202030
rect 355888 199974 355948 200002
rect 356776 199974 357112 200002
rect 357696 199974 357940 200002
rect 358524 199974 358768 200002
rect 359444 199974 359688 200002
rect 360272 199974 360608 200002
rect 361192 199974 361436 200002
rect 362020 199974 362356 200002
rect 362848 199974 362908 200002
rect 363432 200002 363460 202778
rect 363616 202638 363644 357410
rect 363604 202632 363656 202638
rect 363604 202574 363656 202580
rect 363708 202094 363736 358498
rect 364536 222154 364564 360130
rect 365720 360120 365772 360126
rect 365720 360062 365772 360068
rect 364996 358222 365024 360060
rect 364984 358216 365036 358222
rect 364984 358158 365036 358164
rect 364524 222148 364576 222154
rect 364524 222090 364576 222096
rect 364708 212560 364760 212566
rect 364708 212502 364760 212508
rect 364340 202632 364392 202638
rect 364340 202574 364392 202580
rect 363696 202088 363748 202094
rect 363696 202030 363748 202036
rect 364352 200002 364380 202574
rect 364720 200002 364748 212502
rect 365732 200002 365760 360062
rect 367388 358698 367416 360060
rect 367376 358692 367428 358698
rect 367376 358634 367428 358640
rect 369596 358630 369624 360060
rect 369584 358624 369636 358630
rect 369584 358566 369636 358572
rect 371988 358290 372016 360060
rect 374196 358562 374224 360060
rect 374184 358556 374236 358562
rect 374184 358498 374236 358504
rect 376588 358358 376616 360060
rect 378796 358494 378824 360060
rect 380912 360046 381202 360074
rect 378784 358488 378836 358494
rect 378784 358430 378836 358436
rect 376576 358352 376628 358358
rect 376576 358294 376628 358300
rect 371976 358284 372028 358290
rect 371976 358226 372028 358232
rect 380912 340814 380940 360046
rect 383396 358426 383424 360060
rect 385052 360046 385802 360074
rect 383384 358420 383436 358426
rect 383384 358362 383436 358368
rect 385052 340882 385080 360046
rect 387996 358086 388024 360060
rect 390388 358154 390416 360060
rect 390376 358148 390428 358154
rect 390376 358090 390428 358096
rect 387984 358080 388036 358086
rect 387984 358022 388036 358028
rect 385040 340876 385092 340882
rect 385040 340818 385092 340824
rect 380900 340808 380952 340814
rect 380900 340750 380952 340756
rect 390560 227044 390612 227050
rect 390560 226986 390612 226992
rect 390572 219434 390600 226986
rect 390560 219428 390612 219434
rect 390560 219370 390612 219376
rect 390560 209840 390612 209846
rect 390560 209782 390612 209788
rect 375748 202836 375800 202842
rect 375748 202778 375800 202784
rect 374460 202768 374512 202774
rect 374460 202710 374512 202716
rect 367008 202632 367060 202638
rect 367008 202574 367060 202580
rect 367020 200002 367048 202574
rect 374472 200002 374500 202710
rect 375760 200002 375788 202778
rect 376484 202700 376536 202706
rect 376484 202642 376536 202648
rect 376496 200002 376524 202642
rect 390572 202298 390600 209782
rect 390664 202434 390692 366823
rect 390756 357406 390784 366930
rect 390744 357400 390796 357406
rect 390744 357342 390796 357348
rect 390928 357400 390980 357406
rect 390928 357342 390980 357348
rect 390940 356046 390968 357342
rect 390928 356040 390980 356046
rect 390928 355982 390980 355988
rect 390928 346452 390980 346458
rect 390928 346394 390980 346400
rect 390940 340950 390968 346394
rect 390928 340944 390980 340950
rect 390928 340886 390980 340892
rect 390836 340876 390888 340882
rect 390836 340818 390888 340824
rect 390848 338178 390876 340818
rect 390848 338150 390968 338178
rect 390940 336734 390968 338150
rect 390928 336728 390980 336734
rect 390928 336670 390980 336676
rect 390928 327140 390980 327146
rect 390928 327082 390980 327088
rect 390940 321706 390968 327082
rect 390928 321700 390980 321706
rect 390928 321642 390980 321648
rect 390836 321564 390888 321570
rect 390836 321506 390888 321512
rect 390848 318730 390876 321506
rect 390926 318744 390982 318753
rect 390848 318702 390926 318730
rect 390926 318679 390982 318688
rect 390926 309224 390982 309233
rect 390926 309159 390982 309168
rect 390940 309126 390968 309159
rect 390928 309120 390980 309126
rect 390928 309062 390980 309068
rect 390836 299532 390888 299538
rect 390836 299474 390888 299480
rect 390848 299418 390876 299474
rect 390926 299432 390982 299441
rect 390848 299390 390926 299418
rect 390926 299367 390982 299376
rect 390926 289912 390982 289921
rect 390926 289847 390982 289856
rect 390940 289814 390968 289847
rect 390928 289808 390980 289814
rect 390928 289750 390980 289756
rect 390836 280220 390888 280226
rect 390836 280162 390888 280168
rect 390848 280106 390876 280162
rect 390926 280120 390982 280129
rect 390848 280078 390926 280106
rect 390926 280055 390982 280064
rect 390926 270600 390982 270609
rect 390926 270535 390982 270544
rect 390940 270502 390968 270535
rect 390928 270496 390980 270502
rect 390928 270438 390980 270444
rect 390928 263492 390980 263498
rect 390928 263434 390980 263440
rect 390940 260846 390968 263434
rect 390928 260840 390980 260846
rect 390928 260782 390980 260788
rect 390928 253836 390980 253842
rect 390928 253778 390980 253784
rect 390940 251190 390968 253778
rect 390928 251184 390980 251190
rect 390928 251126 390980 251132
rect 391020 241528 391072 241534
rect 391020 241470 391072 241476
rect 391032 231878 391060 241470
rect 390836 231872 390888 231878
rect 390836 231814 390888 231820
rect 391020 231872 391072 231878
rect 391020 231814 391072 231820
rect 390848 227050 390876 231814
rect 390836 227044 390888 227050
rect 390836 226986 390888 226992
rect 390744 219428 390796 219434
rect 390744 219370 390796 219376
rect 390756 209846 390784 219370
rect 390744 209840 390796 209846
rect 390744 209782 390796 209788
rect 391216 202842 391244 556242
rect 395344 556232 395396 556238
rect 395344 556174 395396 556180
rect 391296 518288 391348 518294
rect 391296 518230 391348 518236
rect 391204 202836 391256 202842
rect 391204 202778 391256 202784
rect 391308 202774 391336 518230
rect 393320 407788 393372 407794
rect 393320 407730 393372 407736
rect 391938 387560 391994 387569
rect 391938 387495 391994 387504
rect 391296 202768 391348 202774
rect 391296 202710 391348 202716
rect 390652 202428 390704 202434
rect 390652 202370 390704 202376
rect 390560 202292 390612 202298
rect 390560 202234 390612 202240
rect 391952 202230 391980 387495
rect 393332 384033 393360 407730
rect 393412 406496 393464 406502
rect 393412 406438 393464 406444
rect 393424 390833 393452 406438
rect 393410 390824 393466 390833
rect 393410 390759 393466 390768
rect 393318 384024 393374 384033
rect 393318 383959 393374 383968
rect 393318 377224 393374 377233
rect 393318 377159 393374 377168
rect 392030 370424 392086 370433
rect 392030 370359 392086 370368
rect 392044 202366 392072 370359
rect 393332 202570 393360 377159
rect 393410 373960 393466 373969
rect 393410 373895 393466 373904
rect 393320 202564 393372 202570
rect 393320 202506 393372 202512
rect 392032 202360 392084 202366
rect 392032 202302 392084 202308
rect 391940 202224 391992 202230
rect 391940 202166 391992 202172
rect 393424 202162 393452 373895
rect 393502 363624 393558 363633
rect 393502 363559 393558 363568
rect 393516 202502 393544 363559
rect 395356 202638 395384 556174
rect 398104 518220 398156 518226
rect 398104 518162 398156 518168
rect 398116 202706 398144 518162
rect 416596 389428 416648 389434
rect 416596 389370 416648 389376
rect 401508 389292 401560 389298
rect 401508 389234 401560 389240
rect 401416 337612 401468 337618
rect 401416 337554 401468 337560
rect 401428 202842 401456 337554
rect 400588 202836 400640 202842
rect 400588 202778 400640 202784
rect 401416 202836 401468 202842
rect 401416 202778 401468 202784
rect 398104 202700 398156 202706
rect 398104 202642 398156 202648
rect 395344 202632 395396 202638
rect 395344 202574 395396 202580
rect 393504 202496 393556 202502
rect 393504 202438 393556 202444
rect 393412 202156 393464 202162
rect 393412 202098 393464 202104
rect 400600 200002 400628 202778
rect 401520 202434 401548 389234
rect 413928 374060 413980 374066
rect 413928 374002 413980 374008
rect 412548 357468 412600 357474
rect 412548 357410 412600 357416
rect 411168 337544 411220 337550
rect 411168 337486 411220 337492
rect 408408 337476 408460 337482
rect 408408 337418 408460 337424
rect 400956 202428 401008 202434
rect 400956 202370 401008 202376
rect 401508 202428 401560 202434
rect 401508 202370 401560 202376
rect 400968 200002 400996 202370
rect 408420 200002 408448 337418
rect 411076 202224 411128 202230
rect 411076 202166 411128 202172
rect 409236 202156 409288 202162
rect 409236 202098 409288 202104
rect 409248 200002 409276 202098
rect 410156 201544 410208 201550
rect 410156 201486 410208 201492
rect 410168 200002 410196 201486
rect 363432 199974 363768 200002
rect 364352 199974 364596 200002
rect 364720 199974 365056 200002
rect 365732 199974 365976 200002
rect 366804 199974 367048 200002
rect 374164 199974 374500 200002
rect 375452 199974 375788 200002
rect 376372 199974 376524 200002
rect 400292 199974 400628 200002
rect 400752 199974 400996 200002
rect 408112 199974 408448 200002
rect 408940 199974 409276 200002
rect 409860 199974 410196 200002
rect 411088 200002 411116 202166
rect 411180 201550 411208 337486
rect 411168 201544 411220 201550
rect 411168 201486 411220 201492
rect 412560 200138 412588 357410
rect 413836 337408 413888 337414
rect 413836 337350 413888 337356
rect 413192 202836 413244 202842
rect 413192 202778 413244 202784
rect 412284 200110 412588 200138
rect 412284 200002 412312 200110
rect 413204 200002 413232 202778
rect 413848 200002 413876 337350
rect 413940 202842 413968 374002
rect 416608 202842 416636 389370
rect 418068 389360 418120 389366
rect 418068 389302 418120 389308
rect 416688 389224 416740 389230
rect 416688 389166 416740 389172
rect 413928 202836 413980 202842
rect 413928 202778 413980 202784
rect 415768 202836 415820 202842
rect 415768 202778 415820 202784
rect 416596 202836 416648 202842
rect 416596 202778 416648 202784
rect 414940 202292 414992 202298
rect 414940 202234 414992 202240
rect 414952 200002 414980 202234
rect 415780 200002 415808 202778
rect 416700 202722 416728 389166
rect 418080 202842 418108 389302
rect 417516 202836 417568 202842
rect 417516 202778 417568 202784
rect 418068 202836 418120 202842
rect 418068 202778 418120 202784
rect 416608 202694 416728 202722
rect 416608 200002 416636 202694
rect 417528 200002 417556 202778
rect 411088 199974 411148 200002
rect 411976 199974 412312 200002
rect 412896 199974 413232 200002
rect 413724 199974 413876 200002
rect 414644 199974 414980 200002
rect 415472 199974 415808 200002
rect 416392 199974 416636 200002
rect 417220 199974 417556 200002
rect 238760 199912 238812 199918
rect 238760 199854 238812 199860
rect 239496 199912 239548 199918
rect 243084 199912 243136 199918
rect 239548 199860 239844 199866
rect 239496 199854 239844 199860
rect 243084 199854 243136 199860
rect 243820 199912 243872 199918
rect 243872 199860 244168 199866
rect 243820 199854 244168 199860
rect 239508 199838 239844 199854
rect 243832 199838 244168 199854
rect 134064 195968 134116 195974
rect 134064 195910 134116 195916
rect 133878 180367 133934 180376
rect 133972 180396 134024 180402
rect 133972 180338 134024 180344
rect 134076 180282 134104 195910
rect 133892 180254 134104 180282
rect 133892 176662 133920 180254
rect 133880 176656 133932 176662
rect 133880 176598 133932 176604
rect 134064 176656 134116 176662
rect 134064 176598 134116 176604
rect 133972 172576 134024 172582
rect 133972 172518 134024 172524
rect 133984 162858 134012 172518
rect 133972 162852 134024 162858
rect 133972 162794 134024 162800
rect 133972 143608 134024 143614
rect 133972 143550 134024 143556
rect 133984 143426 134012 143550
rect 133892 143398 134012 143426
rect 133786 140448 133842 140457
rect 133786 140383 133842 140392
rect 133892 138718 133920 143398
rect 133880 138712 133932 138718
rect 133880 138654 133932 138660
rect 133880 125656 133932 125662
rect 133880 125598 133932 125604
rect 133892 122074 133920 125598
rect 133970 123040 134026 123049
rect 133970 122975 134026 122984
rect 133708 122046 133920 122074
rect 133708 120986 133736 122046
rect 133878 121952 133934 121961
rect 133878 121887 133934 121896
rect 133892 121242 133920 121887
rect 133880 121236 133932 121242
rect 133880 121178 133932 121184
rect 133984 121106 134012 122975
rect 133972 121100 134024 121106
rect 133972 121042 134024 121048
rect 133708 120958 133920 120986
rect 134076 120970 134104 176598
rect 433904 157321 433932 699654
rect 433996 159361 434024 700674
rect 434088 161265 434116 700878
rect 434168 700800 434220 700806
rect 434168 700742 434220 700748
rect 434180 163577 434208 700742
rect 434352 700664 434404 700670
rect 434352 700606 434404 700612
rect 434260 700324 434312 700330
rect 434260 700266 434312 700272
rect 434272 169697 434300 700266
rect 434258 169688 434314 169697
rect 434258 169623 434314 169632
rect 434364 165617 434392 700606
rect 434444 700460 434496 700466
rect 434444 700402 434496 700408
rect 438124 700460 438176 700466
rect 438124 700402 438176 700408
rect 434456 167793 434484 700402
rect 434720 681760 434772 681766
rect 434720 681702 434772 681708
rect 434536 294024 434588 294030
rect 434536 293966 434588 293972
rect 434548 186289 434576 293966
rect 434534 186280 434590 186289
rect 434534 186215 434590 186224
rect 434732 172009 434760 681702
rect 434812 623824 434864 623830
rect 434812 623766 434864 623772
rect 434824 173913 434852 623766
rect 436744 438932 436796 438938
rect 436744 438874 436796 438880
rect 436100 355360 436152 355366
rect 436100 355302 436152 355308
rect 434904 336796 434956 336802
rect 434904 336738 434956 336744
rect 434916 184657 434944 336738
rect 435088 251252 435140 251258
rect 435088 251194 435140 251200
rect 434994 196208 435050 196217
rect 434994 196143 435050 196152
rect 434902 184648 434958 184657
rect 434902 184583 434958 184592
rect 434810 173904 434866 173913
rect 434810 173839 434866 173848
rect 434718 172000 434774 172009
rect 434718 171935 434774 171944
rect 434442 167784 434498 167793
rect 434442 167719 434498 167728
rect 434350 165608 434406 165617
rect 434350 165543 434406 165552
rect 434166 163568 434222 163577
rect 434166 163503 434222 163512
rect 434074 161256 434130 161265
rect 434074 161191 434130 161200
rect 433982 159352 434038 159361
rect 433982 159287 434038 159296
rect 433890 157312 433946 157321
rect 433890 157247 433946 157256
rect 133892 118153 133920 120958
rect 134064 120964 134116 120970
rect 134064 120906 134116 120912
rect 388332 120278 388760 120306
rect 164988 120142 165508 120170
rect 200500 120142 201020 120170
rect 202860 120142 203104 120170
rect 134168 120006 134320 120034
rect 134536 120006 134872 120034
rect 135364 120006 135516 120034
rect 135732 120006 136068 120034
rect 133878 118144 133934 118153
rect 133878 118079 133934 118088
rect 133880 113892 133932 113898
rect 133880 113834 133932 113840
rect 133248 38622 133276 41398
rect 133604 41404 133656 41410
rect 133604 41346 133656 41352
rect 133236 38616 133288 38622
rect 133236 38558 133288 38564
rect 133144 31068 133196 31074
rect 133144 31010 133196 31016
rect 132408 30320 132460 30326
rect 132408 30262 132460 30268
rect 133156 22114 133184 31010
rect 132224 22092 132276 22098
rect 133156 22086 133276 22114
rect 132224 22034 132276 22040
rect 133248 12458 133276 22086
rect 133064 12430 133276 12458
rect 131764 8288 131816 8294
rect 131764 8230 131816 8236
rect 131396 7200 131448 7206
rect 131396 7142 131448 7148
rect 130384 4480 130436 4486
rect 130384 4422 130436 4428
rect 131408 480 131436 7142
rect 133064 7138 133092 12430
rect 133788 8288 133840 8294
rect 133788 8230 133840 8236
rect 133052 7132 133104 7138
rect 133052 7074 133104 7080
rect 133144 7132 133196 7138
rect 133144 7074 133196 7080
rect 133156 3330 133184 7074
rect 132592 3324 132644 3330
rect 132592 3266 132644 3272
rect 133144 3324 133196 3330
rect 133144 3266 133196 3272
rect 132604 480 132632 3266
rect 133800 480 133828 8230
rect 133892 7818 133920 113834
rect 133880 7812 133932 7818
rect 133880 7754 133932 7760
rect 134168 7614 134196 120006
rect 134536 113898 134564 120006
rect 134524 113892 134576 113898
rect 134524 113834 134576 113840
rect 135260 113892 135312 113898
rect 135260 113834 135312 113840
rect 134156 7608 134208 7614
rect 134156 7550 134208 7556
rect 134892 7608 134944 7614
rect 134892 7550 134944 7556
rect 134904 480 134932 7550
rect 135272 4826 135300 113834
rect 135364 7682 135392 120006
rect 135444 117496 135496 117502
rect 135444 117438 135496 117444
rect 135352 7676 135404 7682
rect 135352 7618 135404 7624
rect 135456 5098 135484 117438
rect 135732 113898 135760 120006
rect 136698 119762 136726 120020
rect 136652 119734 136726 119762
rect 136836 120006 137356 120034
rect 137572 120006 137908 120034
rect 138216 120006 138552 120034
rect 138860 120006 139196 120034
rect 139596 120006 139748 120034
rect 140056 120006 140392 120034
rect 140792 120006 141036 120034
rect 141252 120006 141588 120034
rect 142232 120006 142384 120034
rect 135720 113892 135772 113898
rect 135720 113834 135772 113840
rect 136088 7812 136140 7818
rect 136088 7754 136140 7760
rect 135444 5092 135496 5098
rect 135444 5034 135496 5040
rect 135260 4820 135312 4826
rect 135260 4762 135312 4768
rect 136100 480 136128 7754
rect 136652 7750 136680 119734
rect 136732 113892 136784 113898
rect 136732 113834 136784 113840
rect 136744 7886 136772 113834
rect 136836 8974 136864 120006
rect 137572 113898 137600 120006
rect 138216 117473 138244 120006
rect 138860 119406 138888 120006
rect 138296 119400 138348 119406
rect 138296 119342 138348 119348
rect 138848 119400 138900 119406
rect 138848 119342 138900 119348
rect 138202 117464 138258 117473
rect 138202 117399 138258 117408
rect 137560 113892 137612 113898
rect 138308 113880 138336 119342
rect 137560 113834 137612 113840
rect 138124 113852 138336 113880
rect 139492 113892 139544 113898
rect 138124 101402 138152 113852
rect 139492 113834 139544 113840
rect 137940 101374 138152 101402
rect 137940 96665 137968 101374
rect 137926 96656 137982 96665
rect 137926 96591 137982 96600
rect 138202 96656 138258 96665
rect 138202 96591 138258 96600
rect 138216 12458 138244 96591
rect 138032 12430 138244 12458
rect 136824 8968 136876 8974
rect 136824 8910 136876 8916
rect 136732 7880 136784 7886
rect 136732 7822 136784 7828
rect 136640 7744 136692 7750
rect 136640 7686 136692 7692
rect 137284 7676 137336 7682
rect 137284 7618 137336 7624
rect 137296 480 137324 7618
rect 138032 3534 138060 12430
rect 138480 5092 138532 5098
rect 138480 5034 138532 5040
rect 138020 3528 138072 3534
rect 138020 3470 138072 3476
rect 138492 480 138520 5034
rect 139504 4894 139532 113834
rect 139492 4888 139544 4894
rect 139492 4830 139544 4836
rect 139596 3466 139624 120006
rect 140056 113898 140084 120006
rect 140792 118697 140820 120006
rect 140778 118688 140834 118697
rect 140778 118623 140834 118632
rect 140792 117337 140820 118623
rect 140778 117328 140834 117337
rect 140778 117263 140834 117272
rect 140962 117328 141018 117337
rect 140962 117263 141018 117272
rect 140044 113892 140096 113898
rect 140044 113834 140096 113840
rect 140780 113892 140832 113898
rect 140780 113834 140832 113840
rect 139676 7744 139728 7750
rect 139676 7686 139728 7692
rect 139584 3460 139636 3466
rect 139584 3402 139636 3408
rect 139688 480 139716 7686
rect 140792 3670 140820 113834
rect 140976 113778 141004 117263
rect 141252 113898 141280 120006
rect 142252 118924 142304 118930
rect 142252 118866 142304 118872
rect 142160 117972 142212 117978
rect 142160 117914 142212 117920
rect 141884 117496 141936 117502
rect 142172 117450 142200 117914
rect 141936 117444 142200 117450
rect 141884 117438 142200 117444
rect 141896 117422 142200 117438
rect 141240 113892 141292 113898
rect 141240 113834 141292 113840
rect 140884 113750 141004 113778
rect 140884 7954 140912 113750
rect 140872 7948 140924 7954
rect 140872 7890 140924 7896
rect 140964 7880 141016 7886
rect 140964 7822 141016 7828
rect 140780 3664 140832 3670
rect 140780 3606 140832 3612
rect 140976 2802 141004 7822
rect 142264 4962 142292 118866
rect 142252 4956 142304 4962
rect 142252 4898 142304 4904
rect 142068 4820 142120 4826
rect 142068 4762 142120 4768
rect 140884 2774 141004 2802
rect 140884 480 140912 2774
rect 142080 480 142108 4762
rect 142356 3602 142384 120006
rect 142540 120006 142876 120034
rect 143092 120006 143428 120034
rect 143552 120006 144072 120034
rect 144380 120006 144716 120034
rect 145116 120006 145268 120034
rect 145576 120006 145912 120034
rect 146404 120006 146556 120034
rect 146772 120006 147108 120034
rect 142540 118930 142568 120006
rect 142528 118924 142580 118930
rect 142528 118866 142580 118872
rect 142802 118688 142858 118697
rect 142802 118623 142858 118632
rect 142816 118153 142844 118623
rect 142802 118144 142858 118153
rect 142802 118079 142858 118088
rect 143092 117978 143120 120006
rect 143080 117972 143132 117978
rect 143080 117914 143132 117920
rect 143264 7948 143316 7954
rect 143264 7890 143316 7896
rect 142344 3596 142396 3602
rect 142344 3538 142396 3544
rect 143276 480 143304 7890
rect 143552 3738 143580 120006
rect 144380 119406 144408 120006
rect 143632 119400 143684 119406
rect 143632 119342 143684 119348
rect 144368 119400 144420 119406
rect 144368 119342 144420 119348
rect 143644 19310 143672 119342
rect 145116 118862 145144 120006
rect 145104 118856 145156 118862
rect 145104 118798 145156 118804
rect 145116 95402 145144 118798
rect 145576 117881 145604 120006
rect 145562 117872 145618 117881
rect 145562 117807 145618 117816
rect 146300 113892 146352 113898
rect 146300 113834 146352 113840
rect 145104 95396 145156 95402
rect 145104 95338 145156 95344
rect 145104 95260 145156 95266
rect 145104 95202 145156 95208
rect 145116 90438 145144 95202
rect 145104 90432 145156 90438
rect 145104 90374 145156 90380
rect 144920 85604 144972 85610
rect 144920 85546 144972 85552
rect 144932 80730 144960 85546
rect 144932 80702 145328 80730
rect 145300 66366 145328 80702
rect 145104 66360 145156 66366
rect 145104 66302 145156 66308
rect 145288 66360 145340 66366
rect 145288 66302 145340 66308
rect 145116 64870 145144 66302
rect 145104 64864 145156 64870
rect 145104 64806 145156 64812
rect 145104 56568 145156 56574
rect 145104 56510 145156 56516
rect 145116 37210 145144 56510
rect 145116 37182 145236 37210
rect 145208 31822 145236 37182
rect 145012 31816 145064 31822
rect 145012 31758 145064 31764
rect 145196 31816 145248 31822
rect 145196 31758 145248 31764
rect 145024 24154 145052 31758
rect 145024 24126 145144 24154
rect 143632 19304 143684 19310
rect 143632 19246 143684 19252
rect 143724 9716 143776 9722
rect 143724 9658 143776 9664
rect 143736 8022 143764 9658
rect 143724 8016 143776 8022
rect 143724 7958 143776 7964
rect 144460 8016 144512 8022
rect 144460 7958 144512 7964
rect 143540 3732 143592 3738
rect 143540 3674 143592 3680
rect 144472 480 144500 7958
rect 145116 5030 145144 24126
rect 145104 5024 145156 5030
rect 145104 4966 145156 4972
rect 145656 4888 145708 4894
rect 145656 4830 145708 4836
rect 145668 480 145696 4830
rect 146312 3874 146340 113834
rect 146300 3868 146352 3874
rect 146300 3810 146352 3816
rect 146404 3806 146432 120006
rect 146772 113898 146800 120006
rect 147738 119762 147766 120020
rect 148060 120006 148396 120034
rect 148520 120006 148948 120034
rect 149072 120006 149592 120034
rect 149900 120006 150236 120034
rect 150452 120006 150788 120034
rect 151188 120006 151432 120034
rect 151832 120006 151984 120034
rect 152108 120006 152628 120034
rect 147738 119734 147812 119762
rect 147784 118794 147812 119734
rect 147772 118788 147824 118794
rect 147772 118730 147824 118736
rect 146760 113892 146812 113898
rect 146760 113834 146812 113840
rect 147784 9042 147812 118730
rect 148060 117434 148088 120006
rect 148048 117428 148100 117434
rect 148048 117370 148100 117376
rect 148520 104922 148548 120006
rect 149072 118726 149100 120006
rect 149060 118720 149112 118726
rect 149060 118662 149112 118668
rect 148232 104916 148284 104922
rect 148232 104858 148284 104864
rect 148508 104916 148560 104922
rect 148508 104858 148560 104864
rect 148244 95266 148272 104858
rect 147956 95260 148008 95266
rect 147956 95202 148008 95208
rect 148232 95260 148284 95266
rect 148232 95202 148284 95208
rect 147968 90386 147996 95202
rect 147968 90358 148088 90386
rect 148060 66473 148088 90358
rect 148046 66464 148102 66473
rect 148046 66399 148102 66408
rect 147954 66328 148010 66337
rect 147954 66263 148010 66272
rect 147968 64870 147996 66263
rect 147956 64864 148008 64870
rect 147956 64806 148008 64812
rect 147956 55276 148008 55282
rect 147956 55218 148008 55224
rect 147968 51814 147996 55218
rect 147956 51808 148008 51814
rect 147956 51750 148008 51756
rect 148140 51808 148192 51814
rect 148140 51750 148192 51756
rect 148152 42090 148180 51750
rect 147864 42084 147916 42090
rect 147864 42026 147916 42032
rect 148140 42084 148192 42090
rect 148140 42026 148192 42032
rect 147876 24206 147904 42026
rect 147864 24200 147916 24206
rect 147864 24142 147916 24148
rect 148048 24200 148100 24206
rect 148048 24142 148100 24148
rect 147772 9036 147824 9042
rect 147772 8978 147824 8984
rect 148060 6186 148088 24142
rect 148048 6180 148100 6186
rect 148048 6122 148100 6128
rect 149072 4865 149100 118662
rect 149900 118386 149928 120006
rect 149888 118380 149940 118386
rect 149888 118322 149940 118328
rect 149244 4956 149296 4962
rect 149244 4898 149296 4904
rect 149058 4856 149114 4865
rect 149058 4791 149114 4800
rect 146392 3800 146444 3806
rect 146392 3742 146444 3748
rect 148048 3664 148100 3670
rect 148048 3606 148100 3612
rect 146852 2848 146904 2854
rect 146852 2790 146904 2796
rect 146864 480 146892 2790
rect 148060 480 148088 3606
rect 149256 480 149284 4898
rect 150452 3942 150480 120006
rect 151188 114578 151216 120006
rect 151832 117745 151860 120006
rect 151818 117736 151874 117745
rect 152108 117688 152136 120006
rect 153258 119762 153286 120020
rect 153488 120006 153824 120034
rect 154132 120006 154468 120034
rect 154684 120006 155112 120034
rect 155328 120006 155664 120034
rect 155972 120006 156308 120034
rect 153258 119734 153332 119762
rect 151818 117671 151874 117680
rect 151924 117660 152136 117688
rect 150900 114572 150952 114578
rect 150900 114514 150952 114520
rect 151176 114572 151228 114578
rect 151176 114514 151228 114520
rect 150912 109018 150940 114514
rect 151924 113914 151952 117660
rect 152004 117564 152056 117570
rect 152004 117506 152056 117512
rect 150728 108990 150940 109018
rect 151832 113886 151952 113914
rect 150728 99482 150756 108990
rect 150716 99476 150768 99482
rect 150716 99418 150768 99424
rect 150624 99340 150676 99346
rect 150624 99282 150676 99288
rect 150636 85678 150664 99282
rect 150624 85672 150676 85678
rect 150624 85614 150676 85620
rect 150532 85604 150584 85610
rect 150532 85546 150584 85552
rect 150544 80782 150572 85546
rect 150532 80776 150584 80782
rect 150532 80718 150584 80724
rect 150716 80776 150768 80782
rect 150716 80718 150768 80724
rect 150728 70514 150756 80718
rect 150716 70508 150768 70514
rect 150716 70450 150768 70456
rect 150624 70372 150676 70378
rect 150624 70314 150676 70320
rect 150636 60738 150664 70314
rect 150544 60722 150664 60738
rect 150532 60716 150664 60722
rect 150584 60710 150664 60716
rect 150716 60716 150768 60722
rect 150532 60658 150584 60664
rect 150716 60658 150768 60664
rect 150728 57934 150756 60658
rect 150716 57928 150768 57934
rect 150716 57870 150768 57876
rect 150808 48340 150860 48346
rect 150808 48282 150860 48288
rect 150820 41478 150848 48282
rect 150808 41472 150860 41478
rect 150808 41414 150860 41420
rect 150808 38616 150860 38622
rect 150808 38558 150860 38564
rect 150820 37262 150848 38558
rect 150808 37256 150860 37262
rect 150808 37198 150860 37204
rect 150716 27668 150768 27674
rect 150716 27610 150768 27616
rect 150728 5166 150756 27610
rect 151832 6254 151860 113886
rect 152016 113778 152044 117506
rect 153200 113892 153252 113898
rect 153200 113834 153252 113840
rect 151924 113750 152044 113778
rect 151820 6248 151872 6254
rect 151820 6190 151872 6196
rect 150716 5160 150768 5166
rect 150716 5102 150768 5108
rect 151924 4146 151952 113750
rect 152740 5024 152792 5030
rect 152740 4966 152792 4972
rect 151912 4140 151964 4146
rect 151912 4082 151964 4088
rect 150440 3936 150492 3942
rect 150440 3878 150492 3884
rect 151544 3800 151596 3806
rect 151544 3742 151596 3748
rect 150440 2916 150492 2922
rect 150440 2858 150492 2864
rect 150452 480 150480 2858
rect 151556 480 151584 3742
rect 152752 480 152780 4966
rect 153212 4010 153240 113834
rect 153304 5234 153332 119734
rect 153488 118017 153516 120006
rect 153474 118008 153530 118017
rect 153474 117943 153530 117952
rect 154132 113898 154160 120006
rect 154120 113892 154172 113898
rect 154120 113834 154172 113840
rect 154684 9110 154712 120006
rect 155328 117570 155356 120006
rect 155316 117564 155368 117570
rect 155316 117506 155368 117512
rect 154672 9104 154724 9110
rect 154672 9046 154724 9052
rect 153936 6180 153988 6186
rect 153936 6122 153988 6128
rect 153292 5228 153344 5234
rect 153292 5170 153344 5176
rect 153200 4004 153252 4010
rect 153200 3946 153252 3952
rect 153948 480 153976 6122
rect 155132 5160 155184 5166
rect 155132 5102 155184 5108
rect 155144 480 155172 5102
rect 155972 4078 156000 120006
rect 156938 119762 156966 120020
rect 156892 119734 156966 119762
rect 157352 120006 157504 120034
rect 157812 120006 158148 120034
rect 156892 117978 156920 119734
rect 157246 118688 157302 118697
rect 157246 118623 157302 118632
rect 157260 118153 157288 118623
rect 157246 118144 157302 118153
rect 157246 118079 157302 118088
rect 156512 117972 156564 117978
rect 156512 117914 156564 117920
rect 156880 117972 156932 117978
rect 156880 117914 156932 117920
rect 156524 109018 156552 117914
rect 157352 117706 157380 120006
rect 157340 117700 157392 117706
rect 157340 117642 157392 117648
rect 157812 114578 157840 120006
rect 158778 119762 158806 120020
rect 159008 120006 159344 120034
rect 159652 120006 159988 120034
rect 160204 120006 160632 120034
rect 160848 120006 161184 120034
rect 161584 120006 161828 120034
rect 162136 120006 162472 120034
rect 162872 120006 163024 120034
rect 163424 120006 163668 120034
rect 158778 119734 158852 119762
rect 157432 114572 157484 114578
rect 157432 114514 157484 114520
rect 157800 114572 157852 114578
rect 157800 114514 157852 114520
rect 156156 108990 156552 109018
rect 156156 100042 156184 108990
rect 157444 103562 157472 114514
rect 157248 103556 157300 103562
rect 157248 103498 157300 103504
rect 157432 103556 157484 103562
rect 157432 103498 157484 103504
rect 156064 100014 156184 100042
rect 156064 93838 156092 100014
rect 156052 93832 156104 93838
rect 156052 93774 156104 93780
rect 157260 90386 157288 103498
rect 157260 90358 157472 90386
rect 156144 84244 156196 84250
rect 156144 84186 156196 84192
rect 156156 84130 156184 84186
rect 156064 84102 156184 84130
rect 156064 74594 156092 84102
rect 157444 75886 157472 90358
rect 157432 75880 157484 75886
rect 157432 75822 157484 75828
rect 156052 74588 156104 74594
rect 156052 74530 156104 74536
rect 156236 74588 156288 74594
rect 156236 74530 156288 74536
rect 156248 70394 156276 74530
rect 156156 70366 156276 70394
rect 156156 60738 156184 70366
rect 157432 66292 157484 66298
rect 157432 66234 157484 66240
rect 156064 60722 156184 60738
rect 156052 60716 156184 60722
rect 156104 60710 156184 60716
rect 156236 60716 156288 60722
rect 156052 60658 156104 60664
rect 156236 60658 156288 60664
rect 156248 51762 156276 60658
rect 156064 51734 156276 51762
rect 156064 48226 156092 51734
rect 156064 48198 156184 48226
rect 156156 46866 156184 48198
rect 157444 46918 157472 66234
rect 156064 46838 156184 46866
rect 157432 46912 157484 46918
rect 157432 46854 157484 46860
rect 156064 38570 156092 46838
rect 156064 38542 156368 38570
rect 156340 27554 156368 38542
rect 157340 37324 157392 37330
rect 157340 37266 157392 37272
rect 157352 29034 157380 37266
rect 157340 29028 157392 29034
rect 157340 28970 157392 28976
rect 157432 29028 157484 29034
rect 157432 28970 157484 28976
rect 157444 27606 157472 28970
rect 157432 27600 157484 27606
rect 156340 27526 156460 27554
rect 157432 27542 157484 27548
rect 156432 22794 156460 27526
rect 156248 22766 156460 22794
rect 156248 5302 156276 22766
rect 157340 9716 157392 9722
rect 157340 9658 157392 9664
rect 157352 9178 157380 9658
rect 157340 9172 157392 9178
rect 157340 9114 157392 9120
rect 158824 8090 158852 119734
rect 159008 117638 159036 120006
rect 158996 117632 159048 117638
rect 158996 117574 159048 117580
rect 159652 115977 159680 120006
rect 159086 115968 159142 115977
rect 159086 115903 159142 115912
rect 159638 115968 159694 115977
rect 159638 115903 159694 115912
rect 159100 100042 159128 115903
rect 159100 100014 159220 100042
rect 159192 77466 159220 100014
rect 159100 77438 159220 77466
rect 159100 64870 159128 77438
rect 159088 64864 159140 64870
rect 159088 64806 159140 64812
rect 159088 55276 159140 55282
rect 159088 55218 159140 55224
rect 159100 51134 159128 55218
rect 159088 51128 159140 51134
rect 159088 51070 159140 51076
rect 159088 50992 159140 50998
rect 159088 50934 159140 50940
rect 159100 29034 159128 50934
rect 159088 29028 159140 29034
rect 159088 28970 159140 28976
rect 159272 29028 159324 29034
rect 159272 28970 159324 28976
rect 159284 19378 159312 28970
rect 159088 19372 159140 19378
rect 159088 19314 159140 19320
rect 159272 19372 159324 19378
rect 159272 19314 159324 19320
rect 158812 8084 158864 8090
rect 158812 8026 158864 8032
rect 156236 5296 156288 5302
rect 156236 5238 156288 5244
rect 158720 5296 158772 5302
rect 158720 5238 158772 5244
rect 156328 5228 156380 5234
rect 156328 5170 156380 5176
rect 155960 4072 156012 4078
rect 155960 4014 156012 4020
rect 156340 480 156368 5170
rect 157524 3868 157576 3874
rect 157524 3810 157576 3816
rect 157536 480 157564 3810
rect 158732 480 158760 5238
rect 159100 3398 159128 19314
rect 160204 8158 160232 120006
rect 160848 117910 160876 120006
rect 160836 117904 160888 117910
rect 160836 117846 160888 117852
rect 161480 113892 161532 113898
rect 161480 113834 161532 113840
rect 161492 9382 161520 113834
rect 161480 9376 161532 9382
rect 161480 9318 161532 9324
rect 161584 9246 161612 120006
rect 162136 113898 162164 120006
rect 162872 117842 162900 120006
rect 162860 117836 162912 117842
rect 162860 117778 162912 117784
rect 163424 115977 163452 120006
rect 164298 119762 164326 120020
rect 164528 120006 164864 120034
rect 164298 119734 164372 119762
rect 163042 115968 163098 115977
rect 163042 115903 163098 115912
rect 163410 115968 163466 115977
rect 163410 115903 163466 115912
rect 162124 113892 162176 113898
rect 162124 113834 162176 113840
rect 163056 93906 163084 115903
rect 162860 93900 162912 93906
rect 162860 93842 162912 93848
rect 163044 93900 163096 93906
rect 163044 93842 163096 93848
rect 162872 84182 162900 93842
rect 162860 84176 162912 84182
rect 162860 84118 162912 84124
rect 162860 74588 162912 74594
rect 162860 74530 162912 74536
rect 162872 64870 162900 74530
rect 162860 64864 162912 64870
rect 162860 64806 162912 64812
rect 163136 64864 163188 64870
rect 163136 64806 163188 64812
rect 163148 19378 163176 64806
rect 162952 19372 163004 19378
rect 162952 19314 163004 19320
rect 163136 19372 163188 19378
rect 163136 19314 163188 19320
rect 162964 9602 162992 19314
rect 162872 9574 162992 9602
rect 161572 9240 161624 9246
rect 161572 9182 161624 9188
rect 160192 8152 160244 8158
rect 160192 8094 160244 8100
rect 162872 6322 162900 9574
rect 164344 9314 164372 119734
rect 164528 118522 164556 120006
rect 164988 119354 165016 120142
rect 164620 119326 165016 119354
rect 165724 120006 166152 120034
rect 166368 120006 166704 120034
rect 167104 120006 167348 120034
rect 167656 120006 167992 120034
rect 168392 120006 168544 120034
rect 168852 120006 169188 120034
rect 169740 120006 169984 120034
rect 164516 118516 164568 118522
rect 164516 118458 164568 118464
rect 164620 113880 164648 119326
rect 164436 113852 164648 113880
rect 164436 9450 164464 113852
rect 164424 9444 164476 9450
rect 164424 9386 164476 9392
rect 164332 9308 164384 9314
rect 164332 9250 164384 9256
rect 162860 6316 162912 6322
rect 162860 6258 162912 6264
rect 165724 5370 165752 120006
rect 166368 117774 166396 120006
rect 166356 117768 166408 117774
rect 166356 117710 166408 117716
rect 167000 113892 167052 113898
rect 167000 113834 167052 113840
rect 167012 5438 167040 113834
rect 167104 6390 167132 120006
rect 167656 113898 167684 120006
rect 168392 118658 168420 120006
rect 168852 119354 168880 120006
rect 168484 119326 168880 119354
rect 168380 118652 168432 118658
rect 168380 118594 168432 118600
rect 167644 113892 167696 113898
rect 167644 113834 167696 113840
rect 168484 12510 168512 119326
rect 169852 113892 169904 113898
rect 169852 113834 169904 113840
rect 168472 12504 168524 12510
rect 168472 12446 168524 12452
rect 168380 9716 168432 9722
rect 168380 9658 168432 9664
rect 168392 9518 168420 9658
rect 168380 9512 168432 9518
rect 168380 9454 168432 9460
rect 169864 6458 169892 113834
rect 169852 6452 169904 6458
rect 169852 6394 169904 6400
rect 167092 6384 167144 6390
rect 167092 6326 167144 6332
rect 169956 5506 169984 120006
rect 170048 120006 170384 120034
rect 170692 120006 171028 120034
rect 171244 120006 171580 120034
rect 171888 120006 172224 120034
rect 172624 120006 172868 120034
rect 173084 120006 173420 120034
rect 173912 120006 174064 120034
rect 174372 120006 174708 120034
rect 175260 120006 175412 120034
rect 170048 118114 170076 120006
rect 170036 118108 170088 118114
rect 170036 118050 170088 118056
rect 170692 113898 170720 120006
rect 170680 113892 170732 113898
rect 170680 113834 170732 113840
rect 169944 5500 169996 5506
rect 169944 5442 169996 5448
rect 167000 5432 167052 5438
rect 167000 5374 167052 5380
rect 170588 5432 170640 5438
rect 170588 5374 170640 5380
rect 165712 5364 165764 5370
rect 165712 5306 165764 5312
rect 167092 5364 167144 5370
rect 167092 5306 167144 5312
rect 163504 4480 163556 4486
rect 163504 4422 163556 4428
rect 159916 4140 159968 4146
rect 159916 4082 159968 4088
rect 159088 3392 159140 3398
rect 159088 3334 159140 3340
rect 159928 480 159956 4082
rect 161112 3936 161164 3942
rect 161112 3878 161164 3884
rect 161124 480 161152 3878
rect 162308 3460 162360 3466
rect 162308 3402 162360 3408
rect 162320 480 162348 3402
rect 163516 480 163544 4422
rect 164700 4344 164752 4350
rect 164700 4286 164752 4292
rect 164712 480 164740 4286
rect 165896 3528 165948 3534
rect 165896 3470 165948 3476
rect 165908 480 165936 3470
rect 167104 480 167132 5306
rect 168196 4140 168248 4146
rect 168196 4082 168248 4088
rect 168208 480 168236 4082
rect 169392 3596 169444 3602
rect 169392 3538 169444 3544
rect 169404 480 169432 3538
rect 170600 480 170628 5374
rect 171244 4758 171272 120006
rect 171888 117978 171916 120006
rect 171876 117972 171928 117978
rect 171876 117914 171928 117920
rect 172520 111648 172572 111654
rect 172520 111590 172572 111596
rect 171232 4752 171284 4758
rect 171232 4694 171284 4700
rect 172532 4690 172560 111590
rect 172624 9450 172652 120006
rect 173084 111654 173112 120006
rect 173912 118182 173940 120006
rect 173900 118176 173952 118182
rect 173900 118118 173952 118124
rect 174372 113218 174400 120006
rect 174544 118176 174596 118182
rect 174544 118118 174596 118124
rect 173900 113212 173952 113218
rect 173900 113154 173952 113160
rect 174360 113212 174412 113218
rect 174360 113154 174412 113160
rect 173072 111648 173124 111654
rect 173072 111590 173124 111596
rect 173912 103494 173940 113154
rect 173900 103488 173952 103494
rect 173900 103430 173952 103436
rect 173992 103420 174044 103426
rect 173992 103362 174044 103368
rect 174004 75954 174032 103362
rect 173992 75948 174044 75954
rect 173992 75890 174044 75896
rect 174084 75948 174136 75954
rect 174084 75890 174136 75896
rect 174096 74526 174124 75890
rect 174084 74520 174136 74526
rect 174084 74462 174136 74468
rect 173992 64932 174044 64938
rect 173992 64874 174044 64880
rect 174004 55282 174032 64874
rect 173992 55276 174044 55282
rect 173992 55218 174044 55224
rect 174084 55276 174136 55282
rect 174084 55218 174136 55224
rect 174096 39370 174124 55218
rect 173900 39364 173952 39370
rect 173900 39306 173952 39312
rect 174084 39364 174136 39370
rect 174084 39306 174136 39312
rect 173912 29730 173940 39306
rect 173912 29702 174032 29730
rect 174004 24834 174032 29702
rect 173912 24806 174032 24834
rect 173912 20058 173940 24806
rect 173900 20052 173952 20058
rect 173900 19994 173952 20000
rect 172612 9444 172664 9450
rect 172612 9386 172664 9392
rect 173992 6928 174044 6934
rect 173992 6870 174044 6876
rect 174004 6526 174032 6870
rect 173992 6520 174044 6526
rect 173992 6462 174044 6468
rect 174176 5500 174228 5506
rect 174176 5442 174228 5448
rect 173900 4752 173952 4758
rect 173900 4694 173952 4700
rect 172520 4684 172572 4690
rect 172520 4626 172572 4632
rect 171784 4004 171836 4010
rect 171784 3946 171836 3952
rect 171796 480 171824 3946
rect 173912 3806 173940 4694
rect 173900 3800 173952 3806
rect 173900 3742 173952 3748
rect 172980 3732 173032 3738
rect 172980 3674 173032 3680
rect 172992 480 173020 3674
rect 174188 480 174216 5442
rect 174556 4146 174584 118118
rect 175384 4622 175412 120006
rect 175568 120006 175904 120034
rect 176212 120006 176548 120034
rect 176764 120006 177100 120034
rect 177408 120006 177744 120034
rect 178052 120006 178388 120034
rect 178604 120006 178940 120034
rect 179432 120006 179584 120034
rect 179892 120006 180228 120034
rect 180780 120006 180932 120034
rect 175568 118454 175596 120006
rect 175556 118448 175608 118454
rect 175556 118390 175608 118396
rect 176212 113218 176240 120006
rect 176568 117972 176620 117978
rect 176568 117914 176620 117920
rect 175556 113212 175608 113218
rect 175556 113154 175608 113160
rect 176200 113212 176252 113218
rect 176200 113154 176252 113160
rect 175568 85626 175596 113154
rect 175646 85640 175702 85649
rect 175568 85598 175646 85626
rect 175646 85575 175702 85584
rect 175830 85504 175886 85513
rect 175830 85439 175886 85448
rect 175844 55282 175872 85439
rect 175648 55276 175700 55282
rect 175648 55218 175700 55224
rect 175832 55276 175884 55282
rect 175832 55218 175884 55224
rect 175660 34490 175688 55218
rect 175568 34462 175688 34490
rect 175568 26314 175596 34462
rect 175556 26308 175608 26314
rect 175556 26250 175608 26256
rect 175556 24880 175608 24886
rect 175556 24822 175608 24828
rect 175568 20074 175596 24822
rect 175568 20046 175688 20074
rect 175372 4616 175424 4622
rect 175372 4558 175424 4564
rect 174544 4140 174596 4146
rect 174544 4082 174596 4088
rect 175372 4140 175424 4146
rect 175372 4082 175424 4088
rect 175384 480 175412 4082
rect 175660 3330 175688 20046
rect 176580 4146 176608 117914
rect 176764 4554 176792 120006
rect 177408 118250 177436 120006
rect 177396 118244 177448 118250
rect 177396 118186 177448 118192
rect 178052 25090 178080 120006
rect 178604 113218 178632 120006
rect 178684 118652 178736 118658
rect 178684 118594 178736 118600
rect 178132 113212 178184 113218
rect 178132 113154 178184 113160
rect 178592 113212 178644 113218
rect 178592 113154 178644 113160
rect 178144 103494 178172 113154
rect 178132 103488 178184 103494
rect 178132 103430 178184 103436
rect 178316 103488 178368 103494
rect 178316 103430 178368 103436
rect 178328 75886 178356 103430
rect 178132 75880 178184 75886
rect 178132 75822 178184 75828
rect 178316 75880 178368 75886
rect 178316 75822 178368 75828
rect 178144 64870 178172 75822
rect 178132 64864 178184 64870
rect 178132 64806 178184 64812
rect 178316 64864 178368 64870
rect 178316 64806 178368 64812
rect 178328 59906 178356 64806
rect 178224 59900 178276 59906
rect 178224 59842 178276 59848
rect 178316 59900 178368 59906
rect 178316 59842 178368 59848
rect 178236 52465 178264 59842
rect 178222 52456 178278 52465
rect 178222 52391 178278 52400
rect 178406 52456 178462 52465
rect 178406 52391 178462 52400
rect 178420 47666 178448 52391
rect 178224 47660 178276 47666
rect 178224 47602 178276 47608
rect 178408 47660 178460 47666
rect 178408 47602 178460 47608
rect 178236 31754 178264 47602
rect 178224 31748 178276 31754
rect 178224 31690 178276 31696
rect 178408 31748 178460 31754
rect 178408 31690 178460 31696
rect 178040 25084 178092 25090
rect 178040 25026 178092 25032
rect 178040 24744 178092 24750
rect 178040 24686 178092 24692
rect 178052 6594 178080 24686
rect 178420 22137 178448 31690
rect 178130 22128 178186 22137
rect 178130 22063 178186 22072
rect 178406 22128 178462 22137
rect 178406 22063 178462 22072
rect 178144 12374 178172 22063
rect 178132 12368 178184 12374
rect 178132 12310 178184 12316
rect 178040 6588 178092 6594
rect 178040 6530 178092 6536
rect 177488 6316 177540 6322
rect 177488 6258 177540 6264
rect 176752 4548 176804 4554
rect 176752 4490 176804 4496
rect 176568 4140 176620 4146
rect 176568 4082 176620 4088
rect 177500 3874 177528 6258
rect 177764 4140 177816 4146
rect 177764 4082 177816 4088
rect 177488 3868 177540 3874
rect 177488 3810 177540 3816
rect 176476 3800 176528 3806
rect 176476 3742 176528 3748
rect 175648 3324 175700 3330
rect 175648 3266 175700 3272
rect 176488 1986 176516 3742
rect 176488 1958 176608 1986
rect 176580 480 176608 1958
rect 177776 480 177804 4082
rect 178696 3942 178724 118594
rect 179328 118108 179380 118114
rect 179328 118050 179380 118056
rect 178684 3936 178736 3942
rect 178684 3878 178736 3884
rect 179340 610 179368 118050
rect 179432 118046 179460 120006
rect 179420 118040 179472 118046
rect 179420 117982 179472 117988
rect 179892 113218 179920 120006
rect 180064 118244 180116 118250
rect 180064 118186 180116 118192
rect 179420 113212 179472 113218
rect 179420 113154 179472 113160
rect 179880 113212 179932 113218
rect 179880 113154 179932 113160
rect 179432 103494 179460 113154
rect 179420 103488 179472 103494
rect 179420 103430 179472 103436
rect 179512 103420 179564 103426
rect 179512 103362 179564 103368
rect 179524 89010 179552 103362
rect 179512 89004 179564 89010
rect 179512 88946 179564 88952
rect 179604 84244 179656 84250
rect 179604 84186 179656 84192
rect 179616 66298 179644 84186
rect 179512 66292 179564 66298
rect 179512 66234 179564 66240
rect 179604 66292 179656 66298
rect 179604 66234 179656 66240
rect 179524 58698 179552 66234
rect 179432 58670 179552 58698
rect 179432 53802 179460 58670
rect 179432 53774 179552 53802
rect 179524 51134 179552 53774
rect 179512 51128 179564 51134
rect 179512 51070 179564 51076
rect 179420 51060 179472 51066
rect 179420 51002 179472 51008
rect 179432 26314 179460 51002
rect 179420 26308 179472 26314
rect 179420 26250 179472 26256
rect 179512 26308 179564 26314
rect 179512 26250 179564 26256
rect 179524 24818 179552 26250
rect 179512 24812 179564 24818
rect 179512 24754 179564 24760
rect 179420 6928 179472 6934
rect 179420 6870 179472 6876
rect 179432 6730 179460 6870
rect 179420 6724 179472 6730
rect 179420 6666 179472 6672
rect 180076 4146 180104 118186
rect 180904 6662 180932 120006
rect 181088 120006 181424 120034
rect 180984 119808 181036 119814
rect 180984 119750 181036 119756
rect 180996 113150 181024 119750
rect 181088 118590 181116 120006
rect 182054 119814 182082 120020
rect 182284 120006 182620 120034
rect 182928 120006 183264 120034
rect 183572 120006 183908 120034
rect 184032 120006 184460 120034
rect 184952 120006 185104 120034
rect 182042 119808 182094 119814
rect 182042 119750 182094 119756
rect 181076 118584 181128 118590
rect 181076 118526 181128 118532
rect 180984 113144 181036 113150
rect 180984 113086 181036 113092
rect 181076 104780 181128 104786
rect 181076 104722 181128 104728
rect 181088 95266 181116 104722
rect 181076 95260 181128 95266
rect 181076 95202 181128 95208
rect 181168 95124 181220 95130
rect 181168 95066 181220 95072
rect 181180 92478 181208 95066
rect 181168 92472 181220 92478
rect 181168 92414 181220 92420
rect 181260 82884 181312 82890
rect 181260 82826 181312 82832
rect 181272 76022 181300 82826
rect 181260 76016 181312 76022
rect 181260 75958 181312 75964
rect 181076 75880 181128 75886
rect 181076 75822 181128 75828
rect 181088 73166 181116 75822
rect 181076 73160 181128 73166
rect 181076 73102 181128 73108
rect 181076 63572 181128 63578
rect 181076 63514 181128 63520
rect 181088 61062 181116 63514
rect 181076 61056 181128 61062
rect 181076 60998 181128 61004
rect 181168 50652 181220 50658
rect 181168 50594 181220 50600
rect 181180 44130 181208 50594
rect 181168 44124 181220 44130
rect 181168 44066 181220 44072
rect 181168 31680 181220 31686
rect 181168 31622 181220 31628
rect 181180 22166 181208 31622
rect 181168 22160 181220 22166
rect 181168 22102 181220 22108
rect 181076 22092 181128 22098
rect 181076 22034 181128 22040
rect 180892 6656 180944 6662
rect 180892 6598 180944 6604
rect 180064 4140 180116 4146
rect 180064 4082 180116 4088
rect 180156 3868 180208 3874
rect 180156 3810 180208 3816
rect 178960 604 179012 610
rect 178960 546 179012 552
rect 179328 604 179380 610
rect 179328 546 179380 552
rect 178972 480 179000 546
rect 180168 480 180196 3810
rect 181088 3330 181116 22034
rect 182284 6798 182312 120006
rect 182928 118318 182956 120006
rect 182916 118312 182968 118318
rect 182916 118254 182968 118260
rect 183468 118040 183520 118046
rect 183468 117982 183520 117988
rect 182272 6792 182324 6798
rect 182272 6734 182324 6740
rect 183480 4146 183508 117982
rect 183572 9518 183600 120006
rect 184032 119354 184060 120006
rect 183756 119326 184060 119354
rect 183756 115938 183784 119326
rect 184848 118312 184900 118318
rect 184848 118254 184900 118260
rect 183744 115932 183796 115938
rect 183744 115874 183796 115880
rect 183928 115932 183980 115938
rect 183928 115874 183980 115880
rect 184756 115932 184808 115938
rect 184756 115874 184808 115880
rect 183940 106321 183968 115874
rect 184768 106321 184796 115874
rect 183650 106312 183706 106321
rect 183650 106247 183706 106256
rect 183926 106312 183982 106321
rect 183926 106247 183982 106256
rect 184754 106312 184810 106321
rect 184754 106247 184810 106256
rect 183664 106214 183692 106247
rect 183652 106208 183704 106214
rect 183652 106150 183704 106156
rect 183928 106208 183980 106214
rect 183928 106150 183980 106156
rect 183940 96665 183968 106150
rect 183742 96656 183798 96665
rect 183742 96591 183798 96600
rect 183926 96656 183982 96665
rect 183926 96591 183982 96600
rect 183756 86970 183784 96591
rect 183744 86964 183796 86970
rect 183744 86906 183796 86912
rect 183928 86964 183980 86970
rect 183928 86906 183980 86912
rect 183940 75886 183968 86906
rect 184860 77382 184888 118254
rect 184952 117609 184980 120006
rect 185734 119814 185762 120020
rect 185124 119808 185176 119814
rect 185124 119750 185176 119756
rect 185722 119808 185774 119814
rect 185722 119750 185774 119756
rect 186286 119762 186314 120020
rect 186608 120006 186944 120034
rect 187068 120006 187496 120034
rect 187712 120006 188140 120034
rect 188448 120006 188784 120034
rect 184938 117600 184994 117609
rect 184938 117535 184994 117544
rect 185136 115954 185164 119750
rect 186286 119734 186360 119762
rect 186228 118448 186280 118454
rect 186228 118390 186280 118396
rect 185584 117700 185636 117706
rect 185584 117642 185636 117648
rect 185044 115938 185164 115954
rect 185032 115932 185164 115938
rect 185084 115926 185164 115932
rect 185032 115874 185084 115880
rect 185044 115843 185072 115874
rect 184938 106312 184994 106321
rect 184938 106247 184994 106256
rect 184952 96642 184980 106247
rect 184952 96614 185072 96642
rect 185044 91746 185072 96614
rect 184952 91718 185072 91746
rect 184952 77466 184980 91718
rect 184952 77438 185072 77466
rect 184848 77376 184900 77382
rect 184848 77318 184900 77324
rect 184848 77172 184900 77178
rect 184848 77114 184900 77120
rect 184756 77104 184808 77110
rect 184756 77046 184808 77052
rect 183928 75880 183980 75886
rect 183928 75822 183980 75828
rect 184768 67658 184796 77046
rect 184756 67652 184808 67658
rect 184756 67594 184808 67600
rect 183744 66360 183796 66366
rect 183744 66302 183796 66308
rect 183756 66230 183784 66302
rect 183744 66224 183796 66230
rect 183744 66166 183796 66172
rect 183744 56636 183796 56642
rect 183744 56578 183796 56584
rect 183756 48385 183784 56578
rect 183742 48376 183798 48385
rect 183742 48311 183798 48320
rect 183650 38720 183706 38729
rect 183650 38655 183706 38664
rect 183664 33810 183692 38655
rect 183664 33782 183784 33810
rect 183756 28966 183784 33782
rect 183744 28960 183796 28966
rect 183744 28902 183796 28908
rect 183744 28824 183796 28830
rect 183744 28766 183796 28772
rect 183756 12510 183784 28766
rect 183744 12504 183796 12510
rect 183744 12446 183796 12452
rect 183652 12436 183704 12442
rect 183652 12378 183704 12384
rect 183664 9654 183692 12378
rect 183652 9648 183704 9654
rect 183652 9590 183704 9596
rect 183560 9512 183612 9518
rect 183560 9454 183612 9460
rect 183560 6248 183612 6254
rect 183560 6190 183612 6196
rect 182548 4140 182600 4146
rect 182548 4082 182600 4088
rect 183468 4140 183520 4146
rect 183468 4082 183520 4088
rect 181076 3324 181128 3330
rect 181076 3266 181128 3272
rect 181352 3188 181404 3194
rect 181352 3130 181404 3136
rect 181364 480 181392 3130
rect 182560 480 182588 4082
rect 183572 4010 183600 6190
rect 183560 4004 183612 4010
rect 183560 3946 183612 3952
rect 183744 3936 183796 3942
rect 183744 3878 183796 3884
rect 183756 480 183784 3878
rect 184860 480 184888 77114
rect 185044 77110 185072 77438
rect 185032 77104 185084 77110
rect 185032 77046 185084 77052
rect 184940 67652 184992 67658
rect 184940 67594 184992 67600
rect 184952 60858 184980 67594
rect 184940 60852 184992 60858
rect 184940 60794 184992 60800
rect 184940 57928 184992 57934
rect 184940 57870 184992 57876
rect 184952 51134 184980 57870
rect 184940 51128 184992 51134
rect 184940 51070 184992 51076
rect 184940 48340 184992 48346
rect 184940 48282 184992 48288
rect 184952 41290 184980 48282
rect 184952 41262 185072 41290
rect 185044 28966 185072 41262
rect 185032 28960 185084 28966
rect 185032 28902 185084 28908
rect 184940 19372 184992 19378
rect 184940 19314 184992 19320
rect 184952 3262 184980 19314
rect 184940 3256 184992 3262
rect 184940 3198 184992 3204
rect 185596 2854 185624 117642
rect 185584 2848 185636 2854
rect 185584 2790 185636 2796
rect 186240 626 186268 118390
rect 186332 6050 186360 119734
rect 186608 118561 186636 120006
rect 187068 119354 187096 120006
rect 186700 119326 187096 119354
rect 186594 118552 186650 118561
rect 186594 118487 186650 118496
rect 186700 113914 186728 119326
rect 186424 113886 186728 113914
rect 186424 21978 186452 113886
rect 186424 21950 186544 21978
rect 186320 6044 186372 6050
rect 186320 5986 186372 5992
rect 186516 5982 186544 21950
rect 186504 5976 186556 5982
rect 186504 5918 186556 5924
rect 187712 5914 187740 120006
rect 188448 118153 188476 120006
rect 189322 119762 189350 120020
rect 189276 119734 189350 119762
rect 189644 120006 189980 120034
rect 190288 120006 190624 120034
rect 190748 120006 191176 120034
rect 191820 120006 191972 120034
rect 188434 118144 188490 118153
rect 188434 118079 188490 118088
rect 188448 117337 188476 118079
rect 187790 117328 187846 117337
rect 187790 117263 187846 117272
rect 188434 117328 188490 117337
rect 188434 117263 188490 117272
rect 187804 8906 187832 117263
rect 189172 113892 189224 113898
rect 189172 113834 189224 113840
rect 187792 8900 187844 8906
rect 187792 8842 187844 8848
rect 187700 5908 187752 5914
rect 187700 5850 187752 5856
rect 189184 5846 189212 113834
rect 189172 5840 189224 5846
rect 189172 5782 189224 5788
rect 187240 4072 187292 4078
rect 187240 4014 187292 4020
rect 186056 598 186268 626
rect 186056 480 186084 598
rect 187252 480 187280 4014
rect 188436 4004 188488 4010
rect 188436 3946 188488 3952
rect 188448 480 188476 3946
rect 189276 3126 189304 119734
rect 189644 113898 189672 120006
rect 190288 117366 190316 120006
rect 190368 118516 190420 118522
rect 190368 118458 190420 118464
rect 190276 117360 190328 117366
rect 190276 117302 190328 117308
rect 189632 113892 189684 113898
rect 189632 113834 189684 113840
rect 190380 3398 190408 118458
rect 190552 117360 190604 117366
rect 190552 117302 190604 117308
rect 190564 116822 190592 117302
rect 190552 116816 190604 116822
rect 190552 116758 190604 116764
rect 190564 8770 190592 116758
rect 190748 86970 190776 120006
rect 191840 113892 191892 113898
rect 191840 113834 191892 113840
rect 190736 86964 190788 86970
rect 190736 86906 190788 86912
rect 190828 77308 190880 77314
rect 190828 77250 190880 77256
rect 190840 67726 190868 77250
rect 190828 67720 190880 67726
rect 190828 67662 190880 67668
rect 190736 67652 190788 67658
rect 190736 67594 190788 67600
rect 190748 66230 190776 67594
rect 190736 66224 190788 66230
rect 190736 66166 190788 66172
rect 190828 66224 190880 66230
rect 190828 66166 190880 66172
rect 190840 46918 190868 66166
rect 190828 46912 190880 46918
rect 190828 46854 190880 46860
rect 190736 29028 190788 29034
rect 190736 28970 190788 28976
rect 190748 19446 190776 28970
rect 190736 19440 190788 19446
rect 190736 19382 190788 19388
rect 190644 18012 190696 18018
rect 190644 17954 190696 17960
rect 190656 9722 190684 17954
rect 190644 9716 190696 9722
rect 190644 9658 190696 9664
rect 190736 9716 190788 9722
rect 190736 9658 190788 9664
rect 190552 8764 190604 8770
rect 190552 8706 190604 8712
rect 190748 8514 190776 9658
rect 190564 8486 190776 8514
rect 190564 5710 190592 8486
rect 190552 5704 190604 5710
rect 190552 5646 190604 5652
rect 190828 4140 190880 4146
rect 190828 4082 190880 4088
rect 189632 3392 189684 3398
rect 189632 3334 189684 3340
rect 190368 3392 190420 3398
rect 190368 3334 190420 3340
rect 189264 3120 189316 3126
rect 189264 3062 189316 3068
rect 189644 480 189672 3334
rect 190840 480 190868 4082
rect 191852 3058 191880 113834
rect 191944 5778 191972 120006
rect 192036 120006 192464 120034
rect 192680 120006 193016 120034
rect 193232 120006 193660 120034
rect 193968 120006 194304 120034
rect 194612 120006 194856 120034
rect 195164 120006 195500 120034
rect 195992 120006 196144 120034
rect 196452 120006 196696 120034
rect 197340 120006 197492 120034
rect 192036 117162 192064 120006
rect 192484 117632 192536 117638
rect 192484 117574 192536 117580
rect 192024 117156 192076 117162
rect 192024 117098 192076 117104
rect 192036 6225 192064 117098
rect 192022 6216 192078 6225
rect 192022 6151 192078 6160
rect 191932 5772 191984 5778
rect 191932 5714 191984 5720
rect 192024 3256 192076 3262
rect 192024 3198 192076 3204
rect 191840 3052 191892 3058
rect 191840 2994 191892 3000
rect 192036 480 192064 3198
rect 192496 2922 192524 117574
rect 192680 113898 192708 120006
rect 192668 113892 192720 113898
rect 192668 113834 192720 113840
rect 193232 5642 193260 120006
rect 193968 118425 193996 120006
rect 193954 118416 194010 118425
rect 193954 118351 194010 118360
rect 194508 118380 194560 118386
rect 194508 118322 194560 118328
rect 193220 5636 193272 5642
rect 193220 5578 193272 5584
rect 194520 3058 194548 118322
rect 194612 7546 194640 120006
rect 195164 119354 195192 120006
rect 194796 119326 195192 119354
rect 194796 109750 194824 119326
rect 195888 118584 195940 118590
rect 195888 118526 195940 118532
rect 194784 109744 194836 109750
rect 194784 109686 194836 109692
rect 194692 104916 194744 104922
rect 194692 104858 194744 104864
rect 194704 104825 194732 104858
rect 194690 104816 194746 104825
rect 194690 104751 194746 104760
rect 194966 104680 195022 104689
rect 194966 104615 195022 104624
rect 194980 95282 195008 104615
rect 194796 95254 195008 95282
rect 194796 89758 194824 95254
rect 194784 89752 194836 89758
rect 194784 89694 194836 89700
rect 194876 89616 194928 89622
rect 194876 89558 194928 89564
rect 194888 85542 194916 89558
rect 194876 85536 194928 85542
rect 194876 85478 194928 85484
rect 194876 75948 194928 75954
rect 194876 75890 194928 75896
rect 194888 70514 194916 75890
rect 194876 70508 194928 70514
rect 194876 70450 194928 70456
rect 194784 70372 194836 70378
rect 194784 70314 194836 70320
rect 194796 66230 194824 70314
rect 194784 66224 194836 66230
rect 194784 66166 194836 66172
rect 195152 56636 195204 56642
rect 195152 56578 195204 56584
rect 195164 48385 195192 56578
rect 194966 48376 195022 48385
rect 194966 48311 195022 48320
rect 195150 48376 195206 48385
rect 195150 48311 195206 48320
rect 194980 46918 195008 48311
rect 194968 46912 195020 46918
rect 194968 46854 195020 46860
rect 194692 37324 194744 37330
rect 194692 37266 194744 37272
rect 194704 31634 194732 37266
rect 194704 31606 194824 31634
rect 194796 22114 194824 31606
rect 194704 22086 194824 22114
rect 194704 21978 194732 22086
rect 194704 21950 194824 21978
rect 194796 8838 194824 21950
rect 194784 8832 194836 8838
rect 194784 8774 194836 8780
rect 194600 7540 194652 7546
rect 194600 7482 194652 7488
rect 193220 3052 193272 3058
rect 193220 2994 193272 3000
rect 194508 3052 194560 3058
rect 194508 2994 194560 3000
rect 192484 2916 192536 2922
rect 192484 2858 192536 2864
rect 193232 480 193260 2994
rect 194416 1352 194468 1358
rect 194416 1294 194468 1300
rect 194428 480 194456 1294
rect 195900 626 195928 118526
rect 195992 117366 196020 120006
rect 195980 117360 196032 117366
rect 195980 117302 196032 117308
rect 196452 116634 196480 120006
rect 197268 117904 197320 117910
rect 197268 117846 197320 117852
rect 196084 116606 196480 116634
rect 196084 7478 196112 116606
rect 196072 7472 196124 7478
rect 196072 7414 196124 7420
rect 197280 3670 197308 117846
rect 197360 116612 197412 116618
rect 197360 116554 197412 116560
rect 196808 3664 196860 3670
rect 196808 3606 196860 3612
rect 197268 3664 197320 3670
rect 197268 3606 197320 3612
rect 195624 598 195928 626
rect 195624 480 195652 598
rect 196820 480 196848 3606
rect 197372 2990 197400 116554
rect 197464 5574 197492 120006
rect 197648 120006 197984 120034
rect 198200 120006 198536 120034
rect 198844 120006 199180 120034
rect 199488 120006 199824 120034
rect 200132 120006 200376 120034
rect 197648 118289 197676 120006
rect 197634 118280 197690 118289
rect 197634 118215 197690 118224
rect 198004 117564 198056 117570
rect 198004 117506 198056 117512
rect 197452 5568 197504 5574
rect 197452 5510 197504 5516
rect 198016 3482 198044 117506
rect 198200 116618 198228 120006
rect 198188 116612 198240 116618
rect 198188 116554 198240 116560
rect 198740 116612 198792 116618
rect 198740 116554 198792 116560
rect 198752 8226 198780 116554
rect 198740 8220 198792 8226
rect 198740 8162 198792 8168
rect 198844 7410 198872 120006
rect 199488 116618 199516 120006
rect 199476 116612 199528 116618
rect 199476 116554 199528 116560
rect 198832 7404 198884 7410
rect 198832 7346 198884 7352
rect 200132 7342 200160 120006
rect 200500 116634 200528 120142
rect 201650 119762 201678 120020
rect 201604 119734 201678 119762
rect 201880 120006 202216 120034
rect 201408 117836 201460 117842
rect 201408 117778 201460 117784
rect 200224 116606 200528 116634
rect 200224 113150 200252 116606
rect 200212 113144 200264 113150
rect 200212 113086 200264 113092
rect 200396 113144 200448 113150
rect 200396 113086 200448 113092
rect 200408 109018 200436 113086
rect 200316 108990 200436 109018
rect 200316 100042 200344 108990
rect 200224 100014 200344 100042
rect 200224 94058 200252 100014
rect 200224 94030 200436 94058
rect 200408 89570 200436 94030
rect 200316 89542 200436 89570
rect 200316 85542 200344 89542
rect 200304 85536 200356 85542
rect 200304 85478 200356 85484
rect 200304 75948 200356 75954
rect 200304 75890 200356 75896
rect 200316 67658 200344 75890
rect 200304 67652 200356 67658
rect 200304 67594 200356 67600
rect 200396 67652 200448 67658
rect 200396 67594 200448 67600
rect 200408 57934 200436 67594
rect 200396 57928 200448 57934
rect 200396 57870 200448 57876
rect 200304 48340 200356 48346
rect 200304 48282 200356 48288
rect 200316 41426 200344 48282
rect 200316 41398 200528 41426
rect 200500 38622 200528 41398
rect 200488 38616 200540 38622
rect 200488 38558 200540 38564
rect 200396 29028 200448 29034
rect 200396 28970 200448 28976
rect 200408 22114 200436 28970
rect 200224 22098 200436 22114
rect 200212 22092 200448 22098
rect 200264 22086 200396 22092
rect 200212 22034 200264 22040
rect 200396 22034 200448 22040
rect 200408 19310 200436 22034
rect 200396 19304 200448 19310
rect 200396 19246 200448 19252
rect 200396 12300 200448 12306
rect 200396 12242 200448 12248
rect 200120 7336 200172 7342
rect 200120 7278 200172 7284
rect 200408 7274 200436 12242
rect 200396 7268 200448 7274
rect 200396 7210 200448 7216
rect 201420 3670 201448 117778
rect 201500 116612 201552 116618
rect 201500 116554 201552 116560
rect 201512 7138 201540 116554
rect 201604 7206 201632 119734
rect 201880 116618 201908 120006
rect 202972 116680 203024 116686
rect 202972 116622 203024 116628
rect 201868 116612 201920 116618
rect 201868 116554 201920 116560
rect 202880 116612 202932 116618
rect 202880 116554 202932 116560
rect 202892 7818 202920 116554
rect 202880 7812 202932 7818
rect 202880 7754 202932 7760
rect 202984 7614 203012 116622
rect 203076 8294 203104 120142
rect 203168 120006 203504 120034
rect 203720 120006 204056 120034
rect 204364 120006 204700 120034
rect 204916 120006 205252 120034
rect 205652 120006 205896 120034
rect 206204 120006 206540 120034
rect 203168 116686 203196 120006
rect 203156 116680 203208 116686
rect 203156 116622 203208 116628
rect 203720 116618 203748 120006
rect 203708 116612 203760 116618
rect 203708 116554 203760 116560
rect 204260 116612 204312 116618
rect 204260 116554 204312 116560
rect 203064 8288 203116 8294
rect 203064 8230 203116 8236
rect 202972 7608 203024 7614
rect 202972 7550 203024 7556
rect 201592 7200 201644 7206
rect 201592 7142 201644 7148
rect 201500 7132 201552 7138
rect 201500 7074 201552 7080
rect 204272 5098 204300 116554
rect 204364 7682 204392 120006
rect 204916 116618 204944 120006
rect 204904 116612 204956 116618
rect 204904 116554 204956 116560
rect 205548 12164 205600 12170
rect 205548 12106 205600 12112
rect 205560 7886 205588 12106
rect 205548 7880 205600 7886
rect 205548 7822 205600 7828
rect 205652 7750 205680 120006
rect 206204 119354 206232 120006
rect 207078 119762 207106 120020
rect 205928 119326 206232 119354
rect 207032 119734 207106 119762
rect 207308 120006 207736 120034
rect 208380 120006 208532 120034
rect 205928 109138 205956 119326
rect 205916 109132 205968 109138
rect 205916 109074 205968 109080
rect 205916 108996 205968 109002
rect 205916 108938 205968 108944
rect 205928 103442 205956 108938
rect 205928 103414 206048 103442
rect 206020 93974 206048 103414
rect 206008 93968 206060 93974
rect 206008 93910 206060 93916
rect 205916 93832 205968 93838
rect 205916 93774 205968 93780
rect 205928 91089 205956 93774
rect 205914 91080 205970 91089
rect 205914 91015 205970 91024
rect 206098 91080 206154 91089
rect 206098 91015 206154 91024
rect 206112 81462 206140 91015
rect 205916 81456 205968 81462
rect 205916 81398 205968 81404
rect 206100 81456 206152 81462
rect 206100 81398 206152 81404
rect 205928 80170 205956 81398
rect 205916 80164 205968 80170
rect 205916 80106 205968 80112
rect 205916 74112 205968 74118
rect 205916 74054 205968 74060
rect 205928 60858 205956 74054
rect 205916 60852 205968 60858
rect 205916 60794 205968 60800
rect 205824 57996 205876 58002
rect 205824 57938 205876 57944
rect 205836 51762 205864 57938
rect 205836 51734 205956 51762
rect 205928 22234 205956 51734
rect 205916 22228 205968 22234
rect 205916 22170 205968 22176
rect 205732 19372 205784 19378
rect 205732 19314 205784 19320
rect 205744 12170 205772 19314
rect 205732 12164 205784 12170
rect 205732 12106 205784 12112
rect 205640 7744 205692 7750
rect 205640 7686 205692 7692
rect 204352 7676 204404 7682
rect 204352 7618 204404 7624
rect 204260 5092 204312 5098
rect 204260 5034 204312 5040
rect 204352 5092 204404 5098
rect 204352 5034 204404 5040
rect 202880 4616 202932 4622
rect 202880 4558 202932 4564
rect 200396 3664 200448 3670
rect 200396 3606 200448 3612
rect 201408 3664 201460 3670
rect 201408 3606 201460 3612
rect 201500 3664 201552 3670
rect 201500 3606 201552 3612
rect 197924 3454 198044 3482
rect 197924 3398 197952 3454
rect 197912 3392 197964 3398
rect 197912 3334 197964 3340
rect 198004 3324 198056 3330
rect 198004 3266 198056 3272
rect 197360 2984 197412 2990
rect 197360 2926 197412 2932
rect 198016 480 198044 3266
rect 199200 3256 199252 3262
rect 199200 3198 199252 3204
rect 199212 480 199240 3198
rect 200408 480 200436 3606
rect 201512 480 201540 3606
rect 202696 3256 202748 3262
rect 202696 3198 202748 3204
rect 202708 480 202736 3198
rect 202892 3058 202920 4558
rect 204260 4548 204312 4554
rect 204260 4490 204312 4496
rect 204272 3330 204300 4490
rect 204364 3670 204392 5034
rect 207032 4826 207060 119734
rect 207308 119354 207336 120006
rect 207124 119326 207336 119354
rect 207124 109138 207152 119326
rect 208308 117768 208360 117774
rect 208308 117710 208360 117716
rect 207112 109132 207164 109138
rect 207112 109074 207164 109080
rect 207112 108996 207164 109002
rect 207112 108938 207164 108944
rect 207124 91050 207152 108938
rect 207112 91044 207164 91050
rect 207112 90986 207164 90992
rect 207204 81456 207256 81462
rect 207204 81398 207256 81404
rect 207216 80170 207244 81398
rect 207204 80164 207256 80170
rect 207204 80106 207256 80112
rect 207204 76628 207256 76634
rect 207204 76570 207256 76576
rect 207216 66230 207244 76570
rect 207204 66224 207256 66230
rect 207204 66166 207256 66172
rect 207112 56636 207164 56642
rect 207112 56578 207164 56584
rect 207124 47054 207152 56578
rect 207112 47048 207164 47054
rect 207112 46990 207164 46996
rect 207204 46980 207256 46986
rect 207204 46922 207256 46928
rect 207216 45558 207244 46922
rect 207204 45552 207256 45558
rect 207204 45494 207256 45500
rect 207204 35964 207256 35970
rect 207204 35906 207256 35912
rect 207216 28966 207244 35906
rect 207204 28960 207256 28966
rect 207204 28902 207256 28908
rect 207296 28960 207348 28966
rect 207296 28902 207348 28908
rect 207308 19417 207336 28902
rect 207294 19408 207350 19417
rect 207294 19343 207350 19352
rect 207294 19272 207350 19281
rect 207294 19207 207350 19216
rect 207308 12322 207336 19207
rect 207216 12294 207336 12322
rect 207216 7954 207244 12294
rect 207204 7948 207256 7954
rect 207204 7890 207256 7896
rect 207020 4820 207072 4826
rect 207020 4762 207072 4768
rect 208216 4820 208268 4826
rect 208216 4762 208268 4768
rect 204352 3664 204404 3670
rect 204352 3606 204404 3612
rect 207480 3664 207532 3670
rect 207480 3606 207532 3612
rect 204260 3324 204312 3330
rect 204260 3266 204312 3272
rect 206284 3120 206336 3126
rect 206284 3062 206336 3068
rect 202880 3052 202932 3058
rect 202880 2994 202932 3000
rect 203892 2984 203944 2990
rect 203892 2926 203944 2932
rect 203904 480 203932 2926
rect 205088 2848 205140 2854
rect 205088 2790 205140 2796
rect 205100 480 205128 2790
rect 206296 480 206324 3062
rect 207492 480 207520 3606
rect 208228 2854 208256 4762
rect 208320 3670 208348 117710
rect 208504 8022 208532 120006
rect 208596 120006 208932 120034
rect 209240 120006 209576 120034
rect 209976 120006 210220 120034
rect 210436 120006 210772 120034
rect 211172 120006 211416 120034
rect 211724 120006 212060 120034
rect 208492 8016 208544 8022
rect 208492 7958 208544 7964
rect 208596 4894 208624 120006
rect 209240 117706 209268 120006
rect 209228 117700 209280 117706
rect 209228 117642 209280 117648
rect 209976 117570 210004 120006
rect 210436 119354 210464 120006
rect 210068 119326 210464 119354
rect 209964 117564 210016 117570
rect 209964 117506 210016 117512
rect 210068 113914 210096 119326
rect 211068 117700 211120 117706
rect 211068 117642 211120 117648
rect 209884 113886 210096 113914
rect 209884 99482 209912 113886
rect 209872 99476 209924 99482
rect 209872 99418 209924 99424
rect 209872 99340 209924 99346
rect 209872 99282 209924 99288
rect 209884 70514 209912 99282
rect 209872 70508 209924 70514
rect 209872 70450 209924 70456
rect 209872 67652 209924 67658
rect 209872 67594 209924 67600
rect 209884 51202 209912 67594
rect 209872 51196 209924 51202
rect 209872 51138 209924 51144
rect 209872 46980 209924 46986
rect 209872 46922 209924 46928
rect 209884 4962 209912 46922
rect 209872 4956 209924 4962
rect 209872 4898 209924 4904
rect 208584 4888 208636 4894
rect 208584 4830 208636 4836
rect 208676 4684 208728 4690
rect 208676 4626 208728 4632
rect 208308 3664 208360 3670
rect 208308 3606 208360 3612
rect 208216 2848 208268 2854
rect 208216 2790 208268 2796
rect 208688 480 208716 4626
rect 211080 3670 211108 117642
rect 211172 117638 211200 120006
rect 211724 119354 211752 120006
rect 212598 119762 212626 120020
rect 211356 119326 211752 119354
rect 212552 119734 212626 119762
rect 212828 120006 213256 120034
rect 211160 117632 211212 117638
rect 211160 117574 211212 117580
rect 211356 105618 211384 119326
rect 211264 105590 211384 105618
rect 211264 100745 211292 105590
rect 211250 100736 211306 100745
rect 211250 100671 211306 100680
rect 211434 100600 211490 100609
rect 211434 100535 211490 100544
rect 211448 81462 211476 100535
rect 211344 81456 211396 81462
rect 211344 81398 211396 81404
rect 211436 81456 211488 81462
rect 211436 81398 211488 81404
rect 211356 75886 211384 81398
rect 211344 75880 211396 75886
rect 211344 75822 211396 75828
rect 211252 66292 211304 66298
rect 211252 66234 211304 66240
rect 211264 64410 211292 66234
rect 211172 64382 211292 64410
rect 211172 56817 211200 64382
rect 212552 57934 212580 119734
rect 212828 119354 212856 120006
rect 213886 119762 213914 120020
rect 214116 120006 214452 120034
rect 214576 120006 215096 120034
rect 215404 120006 215740 120034
rect 215956 120006 216292 120034
rect 216692 120006 216936 120034
rect 217152 120006 217580 120034
rect 213886 119734 213960 119762
rect 212644 119326 212856 119354
rect 212644 110430 212672 119326
rect 213828 117632 213880 117638
rect 213828 117574 213880 117580
rect 213184 117496 213236 117502
rect 213184 117438 213236 117444
rect 212632 110424 212684 110430
rect 212632 110366 212684 110372
rect 212724 100768 212776 100774
rect 212724 100710 212776 100716
rect 212736 91118 212764 100710
rect 212724 91112 212776 91118
rect 212724 91054 212776 91060
rect 212908 91112 212960 91118
rect 212908 91054 212960 91060
rect 212920 86306 212948 91054
rect 212828 86278 212948 86306
rect 212828 73302 212856 86278
rect 212816 73296 212868 73302
rect 212816 73238 212868 73244
rect 212724 73228 212776 73234
rect 212724 73170 212776 73176
rect 212736 68406 212764 73170
rect 212724 68400 212776 68406
rect 212724 68342 212776 68348
rect 212540 57928 212592 57934
rect 212540 57870 212592 57876
rect 212724 57928 212776 57934
rect 212724 57870 212776 57876
rect 211158 56808 211214 56817
rect 211158 56743 211214 56752
rect 211250 56536 211306 56545
rect 211250 56471 211306 56480
rect 211264 46986 211292 56471
rect 212540 51128 212592 51134
rect 212540 51070 212592 51076
rect 211252 46980 211304 46986
rect 211252 46922 211304 46928
rect 211252 45620 211304 45626
rect 211252 45562 211304 45568
rect 211264 45506 211292 45562
rect 211342 45520 211398 45529
rect 211264 45478 211342 45506
rect 211342 45455 211398 45464
rect 211526 45520 211582 45529
rect 211526 45455 211582 45464
rect 211540 40730 211568 45455
rect 211344 40724 211396 40730
rect 211344 40666 211396 40672
rect 211528 40724 211580 40730
rect 211528 40666 211580 40672
rect 211356 27674 211384 40666
rect 211160 27668 211212 27674
rect 211160 27610 211212 27616
rect 211344 27668 211396 27674
rect 211344 27610 211396 27616
rect 211172 19378 211200 27610
rect 211160 19372 211212 19378
rect 211160 19314 211212 19320
rect 211344 19372 211396 19378
rect 211344 19314 211396 19320
rect 211356 12510 211384 19314
rect 211344 12504 211396 12510
rect 211344 12446 211396 12452
rect 211252 12436 211304 12442
rect 211252 12378 211304 12384
rect 211264 4758 211292 12378
rect 212552 5030 212580 51070
rect 212736 38690 212764 57870
rect 212632 38684 212684 38690
rect 212632 38626 212684 38632
rect 212724 38684 212776 38690
rect 212724 38626 212776 38632
rect 212644 38570 212672 38626
rect 212644 38542 212764 38570
rect 212736 22166 212764 38542
rect 212724 22160 212776 22166
rect 212724 22102 212776 22108
rect 212724 22024 212776 22030
rect 212724 21966 212776 21972
rect 212736 6186 212764 21966
rect 212724 6180 212776 6186
rect 212724 6122 212776 6128
rect 212540 5024 212592 5030
rect 212540 4966 212592 4972
rect 212264 4888 212316 4894
rect 212264 4830 212316 4836
rect 211252 4752 211304 4758
rect 211252 4694 211304 4700
rect 209872 3664 209924 3670
rect 209872 3606 209924 3612
rect 211068 3664 211120 3670
rect 211068 3606 211120 3612
rect 209884 480 209912 3606
rect 211068 3052 211120 3058
rect 211068 2994 211120 3000
rect 211080 480 211108 2994
rect 212276 480 212304 4830
rect 213196 2854 213224 117438
rect 213184 2848 213236 2854
rect 213184 2790 213236 2796
rect 213840 626 213868 117574
rect 213932 114034 213960 119734
rect 213920 114028 213972 114034
rect 213920 113970 213972 113976
rect 214116 113898 214144 120006
rect 214196 114028 214248 114034
rect 214196 113970 214248 113976
rect 213920 113892 213972 113898
rect 213920 113834 213972 113840
rect 214104 113892 214156 113898
rect 214104 113834 214156 113840
rect 213932 5234 213960 113834
rect 214208 109154 214236 113970
rect 214024 109126 214236 109154
rect 213920 5228 213972 5234
rect 213920 5170 213972 5176
rect 214024 5166 214052 109126
rect 214576 109070 214604 120006
rect 215300 113892 215352 113898
rect 215300 113834 215352 113840
rect 214104 109064 214156 109070
rect 214104 109006 214156 109012
rect 214564 109064 214616 109070
rect 214564 109006 214616 109012
rect 214116 22098 214144 109006
rect 214104 22092 214156 22098
rect 214104 22034 214156 22040
rect 214196 22024 214248 22030
rect 214196 21966 214248 21972
rect 214208 6322 214236 21966
rect 214196 6316 214248 6322
rect 214196 6258 214248 6264
rect 214012 5160 214064 5166
rect 214012 5102 214064 5108
rect 215312 4282 215340 113834
rect 215404 5302 215432 120006
rect 215956 113898 215984 120006
rect 216692 118658 216720 120006
rect 216680 118652 216732 118658
rect 216680 118594 216732 118600
rect 215944 113892 215996 113898
rect 215944 113834 215996 113840
rect 217152 109018 217180 120006
rect 218118 119762 218146 120020
rect 218440 120006 218776 120034
rect 219420 120006 219664 120034
rect 218118 119734 218192 119762
rect 217324 118652 217376 118658
rect 217324 118594 217376 118600
rect 216876 108990 217180 109018
rect 216876 100722 216904 108990
rect 216784 100694 216904 100722
rect 216784 99414 216812 100694
rect 216772 99408 216824 99414
rect 216772 99350 216824 99356
rect 216680 91112 216732 91118
rect 216680 91054 216732 91060
rect 216692 72434 216720 91054
rect 216692 72406 216812 72434
rect 216784 60722 216812 72406
rect 216772 60716 216824 60722
rect 216772 60658 216824 60664
rect 216956 60716 217008 60722
rect 216956 60658 217008 60664
rect 216968 57934 216996 60658
rect 216956 57928 217008 57934
rect 216956 57870 217008 57876
rect 216864 48340 216916 48346
rect 216864 48282 216916 48288
rect 216876 43602 216904 48282
rect 216784 43574 216904 43602
rect 216784 38690 216812 43574
rect 216680 38684 216732 38690
rect 216680 38626 216732 38632
rect 216772 38684 216824 38690
rect 216772 38626 216824 38632
rect 216692 19378 216720 38626
rect 216680 19372 216732 19378
rect 216680 19314 216732 19320
rect 216956 19372 217008 19378
rect 216956 19314 217008 19320
rect 215392 5296 215444 5302
rect 215392 5238 215444 5244
rect 215852 4956 215904 4962
rect 215852 4898 215904 4904
rect 215300 4276 215352 4282
rect 215300 4218 215352 4224
rect 214656 3596 214708 3602
rect 214656 3538 214708 3544
rect 213472 598 213868 626
rect 213472 480 213500 598
rect 214668 480 214696 3538
rect 215864 480 215892 4898
rect 216968 2922 216996 19314
rect 217048 3324 217100 3330
rect 217048 3266 217100 3272
rect 216956 2916 217008 2922
rect 216956 2858 217008 2864
rect 217060 480 217088 3266
rect 217336 3058 217364 118594
rect 218060 113892 218112 113898
rect 218060 113834 218112 113840
rect 218072 4350 218100 113834
rect 218164 4486 218192 119734
rect 218440 113898 218468 120006
rect 218428 113892 218480 113898
rect 218428 113834 218480 113840
rect 219532 113892 219584 113898
rect 219532 113834 219584 113840
rect 219544 5370 219572 113834
rect 219532 5364 219584 5370
rect 219532 5306 219584 5312
rect 218152 4480 218204 4486
rect 218152 4422 218204 4428
rect 218060 4344 218112 4350
rect 218060 4286 218112 4292
rect 218152 3732 218204 3738
rect 218152 3674 218204 3680
rect 217324 3052 217376 3058
rect 217324 2994 217376 3000
rect 218164 480 218192 3674
rect 219636 3534 219664 120006
rect 219728 120006 219972 120034
rect 220280 120006 220616 120034
rect 220832 120006 221260 120034
rect 221660 120006 221812 120034
rect 222304 120006 222456 120034
rect 222672 120006 223008 120034
rect 219728 113898 219756 120006
rect 220084 118176 220136 118182
rect 220084 118118 220136 118124
rect 219716 113892 219768 113898
rect 219716 113834 219768 113840
rect 220096 3602 220124 118118
rect 220280 117570 220308 120006
rect 220268 117564 220320 117570
rect 220268 117506 220320 117512
rect 220084 3596 220136 3602
rect 220084 3538 220136 3544
rect 219624 3528 219676 3534
rect 219624 3470 219676 3476
rect 219348 3460 219400 3466
rect 219348 3402 219400 3408
rect 219360 480 219388 3402
rect 220544 3052 220596 3058
rect 220544 2994 220596 3000
rect 220556 480 220584 2994
rect 220832 2990 220860 120006
rect 221660 116006 221688 120006
rect 221464 116000 221516 116006
rect 221464 115942 221516 115948
rect 221648 116000 221700 116006
rect 221648 115942 221700 115948
rect 221476 109018 221504 115942
rect 222200 113892 222252 113898
rect 222200 113834 222252 113840
rect 221108 108990 221504 109018
rect 221108 100094 221136 108990
rect 221096 100088 221148 100094
rect 221096 100030 221148 100036
rect 221188 95260 221240 95266
rect 221188 95202 221240 95208
rect 221200 89706 221228 95202
rect 221108 89678 221228 89706
rect 221108 80170 221136 89678
rect 221096 80164 221148 80170
rect 221096 80106 221148 80112
rect 221004 79960 221056 79966
rect 221004 79902 221056 79908
rect 221016 72570 221044 79902
rect 221016 72542 221136 72570
rect 221108 72298 221136 72542
rect 221016 72270 221136 72298
rect 221016 70258 221044 72270
rect 221016 70230 221228 70258
rect 221200 60738 221228 70230
rect 221016 60722 221228 60738
rect 221004 60716 221240 60722
rect 221056 60710 221188 60716
rect 221004 60658 221056 60664
rect 221188 60658 221240 60664
rect 221200 51134 221228 60658
rect 221188 51128 221240 51134
rect 221188 51070 221240 51076
rect 221096 51060 221148 51066
rect 221096 51002 221148 51008
rect 221108 38690 221136 51002
rect 220912 38684 220964 38690
rect 220912 38626 220964 38632
rect 221096 38684 221148 38690
rect 221096 38626 221148 38632
rect 220924 24206 220952 38626
rect 220912 24200 220964 24206
rect 220912 24142 220964 24148
rect 221096 24200 221148 24206
rect 221096 24142 221148 24148
rect 221108 5438 221136 24142
rect 221096 5432 221148 5438
rect 221096 5374 221148 5380
rect 222212 3534 222240 113834
rect 222304 6254 222332 120006
rect 222672 113898 222700 120006
rect 223638 119762 223666 120020
rect 223960 120006 224296 120034
rect 224420 120006 224848 120034
rect 225156 120006 225492 120034
rect 225800 120006 226136 120034
rect 226444 120006 226688 120034
rect 226996 120006 227332 120034
rect 227732 120006 227976 120034
rect 228284 120006 228528 120034
rect 223638 119734 223712 119762
rect 222660 113892 222712 113898
rect 222660 113834 222712 113840
rect 222292 6248 222344 6254
rect 222292 6190 222344 6196
rect 223684 5506 223712 119734
rect 223960 117978 223988 120006
rect 223948 117972 224000 117978
rect 223948 117914 224000 117920
rect 224420 117722 224448 120006
rect 225156 118250 225184 120006
rect 225144 118244 225196 118250
rect 225144 118186 225196 118192
rect 225800 118114 225828 120006
rect 225788 118108 225840 118114
rect 225788 118050 225840 118056
rect 226248 117972 226300 117978
rect 226248 117914 226300 117920
rect 223776 117694 224448 117722
rect 223672 5500 223724 5506
rect 223672 5442 223724 5448
rect 222200 3528 222252 3534
rect 222200 3470 222252 3476
rect 222936 3528 222988 3534
rect 222936 3470 222988 3476
rect 220820 2984 220872 2990
rect 220820 2926 220872 2932
rect 221740 2984 221792 2990
rect 221740 2926 221792 2932
rect 221752 480 221780 2926
rect 222948 480 222976 3470
rect 223776 2922 223804 117694
rect 224224 117564 224276 117570
rect 224224 117506 224276 117512
rect 224236 3738 224264 117506
rect 225604 117360 225656 117366
rect 225604 117302 225656 117308
rect 225328 4140 225380 4146
rect 225328 4082 225380 4088
rect 224224 3732 224276 3738
rect 224224 3674 224276 3680
rect 224132 3596 224184 3602
rect 224132 3538 224184 3544
rect 223764 2916 223816 2922
rect 223764 2858 223816 2864
rect 224144 480 224172 3538
rect 225340 480 225368 4082
rect 225616 3194 225644 117302
rect 226260 4146 226288 117914
rect 226248 4140 226300 4146
rect 226248 4082 226300 4088
rect 226444 3874 226472 120006
rect 226996 117502 227024 120006
rect 227628 118108 227680 118114
rect 227628 118050 227680 118056
rect 226984 117496 227036 117502
rect 226984 117438 227036 117444
rect 227640 4146 227668 118050
rect 227732 118046 227760 120006
rect 227720 118040 227772 118046
rect 227720 117982 227772 117988
rect 228284 115977 228312 120006
rect 229158 119762 229186 120020
rect 229480 120006 229816 120034
rect 229940 120006 230368 120034
rect 230584 120006 231012 120034
rect 231320 120006 231656 120034
rect 231964 120006 232208 120034
rect 232516 120006 232852 120034
rect 233252 120006 233496 120034
rect 233620 120006 234048 120034
rect 229158 119734 229232 119762
rect 229204 118318 229232 119734
rect 229480 118454 229508 120006
rect 229468 118448 229520 118454
rect 229468 118390 229520 118396
rect 229192 118312 229244 118318
rect 229192 118254 229244 118260
rect 229008 118040 229060 118046
rect 229008 117982 229060 117988
rect 228364 117496 228416 117502
rect 228364 117438 228416 117444
rect 227994 115968 228050 115977
rect 227994 115903 228050 115912
rect 228270 115968 228326 115977
rect 228270 115903 228326 115912
rect 228008 109018 228036 115903
rect 227916 108990 228036 109018
rect 227916 101402 227944 108990
rect 227732 101374 227944 101402
rect 227732 96626 227760 101374
rect 227720 96620 227772 96626
rect 227720 96562 227772 96568
rect 227812 89684 227864 89690
rect 227812 89626 227864 89632
rect 227824 86986 227852 89626
rect 227824 86958 227944 86986
rect 227916 82142 227944 86958
rect 227904 82136 227956 82142
rect 227904 82078 227956 82084
rect 227996 77308 228048 77314
rect 227996 77250 228048 77256
rect 228008 60858 228036 77250
rect 227996 60852 228048 60858
rect 227996 60794 228048 60800
rect 227904 60784 227956 60790
rect 227904 60726 227956 60732
rect 227916 53174 227944 60726
rect 227904 53168 227956 53174
rect 227904 53110 227956 53116
rect 227996 48340 228048 48346
rect 227996 48282 228048 48288
rect 228008 22250 228036 48282
rect 227916 22222 228036 22250
rect 227916 22114 227944 22222
rect 227824 22086 227944 22114
rect 227824 21978 227852 22086
rect 227824 21950 227944 21978
rect 226524 4140 226576 4146
rect 226524 4082 226576 4088
rect 227628 4140 227680 4146
rect 227628 4082 227680 4088
rect 227720 4140 227772 4146
rect 227720 4082 227772 4088
rect 226432 3868 226484 3874
rect 226432 3810 226484 3816
rect 225604 3188 225656 3194
rect 225604 3130 225656 3136
rect 226536 480 226564 4082
rect 227732 480 227760 4082
rect 227916 3942 227944 21950
rect 227904 3936 227956 3942
rect 227904 3878 227956 3884
rect 228376 2990 228404 117438
rect 228914 19272 228970 19281
rect 228914 19207 228970 19216
rect 228928 9722 228956 19207
rect 228916 9716 228968 9722
rect 228916 9658 228968 9664
rect 229020 4146 229048 117982
rect 229940 117586 229968 120006
rect 230388 118448 230440 118454
rect 230388 118390 230440 118396
rect 229204 117558 229968 117586
rect 229204 99482 229232 117558
rect 229744 117428 229796 117434
rect 229744 117370 229796 117376
rect 229192 99476 229244 99482
rect 229192 99418 229244 99424
rect 229192 99340 229244 99346
rect 229192 99282 229244 99288
rect 229204 96642 229232 99282
rect 229204 96614 229324 96642
rect 229296 80170 229324 96614
rect 229284 80164 229336 80170
rect 229284 80106 229336 80112
rect 229192 80096 229244 80102
rect 229192 80038 229244 80044
rect 229204 70394 229232 80038
rect 229112 70366 229232 70394
rect 229112 70258 229140 70366
rect 229112 70230 229232 70258
rect 229204 51082 229232 70230
rect 229112 51054 229232 51082
rect 229112 50946 229140 51054
rect 229112 50918 229232 50946
rect 229204 31890 229232 50918
rect 229192 31884 229244 31890
rect 229192 31826 229244 31832
rect 229192 29028 229244 29034
rect 229192 28970 229244 28976
rect 229204 28914 229232 28970
rect 229204 28886 229324 28914
rect 229296 19378 229324 28886
rect 229100 19372 229152 19378
rect 229100 19314 229152 19320
rect 229284 19372 229336 19378
rect 229284 19314 229336 19320
rect 229112 19281 229140 19314
rect 229098 19272 229154 19281
rect 229098 19207 229154 19216
rect 229192 9716 229244 9722
rect 229192 9658 229244 9664
rect 229008 4140 229060 4146
rect 229008 4082 229060 4088
rect 228916 3868 228968 3874
rect 228916 3810 228968 3816
rect 228364 2984 228416 2990
rect 228364 2926 228416 2932
rect 228928 480 228956 3810
rect 229204 3738 229232 9658
rect 229192 3732 229244 3738
rect 229192 3674 229244 3680
rect 229756 3262 229784 117370
rect 229744 3256 229796 3262
rect 229744 3198 229796 3204
rect 230400 610 230428 118390
rect 230584 3806 230612 120006
rect 231320 118522 231348 120006
rect 231308 118516 231360 118522
rect 231308 118458 231360 118464
rect 231768 118312 231820 118318
rect 231768 118254 231820 118260
rect 231122 118008 231178 118017
rect 231122 117943 231178 117952
rect 230572 3800 230624 3806
rect 230572 3742 230624 3748
rect 231136 3126 231164 117943
rect 231780 4146 231808 118254
rect 231860 113892 231912 113898
rect 231860 113834 231912 113840
rect 231308 4140 231360 4146
rect 231308 4082 231360 4088
rect 231768 4140 231820 4146
rect 231768 4082 231820 4088
rect 231124 3120 231176 3126
rect 231124 3062 231176 3068
rect 230112 604 230164 610
rect 230112 546 230164 552
rect 230388 604 230440 610
rect 230388 546 230440 552
rect 230124 480 230152 546
rect 231320 480 231348 4082
rect 231872 3398 231900 113834
rect 231964 4010 231992 120006
rect 232412 117360 232464 117366
rect 232412 117302 232464 117308
rect 232424 113234 232452 117302
rect 232516 113898 232544 120006
rect 233252 118386 233280 120006
rect 233620 119354 233648 120006
rect 234678 119762 234706 120020
rect 233436 119326 233648 119354
rect 234632 119734 234706 119762
rect 235000 120006 235336 120034
rect 235460 120006 235888 120034
rect 236196 120006 236532 120034
rect 236840 120006 237176 120034
rect 237484 120006 237728 120034
rect 238036 120006 238372 120034
rect 238864 120006 239016 120034
rect 239324 120006 239568 120034
rect 233240 118380 233292 118386
rect 233240 118322 233292 118328
rect 233436 115938 233464 119326
rect 234632 118590 234660 119734
rect 234620 118584 234672 118590
rect 234620 118526 234672 118532
rect 234528 118380 234580 118386
rect 234528 118322 234580 118328
rect 233884 117836 233936 117842
rect 233884 117778 233936 117784
rect 233424 115932 233476 115938
rect 233424 115874 233476 115880
rect 233608 115932 233660 115938
rect 233608 115874 233660 115880
rect 232504 113892 232556 113898
rect 232504 113834 232556 113840
rect 232424 113206 232544 113234
rect 231952 4004 232004 4010
rect 231952 3946 232004 3952
rect 231860 3392 231912 3398
rect 231860 3334 231912 3340
rect 232516 3210 232544 113206
rect 233620 106321 233648 115874
rect 233422 106312 233478 106321
rect 233422 106247 233478 106256
rect 233606 106312 233662 106321
rect 233606 106247 233662 106256
rect 233436 104854 233464 106247
rect 233424 104848 233476 104854
rect 233424 104790 233476 104796
rect 233516 95260 233568 95266
rect 233516 95202 233568 95208
rect 233528 87038 233556 95202
rect 233424 87032 233476 87038
rect 233424 86974 233476 86980
rect 233516 87032 233568 87038
rect 233516 86974 233568 86980
rect 233436 86902 233464 86974
rect 233424 86896 233476 86902
rect 233424 86838 233476 86844
rect 233424 77308 233476 77314
rect 233424 77250 233476 77256
rect 233436 67590 233464 77250
rect 233424 67584 233476 67590
rect 233424 67526 233476 67532
rect 233424 62824 233476 62830
rect 233424 62766 233476 62772
rect 233436 41426 233464 62766
rect 233344 41398 233464 41426
rect 233344 41290 233372 41398
rect 233344 41262 233464 41290
rect 233436 29050 233464 41262
rect 233344 29022 233464 29050
rect 233344 22166 233372 29022
rect 233332 22160 233384 22166
rect 233332 22102 233384 22108
rect 233332 19304 233384 19310
rect 233332 19246 233384 19252
rect 233344 4622 233372 19246
rect 233332 4616 233384 4622
rect 233332 4558 233384 4564
rect 233700 4140 233752 4146
rect 233700 4082 233752 4088
rect 232424 3182 232544 3210
rect 232424 3058 232452 3182
rect 232504 3120 232556 3126
rect 232504 3062 232556 3068
rect 232412 3052 232464 3058
rect 232412 2994 232464 3000
rect 232516 480 232544 3062
rect 233712 480 233740 4082
rect 233896 3670 233924 117778
rect 234540 4146 234568 118322
rect 235000 117910 235028 120006
rect 234988 117904 235040 117910
rect 234988 117846 235040 117852
rect 235356 117904 235408 117910
rect 235356 117846 235408 117852
rect 235264 117428 235316 117434
rect 235264 117370 235316 117376
rect 234712 109064 234764 109070
rect 234712 109006 234764 109012
rect 234724 99482 234752 109006
rect 234712 99476 234764 99482
rect 234712 99418 234764 99424
rect 234712 99340 234764 99346
rect 234712 99282 234764 99288
rect 234724 67726 234752 99282
rect 234712 67720 234764 67726
rect 234712 67662 234764 67668
rect 234712 66292 234764 66298
rect 234712 66234 234764 66240
rect 234724 56574 234752 66234
rect 234712 56568 234764 56574
rect 234712 56510 234764 56516
rect 234712 46980 234764 46986
rect 234712 46922 234764 46928
rect 234724 37262 234752 46922
rect 234712 37256 234764 37262
rect 234712 37198 234764 37204
rect 234712 27668 234764 27674
rect 234712 27610 234764 27616
rect 234724 22846 234752 27610
rect 234712 22840 234764 22846
rect 234712 22782 234764 22788
rect 234620 18012 234672 18018
rect 234620 17954 234672 17960
rect 234632 9722 234660 17954
rect 234620 9716 234672 9722
rect 234620 9658 234672 9664
rect 234712 9716 234764 9722
rect 234712 9658 234764 9664
rect 234724 4554 234752 9658
rect 234712 4548 234764 4554
rect 234712 4490 234764 4496
rect 234528 4140 234580 4146
rect 234528 4082 234580 4088
rect 235276 3874 235304 117370
rect 235264 3868 235316 3874
rect 235264 3810 235316 3816
rect 233884 3664 233936 3670
rect 233884 3606 233936 3612
rect 234804 3664 234856 3670
rect 234804 3606 234856 3612
rect 234816 480 234844 3606
rect 235368 3126 235396 117846
rect 235460 109070 235488 120006
rect 236196 118454 236224 120006
rect 236184 118448 236236 118454
rect 236184 118390 236236 118396
rect 236840 118250 236868 120006
rect 236828 118244 236880 118250
rect 236828 118186 236880 118192
rect 237196 118244 237248 118250
rect 237196 118186 237248 118192
rect 235448 109064 235500 109070
rect 235448 109006 235500 109012
rect 236000 3936 236052 3942
rect 236000 3878 236052 3884
rect 235356 3120 235408 3126
rect 235356 3062 235408 3068
rect 236012 480 236040 3878
rect 237208 480 237236 118186
rect 237288 117292 237340 117298
rect 237288 117234 237340 117240
rect 237300 3942 237328 117234
rect 237484 5098 237512 120006
rect 238036 117638 238064 120006
rect 238668 118448 238720 118454
rect 238668 118390 238720 118396
rect 238024 117632 238076 117638
rect 238024 117574 238076 117580
rect 237472 5092 237524 5098
rect 237472 5034 237524 5040
rect 237288 3936 237340 3942
rect 237288 3878 237340 3884
rect 238680 610 238708 118390
rect 238864 117842 238892 120006
rect 238852 117836 238904 117842
rect 238852 117778 238904 117784
rect 239324 115977 239352 120006
rect 240198 119762 240226 120020
rect 240428 120006 240764 120034
rect 240888 120006 241408 120034
rect 241716 120006 242052 120034
rect 242268 120006 242604 120034
rect 243004 120006 243248 120034
rect 243556 120006 243892 120034
rect 244292 120006 244444 120034
rect 244660 120006 245088 120034
rect 240198 119734 240272 119762
rect 240244 118017 240272 119734
rect 240230 118008 240286 118017
rect 240230 117943 240286 117952
rect 240048 117836 240100 117842
rect 240048 117778 240100 117784
rect 238942 115968 238998 115977
rect 238942 115903 238998 115912
rect 239310 115968 239366 115977
rect 239310 115903 239366 115912
rect 238956 106350 238984 115903
rect 238852 106344 238904 106350
rect 238852 106286 238904 106292
rect 238944 106344 238996 106350
rect 238944 106286 238996 106292
rect 238864 101538 238892 106286
rect 238772 101510 238892 101538
rect 238772 96801 238800 101510
rect 238758 96792 238814 96801
rect 238758 96727 238814 96736
rect 238850 96656 238906 96665
rect 238850 96591 238852 96600
rect 238904 96591 238906 96600
rect 238852 96562 238904 96568
rect 238852 89684 238904 89690
rect 238852 89626 238904 89632
rect 238864 86986 238892 89626
rect 238864 86958 238984 86986
rect 238956 81462 238984 86958
rect 238944 81456 238996 81462
rect 238944 81398 238996 81404
rect 238944 77308 238996 77314
rect 238944 77250 238996 77256
rect 238956 60874 238984 77250
rect 238956 60846 239076 60874
rect 239048 53174 239076 60846
rect 238852 53168 238904 53174
rect 238852 53110 238904 53116
rect 239036 53168 239088 53174
rect 239036 53110 239088 53116
rect 238864 45898 238892 53110
rect 238852 45892 238904 45898
rect 238852 45834 238904 45840
rect 238944 41336 238996 41342
rect 238944 41278 238996 41284
rect 238956 37262 238984 41278
rect 238944 37256 238996 37262
rect 238944 37198 238996 37204
rect 238852 27668 238904 27674
rect 238852 27610 238904 27616
rect 238864 21978 238892 27610
rect 238864 21950 238984 21978
rect 238956 4826 238984 21950
rect 238944 4820 238996 4826
rect 238944 4762 238996 4768
rect 240060 4146 240088 117778
rect 240428 117774 240456 120006
rect 240888 119354 240916 120006
rect 240520 119326 240916 119354
rect 240416 117768 240468 117774
rect 240416 117710 240468 117716
rect 240520 113914 240548 119326
rect 241716 117706 241744 120006
rect 242268 118658 242296 120006
rect 242256 118652 242308 118658
rect 242256 118594 242308 118600
rect 241704 117700 241756 117706
rect 241704 117642 241756 117648
rect 241428 117360 241480 117366
rect 241428 117302 241480 117308
rect 240244 113886 240548 113914
rect 240244 99482 240272 113886
rect 240232 99476 240284 99482
rect 240232 99418 240284 99424
rect 240232 99340 240284 99346
rect 240232 99282 240284 99288
rect 240244 70514 240272 99282
rect 240232 70508 240284 70514
rect 240232 70450 240284 70456
rect 240232 67652 240284 67658
rect 240232 67594 240284 67600
rect 240244 58070 240272 67594
rect 240232 58064 240284 58070
rect 240232 58006 240284 58012
rect 240140 56636 240192 56642
rect 240140 56578 240192 56584
rect 240152 48346 240180 56578
rect 240140 48340 240192 48346
rect 240140 48282 240192 48288
rect 240232 48340 240284 48346
rect 240232 48282 240284 48288
rect 240244 12458 240272 48282
rect 240152 12430 240272 12458
rect 240152 4690 240180 12430
rect 240140 4684 240192 4690
rect 240140 4626 240192 4632
rect 239588 4140 239640 4146
rect 239588 4082 239640 4088
rect 240048 4140 240100 4146
rect 240048 4082 240100 4088
rect 238392 604 238444 610
rect 238392 546 238444 552
rect 238668 604 238720 610
rect 238668 546 238720 552
rect 238404 480 238432 546
rect 239600 480 239628 4082
rect 241440 3330 241468 117302
rect 243004 4894 243032 120006
rect 243556 117774 243584 120006
rect 244292 117978 244320 120006
rect 244660 119354 244688 120006
rect 245718 119762 245746 120020
rect 245948 120006 246284 120034
rect 246408 120006 246928 120034
rect 247236 120006 247572 120034
rect 247788 120006 248124 120034
rect 248616 120006 248768 120034
rect 249076 120006 249412 120034
rect 249812 120006 249964 120034
rect 250272 120006 250608 120034
rect 245718 119734 245792 119762
rect 244476 119326 244688 119354
rect 244280 117972 244332 117978
rect 244280 117914 244332 117920
rect 243544 117768 243596 117774
rect 243544 117710 243596 117716
rect 244188 117768 244240 117774
rect 244188 117710 244240 117716
rect 243636 117564 243688 117570
rect 243636 117506 243688 117512
rect 243542 117328 243598 117337
rect 243542 117263 243598 117272
rect 243452 53168 243504 53174
rect 243452 53110 243504 53116
rect 243464 48385 243492 53110
rect 243450 48376 243506 48385
rect 243450 48311 243506 48320
rect 243450 48240 243506 48249
rect 243450 48175 243506 48184
rect 243464 41886 243492 48175
rect 243452 41880 243504 41886
rect 243452 41822 243504 41828
rect 242992 4888 243044 4894
rect 242992 4830 243044 4836
rect 243176 4140 243228 4146
rect 243176 4082 243228 4088
rect 241980 4072 242032 4078
rect 241980 4014 242032 4020
rect 240784 3324 240836 3330
rect 240784 3266 240836 3272
rect 241428 3324 241480 3330
rect 241428 3266 241480 3272
rect 240796 480 240824 3266
rect 241992 480 242020 4014
rect 243188 480 243216 4082
rect 243556 3262 243584 117263
rect 243648 115938 243676 117506
rect 243636 115932 243688 115938
rect 243636 115874 243688 115880
rect 243912 115932 243964 115938
rect 243912 115874 243964 115880
rect 243924 114510 243952 115874
rect 243912 114504 243964 114510
rect 243912 114446 243964 114452
rect 243728 104916 243780 104922
rect 243728 104858 243780 104864
rect 243740 104802 243768 104858
rect 243648 104774 243768 104802
rect 243648 99414 243676 104774
rect 243636 99408 243688 99414
rect 243636 99350 243688 99356
rect 243728 95260 243780 95266
rect 243728 95202 243780 95208
rect 243740 89758 243768 95202
rect 243728 89752 243780 89758
rect 243728 89694 243780 89700
rect 243728 89616 243780 89622
rect 243728 89558 243780 89564
rect 243740 86970 243768 89558
rect 243728 86964 243780 86970
rect 243728 86906 243780 86912
rect 243728 77308 243780 77314
rect 243728 77250 243780 77256
rect 243740 60858 243768 77250
rect 243728 60852 243780 60858
rect 243728 60794 243780 60800
rect 243728 60648 243780 60654
rect 243728 60590 243780 60596
rect 243740 53174 243768 60590
rect 243728 53168 243780 53174
rect 243728 53110 243780 53116
rect 243820 41880 243872 41886
rect 243820 41822 243872 41828
rect 243832 35850 243860 41822
rect 243740 35822 243860 35850
rect 243740 27674 243768 35822
rect 243728 27668 243780 27674
rect 243728 27610 243780 27616
rect 243728 26308 243780 26314
rect 243728 26250 243780 26256
rect 243740 22166 243768 26250
rect 243728 22160 243780 22166
rect 243728 22102 243780 22108
rect 243728 22024 243780 22030
rect 243728 21966 243780 21972
rect 243740 4078 243768 21966
rect 244200 4146 244228 117710
rect 244476 106298 244504 119326
rect 245476 118040 245528 118046
rect 245476 117982 245528 117988
rect 244476 106270 244596 106298
rect 244568 99414 244596 106270
rect 244372 99408 244424 99414
rect 244372 99350 244424 99356
rect 244556 99408 244608 99414
rect 244556 99350 244608 99356
rect 244384 91746 244412 99350
rect 244292 91718 244412 91746
rect 244292 75886 244320 91718
rect 244280 75880 244332 75886
rect 244280 75822 244332 75828
rect 244372 66292 244424 66298
rect 244372 66234 244424 66240
rect 244384 60722 244412 66234
rect 244372 60716 244424 60722
rect 244372 60658 244424 60664
rect 244556 60716 244608 60722
rect 244556 60658 244608 60664
rect 244568 51134 244596 60658
rect 244556 51128 244608 51134
rect 244556 51070 244608 51076
rect 244464 51060 244516 51066
rect 244464 51002 244516 51008
rect 244476 41834 244504 51002
rect 244384 41806 244504 41834
rect 244384 38690 244412 41806
rect 244280 38684 244332 38690
rect 244280 38626 244332 38632
rect 244372 38684 244424 38690
rect 244372 38626 244424 38632
rect 244292 37262 244320 38626
rect 244280 37256 244332 37262
rect 244280 37198 244332 37204
rect 244372 31680 244424 31686
rect 244372 31622 244424 31628
rect 244384 22098 244412 31622
rect 244372 22092 244424 22098
rect 244372 22034 244424 22040
rect 244556 22092 244608 22098
rect 244556 22034 244608 22040
rect 244568 19310 244596 22034
rect 244556 19304 244608 19310
rect 244556 19246 244608 19252
rect 244556 11892 244608 11898
rect 244556 11834 244608 11840
rect 244568 4962 244596 11834
rect 244556 4956 244608 4962
rect 244556 4898 244608 4904
rect 244188 4140 244240 4146
rect 244188 4082 244240 4088
rect 244372 4140 244424 4146
rect 244372 4082 244424 4088
rect 243728 4072 243780 4078
rect 243728 4014 243780 4020
rect 243544 3256 243596 3262
rect 243544 3198 243596 3204
rect 244384 480 244412 4082
rect 245488 4026 245516 117982
rect 245568 117700 245620 117706
rect 245568 117642 245620 117648
rect 245580 4146 245608 117642
rect 245764 117337 245792 119734
rect 245948 117502 245976 120006
rect 246408 119354 246436 120006
rect 246040 119326 246436 119354
rect 245936 117496 245988 117502
rect 245936 117438 245988 117444
rect 245750 117328 245806 117337
rect 245750 117263 245806 117272
rect 246040 109154 246068 119326
rect 247236 118114 247264 120006
rect 247224 118108 247276 118114
rect 247224 118050 247276 118056
rect 247684 117632 247736 117638
rect 247684 117574 247736 117580
rect 246040 109126 246160 109154
rect 246132 108882 246160 109126
rect 246040 108854 246160 108882
rect 246040 99414 246068 108854
rect 245844 99408 245896 99414
rect 245844 99350 245896 99356
rect 246028 99408 246080 99414
rect 246028 99350 246080 99356
rect 245856 89434 245884 99350
rect 245856 89406 245976 89434
rect 245948 86970 245976 89406
rect 245936 86964 245988 86970
rect 245936 86906 245988 86912
rect 245752 77308 245804 77314
rect 245752 77250 245804 77256
rect 245764 75886 245792 77250
rect 245752 75880 245804 75886
rect 245752 75822 245804 75828
rect 245844 66292 245896 66298
rect 245844 66234 245896 66240
rect 245856 60722 245884 66234
rect 245844 60716 245896 60722
rect 245844 60658 245896 60664
rect 246028 60716 246080 60722
rect 246028 60658 246080 60664
rect 246040 51082 246068 60658
rect 245948 51054 246068 51082
rect 245948 43738 245976 51054
rect 245856 43710 245976 43738
rect 245856 38690 245884 43710
rect 245752 38684 245804 38690
rect 245752 38626 245804 38632
rect 245844 38684 245896 38690
rect 245844 38626 245896 38632
rect 245764 37262 245792 38626
rect 245752 37256 245804 37262
rect 245752 37198 245804 37204
rect 245844 31748 245896 31754
rect 245844 31690 245896 31696
rect 245856 22098 245884 31690
rect 245844 22092 245896 22098
rect 245844 22034 245896 22040
rect 246028 22092 246080 22098
rect 246028 22034 246080 22040
rect 246040 11966 246068 22034
rect 246028 11960 246080 11966
rect 246028 11902 246080 11908
rect 246028 11824 246080 11830
rect 246028 11766 246080 11772
rect 245568 4140 245620 4146
rect 245568 4082 245620 4088
rect 245488 3998 245608 4026
rect 245580 480 245608 3998
rect 246040 3466 246068 11766
rect 247696 4146 247724 117574
rect 247788 117570 247816 120006
rect 247776 117564 247828 117570
rect 247776 117506 247828 117512
rect 248328 117496 248380 117502
rect 248328 117438 248380 117444
rect 248340 115938 248368 117438
rect 248328 115932 248380 115938
rect 248328 115874 248380 115880
rect 248512 113892 248564 113898
rect 248512 113834 248564 113840
rect 248328 106344 248380 106350
rect 248328 106286 248380 106292
rect 248340 104854 248368 106286
rect 248328 104848 248380 104854
rect 248328 104790 248380 104796
rect 248236 95260 248288 95266
rect 248236 95202 248288 95208
rect 248248 87174 248276 95202
rect 248236 87168 248288 87174
rect 248236 87110 248288 87116
rect 248328 87032 248380 87038
rect 248328 86974 248380 86980
rect 248340 85542 248368 86974
rect 248328 85536 248380 85542
rect 248328 85478 248380 85484
rect 248328 75948 248380 75954
rect 248328 75890 248380 75896
rect 248340 66230 248368 75890
rect 248328 66224 248380 66230
rect 248328 66166 248380 66172
rect 248328 56636 248380 56642
rect 248328 56578 248380 56584
rect 248340 48346 248368 56578
rect 248328 48340 248380 48346
rect 248328 48282 248380 48288
rect 248328 46980 248380 46986
rect 248328 46922 248380 46928
rect 248340 37262 248368 46922
rect 248328 37256 248380 37262
rect 248328 37198 248380 37204
rect 248328 27668 248380 27674
rect 248328 27610 248380 27616
rect 248340 8362 248368 27610
rect 247960 8356 248012 8362
rect 247960 8298 248012 8304
rect 248328 8356 248380 8362
rect 248328 8298 248380 8304
rect 246764 4140 246816 4146
rect 246764 4082 246816 4088
rect 247684 4140 247736 4146
rect 247684 4082 247736 4088
rect 246028 3460 246080 3466
rect 246028 3402 246080 3408
rect 246776 480 246804 4082
rect 247972 480 248000 8298
rect 248524 3602 248552 113834
rect 248512 3596 248564 3602
rect 248512 3538 248564 3544
rect 248616 3534 248644 120006
rect 248970 118144 249026 118153
rect 248970 118079 249026 118088
rect 248984 117842 249012 118079
rect 248972 117836 249024 117842
rect 248972 117778 249024 117784
rect 249076 113898 249104 120006
rect 249812 118318 249840 120006
rect 249800 118312 249852 118318
rect 249800 118254 249852 118260
rect 250272 118114 250300 120006
rect 251238 119762 251266 120020
rect 251468 120006 251804 120034
rect 252112 120006 252448 120034
rect 252756 120006 253092 120034
rect 253308 120006 253644 120034
rect 253952 120006 254288 120034
rect 254596 120006 254932 120034
rect 255332 120006 255484 120034
rect 255792 120006 256128 120034
rect 251238 119734 251312 119762
rect 250260 118108 250312 118114
rect 250260 118050 250312 118056
rect 251088 117972 251140 117978
rect 251088 117914 251140 117920
rect 249708 117564 249760 117570
rect 249708 117506 249760 117512
rect 249064 113892 249116 113898
rect 249064 113834 249116 113840
rect 249720 4146 249748 117506
rect 250444 117360 250496 117366
rect 250444 117302 250496 117308
rect 249156 4140 249208 4146
rect 249156 4082 249208 4088
rect 249708 4140 249760 4146
rect 249708 4082 249760 4088
rect 248604 3528 248656 3534
rect 248604 3470 248656 3476
rect 249168 480 249196 4082
rect 250456 3670 250484 117302
rect 250444 3664 250496 3670
rect 250444 3606 250496 3612
rect 251100 3398 251128 117914
rect 251284 117842 251312 119734
rect 251468 118318 251496 120006
rect 251456 118312 251508 118318
rect 251456 118254 251508 118260
rect 251548 118312 251600 118318
rect 251548 118254 251600 118260
rect 251560 118153 251588 118254
rect 251546 118144 251602 118153
rect 251546 118079 251602 118088
rect 252112 118046 252140 120006
rect 252756 118590 252784 120006
rect 252744 118584 252796 118590
rect 252744 118526 252796 118532
rect 252468 118108 252520 118114
rect 252468 118050 252520 118056
rect 252100 118040 252152 118046
rect 252100 117982 252152 117988
rect 251272 117836 251324 117842
rect 251272 117778 251324 117784
rect 252480 4146 252508 118050
rect 253308 117434 253336 120006
rect 253952 118386 253980 120006
rect 253940 118380 253992 118386
rect 253940 118322 253992 118328
rect 253296 117428 253348 117434
rect 253296 117370 253348 117376
rect 254596 117366 254624 120006
rect 255332 118522 255360 120006
rect 255320 118516 255372 118522
rect 255320 118458 255372 118464
rect 255792 118454 255820 120006
rect 256758 119762 256786 120020
rect 256712 119734 256786 119762
rect 256988 120006 257324 120034
rect 257632 120006 257968 120034
rect 258276 120006 258520 120034
rect 258828 120006 259164 120034
rect 259472 120006 259808 120034
rect 260024 120006 260360 120034
rect 260852 120006 261004 120034
rect 261312 120006 261648 120034
rect 255780 118448 255832 118454
rect 255780 118390 255832 118396
rect 256608 118380 256660 118386
rect 256608 118322 256660 118328
rect 254676 118244 254728 118250
rect 254676 118186 254728 118192
rect 254584 117360 254636 117366
rect 254584 117302 254636 117308
rect 254688 115682 254716 118186
rect 255228 118040 255280 118046
rect 255228 117982 255280 117988
rect 254596 115654 254716 115682
rect 251456 4140 251508 4146
rect 251456 4082 251508 4088
rect 252468 4140 252520 4146
rect 252468 4082 252520 4088
rect 250352 3392 250404 3398
rect 250352 3334 250404 3340
rect 251088 3392 251140 3398
rect 251088 3334 251140 3340
rect 250364 480 250392 3334
rect 251468 480 251496 4082
rect 253848 3324 253900 3330
rect 253848 3266 253900 3272
rect 252652 3052 252704 3058
rect 252652 2994 252704 3000
rect 252664 480 252692 2994
rect 253860 480 253888 3266
rect 254596 3058 254624 115654
rect 255240 3346 255268 117982
rect 256620 3346 256648 118322
rect 256712 117910 256740 119734
rect 256988 118318 257016 120006
rect 257632 118590 257660 120006
rect 258276 118658 258304 120006
rect 258264 118652 258316 118658
rect 258264 118594 258316 118600
rect 257620 118584 257672 118590
rect 257620 118526 257672 118532
rect 257344 118516 257396 118522
rect 257344 118458 257396 118464
rect 256976 118312 257028 118318
rect 256976 118254 257028 118260
rect 256700 117904 256752 117910
rect 256700 117846 256752 117852
rect 255056 3318 255268 3346
rect 256252 3318 256648 3346
rect 257356 3330 257384 118458
rect 257988 118312 258040 118318
rect 257988 118254 258040 118260
rect 258000 3534 258028 118254
rect 258828 117774 258856 120006
rect 258816 117768 258868 117774
rect 258816 117710 258868 117716
rect 259472 117706 259500 120006
rect 260024 118182 260052 120006
rect 260012 118176 260064 118182
rect 260012 118118 260064 118124
rect 259460 117700 259512 117706
rect 259460 117642 259512 117648
rect 260852 117638 260880 120006
rect 260840 117632 260892 117638
rect 260840 117574 260892 117580
rect 261312 117502 261340 120006
rect 262186 119762 262214 120020
rect 262508 120006 262844 120034
rect 263152 120006 263488 120034
rect 263704 120006 264040 120034
rect 264348 120006 264684 120034
rect 264992 120006 265328 120034
rect 265544 120006 265880 120034
rect 266372 120006 266524 120034
rect 266832 120006 267168 120034
rect 262186 119734 262260 119762
rect 262128 117904 262180 117910
rect 262128 117846 262180 117852
rect 261300 117496 261352 117502
rect 261300 117438 261352 117444
rect 261484 117428 261536 117434
rect 261484 117370 261536 117376
rect 259368 117360 259420 117366
rect 259368 117302 259420 117308
rect 257436 3528 257488 3534
rect 257436 3470 257488 3476
rect 257988 3528 258040 3534
rect 257988 3470 258040 3476
rect 257344 3324 257396 3330
rect 254584 3052 254636 3058
rect 254584 2994 254636 3000
rect 255056 480 255084 3318
rect 256252 480 256280 3318
rect 257344 3266 257396 3272
rect 257448 480 257476 3470
rect 259380 3126 259408 117302
rect 261496 3534 261524 117370
rect 259828 3528 259880 3534
rect 259828 3470 259880 3476
rect 261484 3528 261536 3534
rect 261484 3470 261536 3476
rect 258632 3120 258684 3126
rect 258632 3062 258684 3068
rect 259368 3120 259420 3126
rect 259368 3062 259420 3068
rect 258644 480 258672 3062
rect 259840 480 259868 3470
rect 262140 3262 262168 117846
rect 262232 117570 262260 119734
rect 262508 117978 262536 120006
rect 263152 118114 263180 120006
rect 263704 118250 263732 120006
rect 264348 118522 264376 120006
rect 264336 118516 264388 118522
rect 264336 118458 264388 118464
rect 263692 118244 263744 118250
rect 263692 118186 263744 118192
rect 263140 118108 263192 118114
rect 263140 118050 263192 118056
rect 263416 118108 263468 118114
rect 263416 118050 263468 118056
rect 262496 117972 262548 117978
rect 262496 117914 262548 117920
rect 262220 117564 262272 117570
rect 262220 117506 262272 117512
rect 262220 3528 262272 3534
rect 262220 3470 262272 3476
rect 261024 3256 261076 3262
rect 261024 3198 261076 3204
rect 262128 3256 262180 3262
rect 262128 3198 262180 3204
rect 261036 480 261064 3198
rect 262232 480 262260 3470
rect 263428 480 263456 118050
rect 264992 118046 265020 120006
rect 265544 118386 265572 120006
rect 265532 118380 265584 118386
rect 265532 118322 265584 118328
rect 266372 118318 266400 120006
rect 266360 118312 266412 118318
rect 266360 118254 266412 118260
rect 264980 118040 265032 118046
rect 264980 117982 265032 117988
rect 263508 117972 263560 117978
rect 263508 117914 263560 117920
rect 263520 3534 263548 117914
rect 266268 117564 266320 117570
rect 266268 117506 266320 117512
rect 266280 4146 266308 117506
rect 266832 117366 266860 120006
rect 267706 119762 267734 120020
rect 268028 120006 268364 120034
rect 268672 120006 269008 120034
rect 269224 120006 269560 120034
rect 269868 120006 270204 120034
rect 270512 120006 270848 120034
rect 271064 120006 271400 120034
rect 271892 120006 272044 120034
rect 272444 120006 272688 120034
rect 273240 120006 273392 120034
rect 267706 119734 267780 119762
rect 267648 117496 267700 117502
rect 267648 117438 267700 117444
rect 266820 117360 266872 117366
rect 266820 117302 266872 117308
rect 265808 4140 265860 4146
rect 265808 4082 265860 4088
rect 266268 4140 266320 4146
rect 266268 4082 266320 4088
rect 263508 3528 263560 3534
rect 263508 3470 263560 3476
rect 264612 3120 264664 3126
rect 264612 3062 264664 3068
rect 264624 480 264652 3062
rect 265820 480 265848 4082
rect 267660 3330 267688 117438
rect 267752 117434 267780 119734
rect 268028 117910 268056 120006
rect 268672 117978 268700 120006
rect 269224 118114 269252 120006
rect 269212 118108 269264 118114
rect 269212 118050 269264 118056
rect 268660 117972 268712 117978
rect 268660 117914 268712 117920
rect 268016 117904 268068 117910
rect 268016 117846 268068 117852
rect 267740 117428 267792 117434
rect 267740 117370 267792 117376
rect 269764 117428 269816 117434
rect 269764 117370 269816 117376
rect 268384 117360 268436 117366
rect 268384 117302 268436 117308
rect 268108 4140 268160 4146
rect 268108 4082 268160 4088
rect 267004 3324 267056 3330
rect 267004 3266 267056 3272
rect 267648 3324 267700 3330
rect 267648 3266 267700 3272
rect 267016 480 267044 3266
rect 268120 480 268148 4082
rect 268396 3126 268424 117302
rect 269776 4146 269804 117370
rect 269868 117366 269896 120006
rect 270512 117570 270540 120006
rect 270500 117564 270552 117570
rect 270500 117506 270552 117512
rect 271064 117502 271092 120006
rect 271052 117496 271104 117502
rect 271052 117438 271104 117444
rect 271892 117434 271920 120006
rect 271880 117428 271932 117434
rect 271880 117370 271932 117376
rect 269856 117360 269908 117366
rect 269856 117302 269908 117308
rect 272444 116006 272472 120006
rect 272524 117428 272576 117434
rect 272524 117370 272576 117376
rect 272248 116000 272300 116006
rect 272248 115942 272300 115948
rect 272432 116000 272484 116006
rect 272432 115942 272484 115948
rect 272260 114510 272288 115942
rect 272248 114504 272300 114510
rect 272248 114446 272300 114452
rect 272064 103556 272116 103562
rect 272064 103498 272116 103504
rect 272076 99482 272104 103498
rect 272064 99476 272116 99482
rect 272064 99418 272116 99424
rect 271972 99340 272024 99346
rect 271972 99282 272024 99288
rect 271984 90386 272012 99282
rect 271892 90358 272012 90386
rect 271892 87038 271920 90358
rect 271880 87032 271932 87038
rect 271880 86974 271932 86980
rect 271880 86896 271932 86902
rect 271880 86838 271932 86844
rect 271892 80322 271920 86838
rect 271892 80294 272012 80322
rect 271984 80050 272012 80294
rect 271892 80022 272012 80050
rect 271892 75886 271920 80022
rect 271880 75880 271932 75886
rect 271880 75822 271932 75828
rect 271972 70304 272024 70310
rect 271972 70246 272024 70252
rect 271984 60722 272012 70246
rect 271972 60716 272024 60722
rect 271972 60658 272024 60664
rect 272156 60716 272208 60722
rect 272156 60658 272208 60664
rect 272168 51134 272196 60658
rect 272156 51128 272208 51134
rect 272156 51070 272208 51076
rect 272064 51060 272116 51066
rect 272064 51002 272116 51008
rect 272076 43466 272104 51002
rect 271892 43438 272104 43466
rect 271892 37262 271920 43438
rect 271880 37256 271932 37262
rect 271880 37198 271932 37204
rect 272156 27668 272208 27674
rect 272156 27610 272208 27616
rect 269764 4140 269816 4146
rect 269764 4082 269816 4088
rect 271696 4140 271748 4146
rect 271696 4082 271748 4088
rect 269304 4004 269356 4010
rect 269304 3946 269356 3952
rect 268384 3120 268436 3126
rect 268384 3062 268436 3068
rect 269316 480 269344 3946
rect 270500 3460 270552 3466
rect 270500 3402 270552 3408
rect 270512 480 270540 3402
rect 271708 480 271736 4082
rect 272168 4010 272196 27610
rect 272536 4146 272564 117370
rect 273168 117360 273220 117366
rect 273168 117302 273220 117308
rect 272524 4140 272576 4146
rect 272524 4082 272576 4088
rect 272156 4004 272208 4010
rect 272156 3946 272208 3952
rect 273180 610 273208 117302
rect 273364 3466 273392 120006
rect 273548 120006 273884 120034
rect 274192 120006 274528 120034
rect 274652 120006 275080 120034
rect 275388 120006 275724 120034
rect 276124 120006 276276 120034
rect 276920 120006 277348 120034
rect 277564 120006 277900 120034
rect 278116 120006 278452 120034
rect 278760 120006 279096 120034
rect 279404 120006 279740 120034
rect 279956 120006 280108 120034
rect 280600 120006 280936 120034
rect 281244 120006 281488 120034
rect 281796 120006 282132 120034
rect 282440 120006 282776 120034
rect 283084 120006 283420 120034
rect 283636 120006 283972 120034
rect 284280 120006 284616 120034
rect 284924 120006 285260 120034
rect 273548 117434 273576 120006
rect 273536 117428 273588 117434
rect 273536 117370 273588 117376
rect 274192 117366 274220 120006
rect 274180 117360 274232 117366
rect 274652 117314 274680 120006
rect 274180 117302 274232 117308
rect 274560 117286 274680 117314
rect 274560 4146 274588 117286
rect 275388 104922 275416 120006
rect 274916 104916 274968 104922
rect 274916 104858 274968 104864
rect 275376 104916 275428 104922
rect 275376 104858 275428 104864
rect 274928 100042 274956 104858
rect 274744 100014 274956 100042
rect 274744 89706 274772 100014
rect 274744 89678 274956 89706
rect 274928 86970 274956 89678
rect 274916 86964 274968 86970
rect 274916 86906 274968 86912
rect 274824 77308 274876 77314
rect 274824 77250 274876 77256
rect 274836 18154 274864 77250
rect 276124 57934 276152 120006
rect 276112 57928 276164 57934
rect 276112 57870 276164 57876
rect 276296 57928 276348 57934
rect 276296 57870 276348 57876
rect 276308 48385 276336 57870
rect 276110 48376 276166 48385
rect 276110 48311 276166 48320
rect 276294 48376 276350 48385
rect 276294 48311 276350 48320
rect 276124 46918 276152 48311
rect 276112 46912 276164 46918
rect 276112 46854 276164 46860
rect 276112 37324 276164 37330
rect 276112 37266 276164 37272
rect 276124 27606 276152 37266
rect 276112 27600 276164 27606
rect 276112 27542 276164 27548
rect 274824 18148 274876 18154
rect 274824 18090 274876 18096
rect 276112 18012 276164 18018
rect 276112 17954 276164 17960
rect 276124 12510 276152 17954
rect 276112 12504 276164 12510
rect 276112 12446 276164 12452
rect 276480 12368 276532 12374
rect 276480 12310 276532 12316
rect 275284 9716 275336 9722
rect 275284 9658 275336 9664
rect 274088 4140 274140 4146
rect 274088 4082 274140 4088
rect 274548 4140 274600 4146
rect 274548 4082 274600 4088
rect 273352 3460 273404 3466
rect 273352 3402 273404 3408
rect 272892 604 272944 610
rect 272892 546 272944 552
rect 273168 604 273220 610
rect 273168 546 273220 552
rect 272904 480 272932 546
rect 274100 480 274128 4082
rect 275296 480 275324 9658
rect 276492 480 276520 12310
rect 277320 4146 277348 120006
rect 277872 117366 277900 120006
rect 278424 117434 278452 120006
rect 278412 117428 278464 117434
rect 278412 117370 278464 117376
rect 279068 117366 279096 120006
rect 279712 119354 279740 120006
rect 279712 119326 280016 119354
rect 279148 117428 279200 117434
rect 279148 117370 279200 117376
rect 277860 117360 277912 117366
rect 277860 117302 277912 117308
rect 278872 117360 278924 117366
rect 278872 117302 278924 117308
rect 279056 117360 279108 117366
rect 279056 117302 279108 117308
rect 277308 4140 277360 4146
rect 277308 4082 277360 4088
rect 277676 4140 277728 4146
rect 277676 4082 277728 4088
rect 277688 480 277716 4082
rect 278884 480 278912 117302
rect 279160 4026 279188 117370
rect 279988 109018 280016 119326
rect 280080 117570 280108 120006
rect 280068 117564 280120 117570
rect 280068 117506 280120 117512
rect 280908 117366 280936 120006
rect 280344 117360 280396 117366
rect 280344 117302 280396 117308
rect 280896 117360 280948 117366
rect 280896 117302 280948 117308
rect 281356 117360 281408 117366
rect 281356 117302 281408 117308
rect 279804 108990 280016 109018
rect 279804 103494 279832 108990
rect 279792 103488 279844 103494
rect 279792 103430 279844 103436
rect 279976 103488 280028 103494
rect 279976 103430 280028 103436
rect 279988 93945 280016 103430
rect 279790 93936 279846 93945
rect 279712 93894 279790 93922
rect 279712 93838 279740 93894
rect 279790 93871 279846 93880
rect 279974 93936 280030 93945
rect 279974 93871 280030 93880
rect 279700 93832 279752 93838
rect 279700 93774 279752 93780
rect 279700 84312 279752 84318
rect 279700 84254 279752 84260
rect 279712 84182 279740 84254
rect 279700 84176 279752 84182
rect 279700 84118 279752 84124
rect 279792 74588 279844 74594
rect 279792 74530 279844 74536
rect 279804 70446 279832 74530
rect 279792 70440 279844 70446
rect 279792 70382 279844 70388
rect 279792 70304 279844 70310
rect 279792 70246 279844 70252
rect 279804 60738 279832 70246
rect 279804 60722 279924 60738
rect 279804 60716 279936 60722
rect 279804 60710 279884 60716
rect 279884 60658 279936 60664
rect 280068 60716 280120 60722
rect 280068 60658 280120 60664
rect 280080 57934 280108 60658
rect 280068 57928 280120 57934
rect 280068 57870 280120 57876
rect 279884 48340 279936 48346
rect 279884 48282 279936 48288
rect 279896 31754 279924 48282
rect 279884 31748 279936 31754
rect 279884 31690 279936 31696
rect 280068 31748 280120 31754
rect 280068 31690 280120 31696
rect 280080 28966 280108 31690
rect 280068 28960 280120 28966
rect 280068 28902 280120 28908
rect 279976 19372 280028 19378
rect 279976 19314 280028 19320
rect 279988 12458 280016 19314
rect 279988 12430 280108 12458
rect 280356 12442 280384 117302
rect 280080 4146 280108 12430
rect 280344 12436 280396 12442
rect 280344 12378 280396 12384
rect 281264 12436 281316 12442
rect 281264 12378 281316 12384
rect 280068 4140 280120 4146
rect 280068 4082 280120 4088
rect 279160 3998 280108 4026
rect 280080 480 280108 3998
rect 281276 480 281304 12378
rect 281368 3194 281396 117302
rect 281460 3262 281488 120006
rect 282104 117434 282132 120006
rect 282748 117502 282776 120006
rect 283104 117564 283156 117570
rect 283104 117506 283156 117512
rect 282736 117496 282788 117502
rect 282736 117438 282788 117444
rect 282092 117428 282144 117434
rect 282092 117370 282144 117376
rect 282460 4140 282512 4146
rect 282460 4082 282512 4088
rect 281448 3256 281500 3262
rect 281448 3198 281500 3204
rect 281356 3188 281408 3194
rect 281356 3130 281408 3136
rect 282472 480 282500 4082
rect 283116 3346 283144 117506
rect 283392 117366 283420 120006
rect 283944 118046 283972 120006
rect 284588 118114 284616 120006
rect 284576 118108 284628 118114
rect 284576 118050 284628 118056
rect 283932 118040 283984 118046
rect 283932 117982 283984 117988
rect 284944 117496 284996 117502
rect 284944 117438 284996 117444
rect 283564 117428 283616 117434
rect 283564 117370 283616 117376
rect 283380 117360 283432 117366
rect 283380 117302 283432 117308
rect 283576 3942 283604 117370
rect 284208 117360 284260 117366
rect 284208 117302 284260 117308
rect 284220 4078 284248 117302
rect 284208 4072 284260 4078
rect 284208 4014 284260 4020
rect 283564 3936 283616 3942
rect 283564 3878 283616 3884
rect 284956 3670 284984 117438
rect 285232 117366 285260 120006
rect 285462 119762 285490 120020
rect 286120 120006 286456 120034
rect 286764 120006 287008 120034
rect 287316 120006 287652 120034
rect 287960 120006 288296 120034
rect 288604 120006 288940 120034
rect 289156 120006 289492 120034
rect 289800 120006 290044 120034
rect 290444 120006 290780 120034
rect 285462 119734 285536 119762
rect 285220 117360 285272 117366
rect 285220 117302 285272 117308
rect 284944 3664 284996 3670
rect 284944 3606 284996 3612
rect 285508 3466 285536 119734
rect 286428 117366 286456 120006
rect 285588 117360 285640 117366
rect 285588 117302 285640 117308
rect 286416 117360 286468 117366
rect 286416 117302 286468 117308
rect 286876 117360 286928 117366
rect 286876 117302 286928 117308
rect 285600 4010 285628 117302
rect 285588 4004 285640 4010
rect 285588 3946 285640 3952
rect 286888 3874 286916 117302
rect 286876 3868 286928 3874
rect 286876 3810 286928 3816
rect 286980 3806 287008 120006
rect 287624 117366 287652 120006
rect 287612 117360 287664 117366
rect 287612 117302 287664 117308
rect 287152 3936 287204 3942
rect 287152 3878 287204 3884
rect 286968 3800 287020 3806
rect 286968 3742 287020 3748
rect 285496 3460 285548 3466
rect 285496 3402 285548 3408
rect 283116 3318 283696 3346
rect 283668 480 283696 3318
rect 285956 3256 286008 3262
rect 285956 3198 286008 3204
rect 284760 3188 284812 3194
rect 284760 3130 284812 3136
rect 284772 480 284800 3130
rect 285968 480 285996 3198
rect 287164 480 287192 3878
rect 288268 3738 288296 120006
rect 288912 117910 288940 120006
rect 288900 117904 288952 117910
rect 288900 117846 288952 117852
rect 289464 117502 289492 120006
rect 289452 117496 289504 117502
rect 289452 117438 289504 117444
rect 290016 117434 290044 120006
rect 290096 118040 290148 118046
rect 290096 117982 290148 117988
rect 290004 117428 290056 117434
rect 290004 117370 290056 117376
rect 288348 117360 288400 117366
rect 288348 117302 288400 117308
rect 288360 3942 288388 117302
rect 289544 4072 289596 4078
rect 289544 4014 289596 4020
rect 288348 3936 288400 3942
rect 288348 3878 288400 3884
rect 288256 3732 288308 3738
rect 288256 3674 288308 3680
rect 288348 3664 288400 3670
rect 288348 3606 288400 3612
rect 288360 480 288388 3606
rect 289556 480 289584 4014
rect 290108 610 290136 117982
rect 290752 117366 290780 120006
rect 290982 119762 291010 120020
rect 291640 120006 291976 120034
rect 292284 120006 292436 120034
rect 292836 120006 293172 120034
rect 293480 120006 293816 120034
rect 294032 120006 294368 120034
rect 294676 120006 295012 120034
rect 295320 120006 295656 120034
rect 295872 120006 296208 120034
rect 296516 120006 296668 120034
rect 297160 120006 297496 120034
rect 297712 120006 297956 120034
rect 298356 120006 298692 120034
rect 299000 120006 299428 120034
rect 299552 120006 299888 120034
rect 300196 120006 300532 120034
rect 300840 120006 301176 120034
rect 290936 119734 291010 119762
rect 290740 117360 290792 117366
rect 290740 117302 290792 117308
rect 290936 3534 290964 119734
rect 291384 118108 291436 118114
rect 291384 118050 291436 118056
rect 291108 117428 291160 117434
rect 291108 117370 291160 117376
rect 291016 117360 291068 117366
rect 291016 117302 291068 117308
rect 291028 3670 291056 117302
rect 291016 3664 291068 3670
rect 291016 3606 291068 3612
rect 291120 3602 291148 117370
rect 291108 3596 291160 3602
rect 291108 3538 291160 3544
rect 290924 3528 290976 3534
rect 290924 3470 290976 3476
rect 291396 610 291424 118050
rect 291948 117366 291976 120006
rect 291936 117360 291988 117366
rect 291936 117302 291988 117308
rect 292408 4146 292436 120006
rect 293144 117910 293172 120006
rect 293788 118250 293816 120006
rect 293776 118244 293828 118250
rect 293776 118186 293828 118192
rect 294340 117978 294368 120006
rect 294328 117972 294380 117978
rect 294328 117914 294380 117920
rect 293132 117904 293184 117910
rect 293132 117846 293184 117852
rect 293868 117904 293920 117910
rect 293868 117846 293920 117852
rect 292488 117360 292540 117366
rect 292488 117302 292540 117308
rect 292396 4140 292448 4146
rect 292396 4082 292448 4088
rect 292500 3330 292528 117302
rect 293132 4004 293184 4010
rect 293132 3946 293184 3952
rect 292488 3324 292540 3330
rect 292488 3266 292540 3272
rect 290096 604 290148 610
rect 290096 546 290148 552
rect 290740 604 290792 610
rect 290740 546 290792 552
rect 291384 604 291436 610
rect 291384 546 291436 552
rect 291936 604 291988 610
rect 291936 546 291988 552
rect 290752 480 290780 546
rect 291948 480 291976 546
rect 293144 480 293172 3946
rect 293880 3398 293908 117846
rect 294984 117638 295012 120006
rect 295628 118182 295656 120006
rect 296180 118318 296208 120006
rect 296168 118312 296220 118318
rect 296168 118254 296220 118260
rect 295616 118176 295668 118182
rect 295616 118118 295668 118124
rect 296640 118114 296668 120006
rect 296628 118108 296680 118114
rect 296628 118050 296680 118056
rect 297468 117978 297496 120006
rect 295248 117972 295300 117978
rect 295248 117914 295300 117920
rect 297456 117972 297508 117978
rect 297456 117914 297508 117920
rect 294972 117632 295024 117638
rect 294972 117574 295024 117580
rect 294604 117496 294656 117502
rect 294604 117438 294656 117444
rect 294328 3460 294380 3466
rect 294328 3402 294380 3408
rect 293868 3392 293920 3398
rect 293868 3334 293920 3340
rect 294340 480 294368 3402
rect 294616 3262 294644 117438
rect 295260 3466 295288 117914
rect 297364 117836 297416 117842
rect 297364 117778 297416 117784
rect 295524 3868 295576 3874
rect 295524 3810 295576 3816
rect 295248 3460 295300 3466
rect 295248 3402 295300 3408
rect 294604 3256 294656 3262
rect 294604 3198 294656 3204
rect 295536 480 295564 3810
rect 296720 3800 296772 3806
rect 296720 3742 296772 3748
rect 296732 480 296760 3742
rect 297376 3194 297404 117778
rect 297928 4078 297956 120006
rect 298664 118046 298692 120006
rect 298652 118040 298704 118046
rect 298652 117982 298704 117988
rect 298008 117972 298060 117978
rect 298008 117914 298060 117920
rect 298020 4078 298048 117914
rect 297916 4072 297968 4078
rect 297916 4014 297968 4020
rect 298008 4072 298060 4078
rect 298008 4014 298060 4020
rect 297916 3936 297968 3942
rect 297916 3878 297968 3884
rect 297364 3188 297416 3194
rect 297364 3130 297416 3136
rect 297928 480 297956 3878
rect 299400 3874 299428 120006
rect 299860 117570 299888 120006
rect 300504 117978 300532 120006
rect 300492 117972 300544 117978
rect 300492 117914 300544 117920
rect 299848 117564 299900 117570
rect 299848 117506 299900 117512
rect 301148 117366 301176 120006
rect 301378 119762 301406 120020
rect 302036 120006 302188 120034
rect 302680 120006 303016 120034
rect 303232 120006 303476 120034
rect 303876 120006 304212 120034
rect 304520 120006 304856 120034
rect 305072 120006 305408 120034
rect 305716 120006 306052 120034
rect 306360 120006 306696 120034
rect 306912 120006 307248 120034
rect 307556 120006 307708 120034
rect 308200 120006 308536 120034
rect 308752 120006 309088 120034
rect 309396 120006 309732 120034
rect 310040 120006 310468 120034
rect 310592 120006 310928 120034
rect 311236 120006 311572 120034
rect 301378 119734 301452 119762
rect 301136 117360 301188 117366
rect 301136 117302 301188 117308
rect 301424 116006 301452 119734
rect 302160 117774 302188 120006
rect 302884 118244 302936 118250
rect 302884 118186 302936 118192
rect 302148 117768 302200 117774
rect 302148 117710 302200 117716
rect 302148 117360 302200 117366
rect 302148 117302 302200 117308
rect 301412 116000 301464 116006
rect 301412 115942 301464 115948
rect 301596 116000 301648 116006
rect 301596 115942 301648 115948
rect 301608 109018 301636 115942
rect 301608 108990 301728 109018
rect 301700 108882 301728 108990
rect 301700 108854 302004 108882
rect 301976 106282 302004 108854
rect 301964 106276 302016 106282
rect 301964 106218 302016 106224
rect 301964 99340 302016 99346
rect 301964 99282 302016 99288
rect 301976 96642 302004 99282
rect 301976 96614 302096 96642
rect 302068 89706 302096 96614
rect 301884 89678 302096 89706
rect 301884 77382 301912 89678
rect 301872 77376 301924 77382
rect 301872 77318 301924 77324
rect 302056 77376 302108 77382
rect 302056 77318 302108 77324
rect 302068 77178 302096 77318
rect 302056 77172 302108 77178
rect 302056 77114 302108 77120
rect 301964 67652 302016 67658
rect 301964 67594 302016 67600
rect 301976 60738 302004 67594
rect 301792 60710 302004 60738
rect 301792 57934 301820 60710
rect 301780 57928 301832 57934
rect 301780 57870 301832 57876
rect 301872 48340 301924 48346
rect 301872 48282 301924 48288
rect 301884 41426 301912 48282
rect 301884 41398 302004 41426
rect 301976 31890 302004 41398
rect 301964 31884 302016 31890
rect 301964 31826 302016 31832
rect 302056 31748 302108 31754
rect 302056 31690 302108 31696
rect 302068 26353 302096 31690
rect 301870 26344 301926 26353
rect 301870 26279 301926 26288
rect 302054 26344 302110 26353
rect 302054 26279 302110 26288
rect 301884 26246 301912 26279
rect 301872 26240 301924 26246
rect 301872 26182 301924 26188
rect 302056 8356 302108 8362
rect 302056 8298 302108 8304
rect 299388 3868 299440 3874
rect 299388 3810 299440 3816
rect 302068 3806 302096 8298
rect 302160 3942 302188 117302
rect 302148 3936 302200 3942
rect 302148 3878 302200 3884
rect 302056 3800 302108 3806
rect 302056 3742 302108 3748
rect 299112 3732 299164 3738
rect 299112 3674 299164 3680
rect 299124 480 299152 3674
rect 302608 3596 302660 3602
rect 302608 3538 302660 3544
rect 301412 3256 301464 3262
rect 301412 3198 301464 3204
rect 300308 3188 300360 3194
rect 300308 3130 300360 3136
rect 300320 480 300348 3130
rect 301424 480 301452 3198
rect 302620 480 302648 3538
rect 302896 3194 302924 118186
rect 302988 117366 303016 120006
rect 302976 117360 303028 117366
rect 302976 117302 303028 117308
rect 303448 3602 303476 120006
rect 304184 117706 304212 120006
rect 304828 117910 304856 120006
rect 304816 117904 304868 117910
rect 304816 117846 304868 117852
rect 304172 117700 304224 117706
rect 304172 117642 304224 117648
rect 305380 117366 305408 120006
rect 306024 118658 306052 120006
rect 306012 118652 306064 118658
rect 306012 118594 306064 118600
rect 305644 118312 305696 118318
rect 305644 118254 305696 118260
rect 303528 117360 303580 117366
rect 303528 117302 303580 117308
rect 305368 117360 305420 117366
rect 305368 117302 305420 117308
rect 303540 3738 303568 117302
rect 303528 3732 303580 3738
rect 303528 3674 303580 3680
rect 303804 3664 303856 3670
rect 303804 3606 303856 3612
rect 303436 3596 303488 3602
rect 303436 3538 303488 3544
rect 302884 3188 302936 3194
rect 302884 3130 302936 3136
rect 303816 480 303844 3606
rect 305656 3534 305684 118254
rect 306668 117502 306696 120006
rect 307220 118318 307248 120006
rect 307208 118312 307260 118318
rect 307208 118254 307260 118260
rect 307680 118250 307708 120006
rect 308508 118454 308536 120006
rect 308496 118448 308548 118454
rect 308496 118390 308548 118396
rect 307668 118244 307720 118250
rect 307668 118186 307720 118192
rect 308404 118176 308456 118182
rect 308404 118118 308456 118124
rect 306656 117496 306708 117502
rect 306656 117438 306708 117444
rect 306288 117360 306340 117366
rect 306288 117302 306340 117308
rect 306300 3670 306328 117302
rect 307392 4140 307444 4146
rect 307392 4082 307444 4088
rect 306288 3664 306340 3670
rect 306288 3606 306340 3612
rect 305000 3528 305052 3534
rect 305000 3470 305052 3476
rect 305644 3528 305696 3534
rect 305644 3470 305696 3476
rect 306288 3528 306340 3534
rect 306288 3470 306340 3476
rect 305012 480 305040 3470
rect 306300 3330 306328 3470
rect 306196 3324 306248 3330
rect 306196 3266 306248 3272
rect 306288 3324 306340 3330
rect 306288 3266 306340 3272
rect 306208 480 306236 3266
rect 307404 480 307432 4082
rect 308416 2990 308444 118118
rect 309060 3534 309088 120006
rect 309704 118590 309732 120006
rect 309692 118584 309744 118590
rect 309692 118526 309744 118532
rect 310440 4962 310468 120006
rect 310900 118522 310928 120006
rect 310888 118516 310940 118522
rect 310888 118458 310940 118464
rect 311544 118386 311572 120006
rect 311774 119762 311802 120020
rect 312432 120006 312768 120034
rect 311774 119734 311848 119762
rect 311532 118380 311584 118386
rect 311532 118322 311584 118328
rect 311820 117910 311848 119734
rect 311808 117904 311860 117910
rect 311808 117846 311860 117852
rect 311900 117632 311952 117638
rect 311900 117574 311952 117580
rect 310428 4956 310480 4962
rect 310428 4898 310480 4904
rect 309048 3528 309100 3534
rect 309048 3470 309100 3476
rect 310980 3460 311032 3466
rect 310980 3402 311032 3408
rect 308588 3392 308640 3398
rect 308588 3334 308640 3340
rect 308404 2984 308456 2990
rect 308404 2926 308456 2932
rect 308600 480 308628 3334
rect 309784 3188 309836 3194
rect 309784 3130 309836 3136
rect 309796 480 309824 3130
rect 310992 480 311020 3402
rect 311912 626 311940 117574
rect 312740 117366 312768 120006
rect 313062 119762 313090 120020
rect 313628 120006 313964 120034
rect 314272 120006 314608 120034
rect 314916 120006 315252 120034
rect 315468 120006 315988 120034
rect 316112 120006 316448 120034
rect 316756 120006 317092 120034
rect 313062 119734 313136 119762
rect 312728 117360 312780 117366
rect 312728 117302 312780 117308
rect 313108 4826 313136 119734
rect 313936 117366 313964 120006
rect 314580 117638 314608 120006
rect 314844 118108 314896 118114
rect 314844 118050 314896 118056
rect 314568 117632 314620 117638
rect 314568 117574 314620 117580
rect 313188 117360 313240 117366
rect 313188 117302 313240 117308
rect 313924 117360 313976 117366
rect 313924 117302 313976 117308
rect 314568 117360 314620 117366
rect 314568 117302 314620 117308
rect 313096 4820 313148 4826
rect 313096 4762 313148 4768
rect 313200 3466 313228 117302
rect 314580 4894 314608 117302
rect 314568 4888 314620 4894
rect 314568 4830 314620 4836
rect 313188 3460 313240 3466
rect 313188 3402 313240 3408
rect 314856 3346 314884 118050
rect 315224 117366 315252 120006
rect 315304 117564 315356 117570
rect 315304 117506 315356 117512
rect 315212 117360 315264 117366
rect 315212 117302 315264 117308
rect 315316 4146 315344 117506
rect 315856 117360 315908 117366
rect 315856 117302 315908 117308
rect 315868 5914 315896 117302
rect 315960 5982 315988 120006
rect 316420 117434 316448 120006
rect 316408 117428 316460 117434
rect 316408 117370 316460 117376
rect 317064 117366 317092 120006
rect 317156 120006 317308 120034
rect 317952 120006 318288 120034
rect 318596 120006 318748 120034
rect 319148 120006 319484 120034
rect 319792 120006 320128 120034
rect 320436 120006 320772 120034
rect 320988 120006 321508 120034
rect 321632 120006 321968 120034
rect 322276 120006 322428 120034
rect 317052 117360 317104 117366
rect 317052 117302 317104 117308
rect 317156 6866 317184 120006
rect 318260 117434 318288 120006
rect 317328 117428 317380 117434
rect 317328 117370 317380 117376
rect 318248 117428 318300 117434
rect 318248 117370 318300 117376
rect 317236 117360 317288 117366
rect 317236 117302 317288 117308
rect 317144 6860 317196 6866
rect 317144 6802 317196 6808
rect 317248 6050 317276 117302
rect 317236 6044 317288 6050
rect 317236 5986 317288 5992
rect 315948 5976 316000 5982
rect 315948 5918 316000 5924
rect 315856 5908 315908 5914
rect 315856 5850 315908 5856
rect 315304 4140 315356 4146
rect 315304 4082 315356 4088
rect 315856 4140 315908 4146
rect 315856 4082 315908 4088
rect 314568 3324 314620 3330
rect 314856 3318 315804 3346
rect 314568 3266 314620 3272
rect 313372 2984 313424 2990
rect 313372 2926 313424 2932
rect 311912 598 312216 626
rect 312188 480 312216 598
rect 313384 480 313412 2926
rect 314580 480 314608 3266
rect 315776 480 315804 3318
rect 315868 3262 315896 4082
rect 316960 4072 317012 4078
rect 316960 4014 317012 4020
rect 315856 3256 315908 3262
rect 315856 3198 315908 3204
rect 316972 480 317000 4014
rect 317340 3330 317368 117370
rect 318720 6118 318748 120006
rect 318984 118040 319036 118046
rect 318984 117982 319036 117988
rect 318708 6112 318760 6118
rect 318708 6054 318760 6060
rect 318064 4004 318116 4010
rect 318064 3946 318116 3952
rect 317328 3324 317380 3330
rect 317328 3266 317380 3272
rect 318076 480 318104 3946
rect 318996 610 319024 117982
rect 319456 117366 319484 120006
rect 320100 117502 320128 120006
rect 320088 117496 320140 117502
rect 320088 117438 320140 117444
rect 320744 117366 320772 120006
rect 320824 117564 320876 117570
rect 320824 117506 320876 117512
rect 319444 117360 319496 117366
rect 319444 117302 319496 117308
rect 320088 117360 320140 117366
rect 320088 117302 320140 117308
rect 320732 117360 320784 117366
rect 320732 117302 320784 117308
rect 320100 3398 320128 117302
rect 320456 3868 320508 3874
rect 320456 3810 320508 3816
rect 320088 3392 320140 3398
rect 320088 3334 320140 3340
rect 318984 604 319036 610
rect 318984 546 319036 552
rect 319260 604 319312 610
rect 319260 546 319312 552
rect 319272 480 319300 546
rect 320468 480 320496 3810
rect 320836 3194 320864 117506
rect 321376 117360 321428 117366
rect 321376 117302 321428 117308
rect 321388 4214 321416 117302
rect 321376 4208 321428 4214
rect 321376 4150 321428 4156
rect 321480 4146 321508 120006
rect 321940 118046 321968 120006
rect 321928 118040 321980 118046
rect 321928 117982 321980 117988
rect 321744 117972 321796 117978
rect 321744 117914 321796 117920
rect 321756 12442 321784 117914
rect 322204 117428 322256 117434
rect 322204 117370 322256 117376
rect 321744 12436 321796 12442
rect 321744 12378 321796 12384
rect 321468 4140 321520 4146
rect 321468 4082 321520 4088
rect 322216 3262 322244 117370
rect 322400 116006 322428 120006
rect 322814 119762 322842 120020
rect 323472 120006 323808 120034
rect 322814 119734 322888 119762
rect 322388 116000 322440 116006
rect 322388 115942 322440 115948
rect 322572 116000 322624 116006
rect 322572 115942 322624 115948
rect 322584 109018 322612 115942
rect 322584 108990 322704 109018
rect 322676 106282 322704 108990
rect 322664 106276 322716 106282
rect 322664 106218 322716 106224
rect 322664 99340 322716 99346
rect 322664 99282 322716 99288
rect 322676 96642 322704 99282
rect 322676 96614 322796 96642
rect 322768 89758 322796 96614
rect 322572 89752 322624 89758
rect 322756 89752 322808 89758
rect 322624 89700 322704 89706
rect 322572 89694 322704 89700
rect 322756 89694 322808 89700
rect 322584 89678 322704 89694
rect 322676 86970 322704 89678
rect 322664 86964 322716 86970
rect 322664 86906 322716 86912
rect 322756 77308 322808 77314
rect 322756 77250 322808 77256
rect 322768 66298 322796 77250
rect 322664 66292 322716 66298
rect 322664 66234 322716 66240
rect 322756 66292 322808 66298
rect 322756 66234 322808 66240
rect 322676 60738 322704 66234
rect 322676 60710 322796 60738
rect 322768 57934 322796 60710
rect 322756 57928 322808 57934
rect 322756 57870 322808 57876
rect 322664 48340 322716 48346
rect 322664 48282 322716 48288
rect 322676 41426 322704 48282
rect 322676 41398 322796 41426
rect 322768 38622 322796 41398
rect 322756 38616 322808 38622
rect 322756 38558 322808 38564
rect 322664 29028 322716 29034
rect 322664 28970 322716 28976
rect 322676 22114 322704 28970
rect 322676 22086 322796 22114
rect 322768 12458 322796 22086
rect 322584 12430 322796 12458
rect 322584 4282 322612 12430
rect 322756 12368 322808 12374
rect 322756 12310 322808 12316
rect 322572 4276 322624 4282
rect 322572 4218 322624 4224
rect 322768 3890 322796 12310
rect 322860 4078 322888 119734
rect 323780 117366 323808 120006
rect 324102 119762 324130 120020
rect 324668 120006 325004 120034
rect 325312 120006 325464 120034
rect 325956 120006 326292 120034
rect 326508 120006 326936 120034
rect 327152 120006 327488 120034
rect 327796 120006 328132 120034
rect 324102 119734 324176 119762
rect 323768 117360 323820 117366
rect 323768 117302 323820 117308
rect 324148 4350 324176 119734
rect 324976 117502 325004 120006
rect 325436 117638 325464 120006
rect 325424 117632 325476 117638
rect 325424 117574 325476 117580
rect 324964 117496 325016 117502
rect 324964 117438 325016 117444
rect 326264 117366 326292 120006
rect 326344 117496 326396 117502
rect 326344 117438 326396 117444
rect 324228 117360 324280 117366
rect 324228 117302 324280 117308
rect 326252 117360 326304 117366
rect 326252 117302 326304 117308
rect 324136 4344 324188 4350
rect 324136 4286 324188 4292
rect 322848 4072 322900 4078
rect 322848 4014 322900 4020
rect 324240 4010 324268 117302
rect 325700 114572 325752 114578
rect 325700 114514 325752 114520
rect 325712 104854 325740 114514
rect 325700 104848 325752 104854
rect 325700 104790 325752 104796
rect 325700 95260 325752 95266
rect 325700 95202 325752 95208
rect 325712 85542 325740 95202
rect 325700 85536 325752 85542
rect 325700 85478 325752 85484
rect 325700 75948 325752 75954
rect 325700 75890 325752 75896
rect 325712 66230 325740 75890
rect 325700 66224 325752 66230
rect 325700 66166 325752 66172
rect 325516 56636 325568 56642
rect 325516 56578 325568 56584
rect 325528 48385 325556 56578
rect 325514 48376 325570 48385
rect 325514 48311 325570 48320
rect 325698 48376 325754 48385
rect 325698 48311 325754 48320
rect 325712 46918 325740 48311
rect 325700 46912 325752 46918
rect 325700 46854 325752 46860
rect 325700 29096 325752 29102
rect 325700 29038 325752 29044
rect 325712 27606 325740 29038
rect 325700 27600 325752 27606
rect 325700 27542 325752 27548
rect 326252 9716 326304 9722
rect 326252 9658 326304 9664
rect 326264 9602 326292 9658
rect 326172 9574 326292 9602
rect 324228 4004 324280 4010
rect 324228 3946 324280 3952
rect 324044 3936 324096 3942
rect 322768 3862 322888 3890
rect 324044 3878 324096 3884
rect 321652 3256 321704 3262
rect 321652 3198 321704 3204
rect 322204 3256 322256 3262
rect 322204 3198 322256 3204
rect 320824 3188 320876 3194
rect 320824 3130 320876 3136
rect 321664 480 321692 3198
rect 322860 480 322888 3862
rect 324056 480 324084 3878
rect 326172 3806 326200 9574
rect 326356 3942 326384 117438
rect 326908 6798 326936 120006
rect 327460 117366 327488 120006
rect 328104 117502 328132 120006
rect 328196 120006 328348 120034
rect 328992 120006 329328 120034
rect 329544 120006 329788 120034
rect 330188 120006 330524 120034
rect 330832 120006 331168 120034
rect 331384 120006 331720 120034
rect 332028 120006 332456 120034
rect 332672 120006 333008 120034
rect 333224 120006 333560 120034
rect 328092 117496 328144 117502
rect 328092 117438 328144 117444
rect 326988 117360 327040 117366
rect 326988 117302 327040 117308
rect 327448 117360 327500 117366
rect 327448 117302 327500 117308
rect 326896 6792 326948 6798
rect 326896 6734 326948 6740
rect 327000 4418 327028 117302
rect 328196 6730 328224 120006
rect 329300 117774 329328 120006
rect 329288 117768 329340 117774
rect 329288 117710 329340 117716
rect 328276 117496 328328 117502
rect 328276 117438 328328 117444
rect 328184 6724 328236 6730
rect 328184 6666 328236 6672
rect 328288 4486 328316 117438
rect 328368 117360 328420 117366
rect 328368 117302 328420 117308
rect 328276 4480 328328 4486
rect 328276 4422 328328 4428
rect 326988 4412 327040 4418
rect 326988 4354 327040 4360
rect 326344 3936 326396 3942
rect 326344 3878 326396 3884
rect 328380 3874 328408 117302
rect 329760 4622 329788 120006
rect 329840 117700 329892 117706
rect 329840 117642 329892 117648
rect 329748 4616 329800 4622
rect 329748 4558 329800 4564
rect 328368 3868 328420 3874
rect 328368 3810 328420 3816
rect 325240 3800 325292 3806
rect 325240 3742 325292 3748
rect 326160 3800 326212 3806
rect 326160 3742 326212 3748
rect 325252 480 325280 3742
rect 327632 3732 327684 3738
rect 327632 3674 327684 3680
rect 326436 604 326488 610
rect 326436 546 326488 552
rect 326448 480 326476 546
rect 327644 480 327672 3674
rect 328828 3596 328880 3602
rect 328828 3538 328880 3544
rect 328840 480 328868 3538
rect 329852 626 329880 117642
rect 330496 117638 330524 120006
rect 330484 117632 330536 117638
rect 330484 117574 330536 117580
rect 331036 117632 331088 117638
rect 331036 117574 331088 117580
rect 331048 6662 331076 117574
rect 331036 6656 331088 6662
rect 331036 6598 331088 6604
rect 331140 3602 331168 120006
rect 331312 117836 331364 117842
rect 331312 117778 331364 117784
rect 331128 3596 331180 3602
rect 331128 3538 331180 3544
rect 331324 626 331352 117778
rect 331692 117366 331720 120006
rect 331680 117360 331732 117366
rect 331680 117302 331732 117308
rect 332428 6594 332456 120006
rect 332876 118652 332928 118658
rect 332876 118594 332928 118600
rect 332508 117360 332560 117366
rect 332508 117302 332560 117308
rect 332416 6588 332468 6594
rect 332416 6530 332468 6536
rect 332520 4554 332548 117302
rect 332508 4548 332560 4554
rect 332508 4490 332560 4496
rect 332416 3664 332468 3670
rect 332416 3606 332468 3612
rect 329852 598 330064 626
rect 330036 480 330064 598
rect 331232 598 331352 626
rect 331232 480 331260 598
rect 332428 480 332456 3606
rect 332888 610 332916 118594
rect 332980 117842 333008 120006
rect 332968 117836 333020 117842
rect 332968 117778 333020 117784
rect 333532 117366 333560 120006
rect 333716 120006 333868 120034
rect 334512 120006 334848 120034
rect 335064 120006 335216 120034
rect 335708 120006 336044 120034
rect 336352 120006 336688 120034
rect 336904 120006 337240 120034
rect 337548 120006 337976 120034
rect 338192 120006 338528 120034
rect 338744 120006 339080 120034
rect 333520 117360 333572 117366
rect 333520 117302 333572 117308
rect 333716 6458 333744 120006
rect 334820 118454 334848 120006
rect 334808 118448 334860 118454
rect 334808 118390 334860 118396
rect 334624 118312 334676 118318
rect 334624 118254 334676 118260
rect 333980 117904 334032 117910
rect 333980 117846 334032 117852
rect 333888 117836 333940 117842
rect 333888 117778 333940 117784
rect 333796 117360 333848 117366
rect 333796 117302 333848 117308
rect 333704 6452 333756 6458
rect 333704 6394 333756 6400
rect 333808 4690 333836 117302
rect 333796 4684 333848 4690
rect 333796 4626 333848 4632
rect 333900 3738 333928 117778
rect 333888 3732 333940 3738
rect 333888 3674 333940 3680
rect 333992 3346 334020 117846
rect 334636 3806 334664 118254
rect 335188 5506 335216 120006
rect 335268 118448 335320 118454
rect 335268 118390 335320 118396
rect 335176 5500 335228 5506
rect 335176 5442 335228 5448
rect 334624 3800 334676 3806
rect 334624 3742 334676 3748
rect 335280 3670 335308 118390
rect 336016 117366 336044 120006
rect 336660 118318 336688 120006
rect 336648 118312 336700 118318
rect 336648 118254 336700 118260
rect 336924 118244 336976 118250
rect 336924 118186 336976 118192
rect 336004 117360 336056 117366
rect 336004 117302 336056 117308
rect 336648 117360 336700 117366
rect 336648 117302 336700 117308
rect 336660 6526 336688 117302
rect 336648 6520 336700 6526
rect 336648 6462 336700 6468
rect 335912 3800 335964 3806
rect 335912 3742 335964 3748
rect 335268 3664 335320 3670
rect 335268 3606 335320 3612
rect 333992 3318 334756 3346
rect 332876 604 332928 610
rect 332876 546 332928 552
rect 333612 604 333664 610
rect 333612 546 333664 552
rect 333624 480 333652 546
rect 334728 480 334756 3318
rect 335924 480 335952 3742
rect 336936 610 336964 118186
rect 337212 117366 337240 120006
rect 337200 117360 337252 117366
rect 337200 117302 337252 117308
rect 337948 6390 337976 120006
rect 338396 118584 338448 118590
rect 338396 118526 338448 118532
rect 338028 117360 338080 117366
rect 338028 117302 338080 117308
rect 337936 6384 337988 6390
rect 337936 6326 337988 6332
rect 338040 4758 338068 117302
rect 338028 4752 338080 4758
rect 338028 4694 338080 4700
rect 338408 626 338436 118526
rect 338500 118250 338528 120006
rect 338488 118244 338540 118250
rect 338488 118186 338540 118192
rect 339052 117366 339080 120006
rect 339374 119762 339402 120020
rect 340032 120006 340368 120034
rect 340584 120006 340736 120034
rect 341228 120006 341564 120034
rect 341872 120006 342208 120034
rect 342424 120006 342760 120034
rect 343068 120006 343496 120034
rect 343712 120006 344048 120034
rect 344264 120006 344600 120034
rect 339328 119734 339402 119762
rect 339040 117360 339092 117366
rect 339040 117302 339092 117308
rect 339328 6254 339356 119734
rect 339592 118652 339644 118658
rect 339592 118594 339644 118600
rect 339408 117360 339460 117366
rect 339408 117302 339460 117308
rect 339316 6248 339368 6254
rect 339316 6190 339368 6196
rect 339420 5438 339448 117302
rect 339408 5432 339460 5438
rect 339408 5374 339460 5380
rect 339500 3528 339552 3534
rect 339500 3470 339552 3476
rect 336924 604 336976 610
rect 336924 546 336976 552
rect 337108 604 337160 610
rect 337108 546 337160 552
rect 338316 598 338436 626
rect 337120 480 337148 546
rect 338316 480 338344 598
rect 339512 480 339540 3470
rect 339604 3346 339632 118594
rect 340340 117366 340368 120006
rect 340328 117360 340380 117366
rect 340328 117302 340380 117308
rect 340708 5370 340736 120006
rect 341340 118516 341392 118522
rect 341340 118458 341392 118464
rect 340788 117360 340840 117366
rect 340788 117302 340840 117308
rect 340696 5364 340748 5370
rect 340696 5306 340748 5312
rect 339604 3318 340736 3346
rect 340708 480 340736 3318
rect 340800 2854 340828 117302
rect 341352 115938 341380 118458
rect 341536 117366 341564 120006
rect 342180 118454 342208 120006
rect 342168 118448 342220 118454
rect 342168 118390 342220 118396
rect 342732 117366 342760 120006
rect 341524 117360 341576 117366
rect 341524 117302 341576 117308
rect 342168 117360 342220 117366
rect 342168 117302 342220 117308
rect 342720 117360 342772 117366
rect 342720 117302 342772 117308
rect 341064 115932 341116 115938
rect 341064 115874 341116 115880
rect 341340 115932 341392 115938
rect 341340 115874 341392 115880
rect 341076 106321 341104 115874
rect 341062 106312 341118 106321
rect 341062 106247 341118 106256
rect 341246 106312 341302 106321
rect 341246 106247 341302 106256
rect 341260 99414 341288 106247
rect 341248 99408 341300 99414
rect 341248 99350 341300 99356
rect 341340 99340 341392 99346
rect 341340 99282 341392 99288
rect 341352 96626 341380 99282
rect 341064 96620 341116 96626
rect 341064 96562 341116 96568
rect 341340 96620 341392 96626
rect 341340 96562 341392 96568
rect 341076 87009 341104 96562
rect 341062 87000 341118 87009
rect 341062 86935 341118 86944
rect 341246 87000 341302 87009
rect 341246 86935 341302 86944
rect 341260 79914 341288 86935
rect 341260 79886 341380 79914
rect 341352 77178 341380 79886
rect 341340 77172 341392 77178
rect 341340 77114 341392 77120
rect 341432 67652 341484 67658
rect 341432 67594 341484 67600
rect 341444 60738 341472 67594
rect 341444 60710 341564 60738
rect 341536 51202 341564 60710
rect 341524 51196 341576 51202
rect 341524 51138 341576 51144
rect 341524 45620 341576 45626
rect 341524 45562 341576 45568
rect 341536 45490 341564 45562
rect 341524 45484 341576 45490
rect 341524 45426 341576 45432
rect 341432 38276 341484 38282
rect 341432 38218 341484 38224
rect 341444 31686 341472 38218
rect 341432 31680 341484 31686
rect 341432 31622 341484 31628
rect 341524 31680 341576 31686
rect 341524 31622 341576 31628
rect 341536 12458 341564 31622
rect 341536 12430 341656 12458
rect 341628 3602 341656 12430
rect 342180 6322 342208 117302
rect 342168 6316 342220 6322
rect 342168 6258 342220 6264
rect 343468 6186 343496 120006
rect 343916 118380 343968 118386
rect 343916 118322 343968 118328
rect 343548 117360 343600 117366
rect 343548 117302 343600 117308
rect 343456 6180 343508 6186
rect 343456 6122 343508 6128
rect 343560 5302 343588 117302
rect 343548 5296 343600 5302
rect 343548 5238 343600 5244
rect 341892 4956 341944 4962
rect 341892 4898 341944 4904
rect 341616 3596 341668 3602
rect 341616 3538 341668 3544
rect 340788 2848 340840 2854
rect 340788 2790 340840 2796
rect 341904 480 341932 4898
rect 343088 3596 343140 3602
rect 343088 3538 343140 3544
rect 343100 480 343128 3538
rect 343928 610 343956 118322
rect 344020 117434 344048 120006
rect 344008 117428 344060 117434
rect 344008 117370 344060 117376
rect 344572 117366 344600 120006
rect 344756 120006 344908 120034
rect 345552 120006 345888 120034
rect 346104 120006 346348 120034
rect 346748 120006 347084 120034
rect 347300 120006 347636 120034
rect 347944 120006 348280 120034
rect 348588 120006 349016 120034
rect 349140 120006 349476 120034
rect 349784 120006 350120 120034
rect 344560 117360 344612 117366
rect 344560 117302 344612 117308
rect 344756 7750 344784 120006
rect 345860 118658 345888 120006
rect 345848 118652 345900 118658
rect 345848 118594 345900 118600
rect 345112 118176 345164 118182
rect 345112 118118 345164 118124
rect 344928 117428 344980 117434
rect 344928 117370 344980 117376
rect 344836 117360 344888 117366
rect 344836 117302 344888 117308
rect 344744 7744 344796 7750
rect 344744 7686 344796 7692
rect 344848 5234 344876 117302
rect 344836 5228 344888 5234
rect 344836 5170 344888 5176
rect 344940 3534 344968 117370
rect 344928 3528 344980 3534
rect 344928 3470 344980 3476
rect 345124 626 345152 118118
rect 346320 5166 346348 120006
rect 347056 117366 347084 120006
rect 347608 118522 347636 120006
rect 347596 118516 347648 118522
rect 347596 118458 347648 118464
rect 348252 117366 348280 120006
rect 347044 117360 347096 117366
rect 347044 117302 347096 117308
rect 347688 117360 347740 117366
rect 347688 117302 347740 117308
rect 348240 117360 348292 117366
rect 348240 117302 348292 117308
rect 347700 7682 347728 117302
rect 347688 7676 347740 7682
rect 347688 7618 347740 7624
rect 348988 7614 349016 120006
rect 349448 118182 349476 120006
rect 349436 118176 349488 118182
rect 349436 118118 349488 118124
rect 350092 117366 350120 120006
rect 350414 119762 350442 120020
rect 350980 120006 351316 120034
rect 351624 120006 351776 120034
rect 352268 120006 352604 120034
rect 352820 120006 353156 120034
rect 353464 120006 353800 120034
rect 354108 120006 354536 120034
rect 354660 120006 354996 120034
rect 355304 120006 355640 120034
rect 350368 119734 350442 119762
rect 349068 117360 349120 117366
rect 349068 117302 349120 117308
rect 350080 117360 350132 117366
rect 350080 117302 350132 117308
rect 348976 7608 349028 7614
rect 348976 7550 349028 7556
rect 346308 5160 346360 5166
rect 346308 5102 346360 5108
rect 349080 5098 349108 117302
rect 350368 9178 350396 119734
rect 351288 117366 351316 120006
rect 350448 117360 350500 117366
rect 350448 117302 350500 117308
rect 351276 117360 351328 117366
rect 351276 117302 351328 117308
rect 350356 9172 350408 9178
rect 350356 9114 350408 9120
rect 349068 5092 349120 5098
rect 349068 5034 349120 5040
rect 350460 5030 350488 117302
rect 351368 5908 351420 5914
rect 351368 5850 351420 5856
rect 350448 5024 350500 5030
rect 350448 4966 350500 4972
rect 349068 4888 349120 4894
rect 349068 4830 349120 4836
rect 347872 4820 347924 4826
rect 347872 4762 347924 4768
rect 346676 3460 346728 3466
rect 346676 3402 346728 3408
rect 343916 604 343968 610
rect 343916 546 343968 552
rect 344284 604 344336 610
rect 345124 598 345520 626
rect 344284 546 344336 552
rect 344296 480 344324 546
rect 345492 480 345520 598
rect 346688 480 346716 3402
rect 347884 480 347912 4762
rect 349080 480 349108 4830
rect 350264 3188 350316 3194
rect 350264 3130 350316 3136
rect 350276 480 350304 3130
rect 351380 480 351408 5850
rect 351748 4894 351776 120006
rect 352576 117366 352604 120006
rect 353128 117910 353156 120006
rect 353116 117904 353168 117910
rect 353116 117846 353168 117852
rect 353772 117366 353800 120006
rect 354312 118108 354364 118114
rect 354312 118050 354364 118056
rect 354324 117978 354352 118050
rect 354312 117972 354364 117978
rect 354312 117914 354364 117920
rect 351828 117360 351880 117366
rect 351828 117302 351880 117308
rect 352564 117360 352616 117366
rect 352564 117302 352616 117308
rect 353208 117360 353260 117366
rect 353208 117302 353260 117308
rect 353760 117360 353812 117366
rect 353760 117302 353812 117308
rect 351736 4888 351788 4894
rect 351736 4830 351788 4836
rect 351840 3466 351868 117302
rect 353220 9110 353248 117302
rect 353208 9104 353260 9110
rect 353208 9046 353260 9052
rect 354508 9042 354536 120006
rect 354968 117638 354996 120006
rect 354956 117632 355008 117638
rect 354956 117574 355008 117580
rect 355612 117366 355640 120006
rect 355934 119762 355962 120020
rect 356500 120006 356836 120034
rect 357144 120006 357388 120034
rect 357788 120006 358124 120034
rect 358340 120006 358768 120034
rect 358984 120006 359320 120034
rect 359628 120006 360056 120034
rect 360180 120006 360516 120034
rect 360824 120006 361160 120034
rect 355888 119734 355962 119762
rect 354588 117360 354640 117366
rect 354588 117302 354640 117308
rect 355600 117360 355652 117366
rect 355600 117302 355652 117308
rect 354496 9036 354548 9042
rect 354496 8978 354548 8984
rect 352564 5976 352616 5982
rect 352564 5918 352616 5924
rect 351828 3460 351880 3466
rect 351828 3402 351880 3408
rect 352576 480 352604 5918
rect 354600 4962 354628 117302
rect 355888 8974 355916 119734
rect 356808 117706 356836 120006
rect 356796 117700 356848 117706
rect 356796 117642 356848 117648
rect 355968 117360 356020 117366
rect 355968 117302 356020 117308
rect 355876 8968 355928 8974
rect 355876 8910 355928 8916
rect 354956 6044 355008 6050
rect 354956 5986 355008 5992
rect 354588 4956 354640 4962
rect 354588 4898 354640 4904
rect 353760 3324 353812 3330
rect 353760 3266 353812 3272
rect 353772 480 353800 3266
rect 354968 480 354996 5986
rect 355980 4826 356008 117302
rect 356152 6860 356204 6866
rect 356152 6802 356204 6808
rect 355968 4820 356020 4826
rect 355968 4762 356020 4768
rect 356164 480 356192 6802
rect 357360 4865 357388 120006
rect 357992 117768 358044 117774
rect 357992 117710 358044 117716
rect 358004 103578 358032 117710
rect 358096 117570 358124 120006
rect 358176 117972 358228 117978
rect 358176 117914 358228 117920
rect 358084 117564 358136 117570
rect 358084 117506 358136 117512
rect 358004 103550 358124 103578
rect 358096 99362 358124 103550
rect 358004 99334 358124 99362
rect 358004 80170 358032 99334
rect 357992 80164 358044 80170
rect 357992 80106 358044 80112
rect 357992 79960 358044 79966
rect 357992 79902 358044 79908
rect 358004 70394 358032 79902
rect 357912 70366 358032 70394
rect 357912 70258 357940 70366
rect 357912 70230 358032 70258
rect 358004 51082 358032 70230
rect 357912 51066 358032 51082
rect 357900 51060 358032 51066
rect 357952 51054 358032 51060
rect 358084 51060 358136 51066
rect 357900 51002 357952 51008
rect 358084 51002 358136 51008
rect 357912 50971 357940 51002
rect 358096 48278 358124 51002
rect 358084 48272 358136 48278
rect 358084 48214 358136 48220
rect 357992 38684 358044 38690
rect 357992 38626 358044 38632
rect 358004 29102 358032 38626
rect 357992 29096 358044 29102
rect 357992 29038 358044 29044
rect 357716 26376 357768 26382
rect 357716 26318 357768 26324
rect 357728 26246 357756 26318
rect 357716 26240 357768 26246
rect 357716 26182 357768 26188
rect 357900 22024 357952 22030
rect 357900 21966 357952 21972
rect 357912 8362 357940 21966
rect 357808 8356 357860 8362
rect 357808 8298 357860 8304
rect 357900 8356 357952 8362
rect 357900 8298 357952 8304
rect 357346 4856 357402 4865
rect 357346 4791 357402 4800
rect 357820 3330 357848 8298
rect 358188 3602 358216 117914
rect 358636 117564 358688 117570
rect 358636 117506 358688 117512
rect 358648 8498 358676 117506
rect 358636 8492 358688 8498
rect 358636 8434 358688 8440
rect 358740 7206 358768 120006
rect 359292 117638 359320 120006
rect 359280 117632 359332 117638
rect 359280 117574 359332 117580
rect 360028 8566 360056 120006
rect 360488 117638 360516 120006
rect 360108 117632 360160 117638
rect 360108 117574 360160 117580
rect 360476 117632 360528 117638
rect 360476 117574 360528 117580
rect 360016 8560 360068 8566
rect 360016 8502 360068 8508
rect 358728 7200 358780 7206
rect 358728 7142 358780 7148
rect 360120 7138 360148 117574
rect 361132 117366 361160 120006
rect 361454 119762 361482 120020
rect 362020 120006 362356 120034
rect 362664 120006 362908 120034
rect 363308 120006 363644 120034
rect 363860 120006 364104 120034
rect 364504 120006 364840 120034
rect 365056 120006 365576 120034
rect 365700 120006 366036 120034
rect 366344 120006 366680 120034
rect 361408 119734 361482 119762
rect 361120 117360 361172 117366
rect 361120 117302 361172 117308
rect 361408 8702 361436 119734
rect 362328 118590 362356 120006
rect 362316 118584 362368 118590
rect 362316 118526 362368 118532
rect 361488 117360 361540 117366
rect 361488 117302 361540 117308
rect 361396 8696 361448 8702
rect 361396 8638 361448 8644
rect 361500 7274 361528 117302
rect 362880 7342 362908 120006
rect 363512 118040 363564 118046
rect 363512 117982 363564 117988
rect 363524 117178 363552 117982
rect 363616 117366 363644 120006
rect 364076 117774 364104 120006
rect 364064 117768 364116 117774
rect 364064 117710 364116 117716
rect 364812 117366 364840 120006
rect 363604 117360 363656 117366
rect 363604 117302 363656 117308
rect 364248 117360 364300 117366
rect 364248 117302 364300 117308
rect 364800 117360 364852 117366
rect 364800 117302 364852 117308
rect 363524 117150 363644 117178
rect 362868 7336 362920 7342
rect 362868 7278 362920 7284
rect 361488 7268 361540 7274
rect 361488 7210 361540 7216
rect 360108 7132 360160 7138
rect 360108 7074 360160 7080
rect 358544 6112 358596 6118
rect 358544 6054 358596 6060
rect 358176 3596 358228 3602
rect 358176 3538 358228 3544
rect 357808 3324 357860 3330
rect 357808 3266 357860 3272
rect 357348 3256 357400 3262
rect 357348 3198 357400 3204
rect 357360 480 357388 3198
rect 358556 480 358584 6054
rect 362132 4208 362184 4214
rect 362132 4150 362184 4156
rect 360936 3596 360988 3602
rect 360936 3538 360988 3544
rect 359740 3392 359792 3398
rect 359740 3334 359792 3340
rect 359752 480 359780 3334
rect 360948 480 360976 3538
rect 362144 480 362172 4150
rect 363616 4146 363644 117150
rect 364260 8634 364288 117302
rect 365548 8770 365576 120006
rect 366008 118386 366036 120006
rect 365996 118380 366048 118386
rect 365996 118322 366048 118328
rect 366652 117366 366680 120006
rect 366882 119762 366910 120020
rect 367540 120006 367876 120034
rect 368184 120006 368428 120034
rect 368736 120006 369072 120034
rect 369380 120006 369716 120034
rect 370024 120006 370360 120034
rect 370576 120006 371096 120034
rect 371220 120006 371556 120034
rect 371864 120006 372200 120034
rect 366882 119734 366956 119762
rect 365628 117360 365680 117366
rect 365628 117302 365680 117308
rect 366640 117360 366692 117366
rect 366640 117302 366692 117308
rect 365536 8764 365588 8770
rect 365536 8706 365588 8712
rect 364248 8628 364300 8634
rect 364248 8570 364300 8576
rect 365640 7410 365668 117302
rect 366928 8838 366956 119734
rect 367848 117502 367876 120006
rect 367836 117496 367888 117502
rect 367836 117438 367888 117444
rect 367008 117360 367060 117366
rect 367008 117302 367060 117308
rect 366916 8832 366968 8838
rect 366916 8774 366968 8780
rect 367020 7478 367048 117302
rect 368400 9654 368428 120006
rect 369044 117366 369072 120006
rect 369688 118182 369716 120006
rect 369676 118176 369728 118182
rect 369676 118118 369728 118124
rect 369216 118108 369268 118114
rect 369216 118050 369268 118056
rect 369124 117564 369176 117570
rect 369124 117506 369176 117512
rect 369032 117360 369084 117366
rect 369032 117302 369084 117308
rect 368388 9648 368440 9654
rect 368388 9590 368440 9596
rect 367008 7472 367060 7478
rect 367008 7414 367060 7420
rect 365628 7404 365680 7410
rect 365628 7346 365680 7352
rect 369136 6882 369164 117506
rect 368952 6854 369164 6882
rect 365720 4276 365772 4282
rect 365720 4218 365772 4224
rect 363328 4140 363380 4146
rect 363328 4082 363380 4088
rect 363604 4140 363656 4146
rect 363604 4082 363656 4088
rect 364524 4140 364576 4146
rect 364524 4082 364576 4088
rect 363340 480 363368 4082
rect 364536 480 364564 4082
rect 365732 480 365760 4218
rect 368020 4004 368072 4010
rect 368020 3946 368072 3952
rect 366916 3596 366968 3602
rect 366916 3538 366968 3544
rect 366928 480 366956 3538
rect 368032 480 368060 3946
rect 368952 2922 368980 6854
rect 369124 4344 369176 4350
rect 369124 4286 369176 4292
rect 368940 2916 368992 2922
rect 368940 2858 368992 2864
rect 369136 2258 369164 4286
rect 369228 3602 369256 118050
rect 370332 117366 370360 120006
rect 369768 117360 369820 117366
rect 369768 117302 369820 117308
rect 370320 117360 370372 117366
rect 370320 117302 370372 117308
rect 369780 8906 369808 117302
rect 371068 10742 371096 120006
rect 371528 117434 371556 120006
rect 371516 117428 371568 117434
rect 371516 117370 371568 117376
rect 372172 117366 372200 120006
rect 372402 119762 372430 120020
rect 373060 120006 373396 120034
rect 373704 120006 373948 120034
rect 374256 120006 374592 120034
rect 374900 120006 375328 120034
rect 375544 120006 375880 120034
rect 376096 120006 376616 120034
rect 376740 120006 377076 120034
rect 377384 120006 377720 120034
rect 372356 119734 372430 119762
rect 371148 117360 371200 117366
rect 371148 117302 371200 117308
rect 372160 117360 372212 117366
rect 372160 117302 372212 117308
rect 371056 10736 371108 10742
rect 371056 10678 371108 10684
rect 371160 9586 371188 117302
rect 372356 10674 372384 119734
rect 373368 118114 373396 120006
rect 373356 118108 373408 118114
rect 373356 118050 373408 118056
rect 372528 117428 372580 117434
rect 372528 117370 372580 117376
rect 372436 117360 372488 117366
rect 372436 117302 372488 117308
rect 372344 10668 372396 10674
rect 372344 10610 372396 10616
rect 371148 9580 371200 9586
rect 371148 9522 371200 9528
rect 372448 9518 372476 117302
rect 372436 9512 372488 9518
rect 372436 9454 372488 9460
rect 369768 8900 369820 8906
rect 369768 8842 369820 8848
rect 370412 3936 370464 3942
rect 370412 3878 370464 3884
rect 369216 3596 369268 3602
rect 369216 3538 369268 3544
rect 369136 2230 369256 2258
rect 369228 480 369256 2230
rect 370424 480 370452 3878
rect 371608 3596 371660 3602
rect 371608 3538 371660 3544
rect 371620 480 371648 3538
rect 372540 3126 372568 117370
rect 373920 5642 373948 120006
rect 374564 117366 374592 120006
rect 374644 118312 374696 118318
rect 374644 118254 374696 118260
rect 374552 117360 374604 117366
rect 374552 117302 374604 117308
rect 374000 6792 374052 6798
rect 374000 6734 374052 6740
rect 373908 5636 373960 5642
rect 373908 5578 373960 5584
rect 372804 4412 372856 4418
rect 372804 4354 372856 4360
rect 372528 3120 372580 3126
rect 372528 3062 372580 3068
rect 372816 480 372844 4354
rect 374012 480 374040 6734
rect 374656 3942 374684 118254
rect 375196 117360 375248 117366
rect 375196 117302 375248 117308
rect 375208 10606 375236 117302
rect 375196 10600 375248 10606
rect 375196 10542 375248 10548
rect 374644 3936 374696 3942
rect 374644 3878 374696 3884
rect 375196 3868 375248 3874
rect 375196 3810 375248 3816
rect 375208 480 375236 3810
rect 375300 3194 375328 120006
rect 375852 117366 375880 120006
rect 376024 118516 376076 118522
rect 376024 118458 376076 118464
rect 375840 117360 375892 117366
rect 375840 117302 375892 117308
rect 375288 3188 375340 3194
rect 375288 3130 375340 3136
rect 376036 2990 376064 118458
rect 376588 10538 376616 120006
rect 377048 118318 377076 120006
rect 377036 118312 377088 118318
rect 377036 118254 377088 118260
rect 377404 117496 377456 117502
rect 377404 117438 377456 117444
rect 376668 117360 376720 117366
rect 376668 117302 376720 117308
rect 376576 10532 376628 10538
rect 376576 10474 376628 10480
rect 376680 5574 376708 117302
rect 376668 5568 376720 5574
rect 376668 5510 376720 5516
rect 376392 4480 376444 4486
rect 376392 4422 376444 4428
rect 376024 2984 376076 2990
rect 376024 2926 376076 2932
rect 376404 480 376432 4422
rect 377416 3058 377444 117438
rect 377692 117366 377720 120006
rect 377922 119762 377950 120020
rect 378580 120006 378916 120034
rect 379224 120006 379376 120034
rect 379776 120006 380112 120034
rect 380420 120006 380756 120034
rect 381064 120006 381400 120034
rect 381616 120006 382136 120034
rect 382260 120006 382596 120034
rect 382812 120006 382964 120034
rect 377922 119734 377996 119762
rect 377680 117360 377732 117366
rect 377680 117302 377732 117308
rect 377968 10470 377996 119734
rect 378888 117366 378916 120006
rect 378048 117360 378100 117366
rect 378048 117302 378100 117308
rect 378876 117360 378928 117366
rect 378876 117302 378928 117308
rect 377956 10464 378008 10470
rect 377956 10406 378008 10412
rect 377588 6724 377640 6730
rect 377588 6666 377640 6672
rect 377404 3052 377456 3058
rect 377404 2994 377456 3000
rect 377600 480 377628 6666
rect 378060 5710 378088 117302
rect 379348 5846 379376 120006
rect 380084 117366 380112 120006
rect 380728 117978 380756 120006
rect 380716 117972 380768 117978
rect 380716 117914 380768 117920
rect 381372 117366 381400 120006
rect 379428 117360 379480 117366
rect 379428 117302 379480 117308
rect 380072 117360 380124 117366
rect 380072 117302 380124 117308
rect 380808 117360 380860 117366
rect 380808 117302 380860 117308
rect 381360 117360 381412 117366
rect 381360 117302 381412 117308
rect 379336 5840 379388 5846
rect 379336 5782 379388 5788
rect 378048 5704 378100 5710
rect 378048 5646 378100 5652
rect 378784 3324 378836 3330
rect 378784 3266 378836 3272
rect 378796 480 378824 3266
rect 379440 3262 379468 117302
rect 380820 10402 380848 117302
rect 380808 10396 380860 10402
rect 380808 10338 380860 10344
rect 382108 10334 382136 120006
rect 382568 117366 382596 120006
rect 382188 117360 382240 117366
rect 382188 117302 382240 117308
rect 382556 117360 382608 117366
rect 382556 117302 382608 117308
rect 382096 10328 382148 10334
rect 382096 10270 382148 10276
rect 381176 6656 381228 6662
rect 381176 6598 381228 6604
rect 379980 4616 380032 4622
rect 379980 4558 380032 4564
rect 379428 3256 379480 3262
rect 379428 3198 379480 3204
rect 379992 480 380020 4558
rect 381188 480 381216 6598
rect 382200 5778 382228 117302
rect 382936 116006 382964 120006
rect 383442 119762 383470 120020
rect 384100 120006 384436 120034
rect 384652 120006 384988 120034
rect 385296 120006 385632 120034
rect 385940 120006 386276 120034
rect 386492 120006 386828 120034
rect 387136 120006 387656 120034
rect 387780 120006 388116 120034
rect 383442 119734 383516 119762
rect 382924 116000 382976 116006
rect 382924 115942 382976 115948
rect 383108 116000 383160 116006
rect 383108 115942 383160 115948
rect 383120 109018 383148 115942
rect 383120 108990 383332 109018
rect 383304 99482 383332 108990
rect 383292 99476 383344 99482
rect 383292 99418 383344 99424
rect 383200 99340 383252 99346
rect 383200 99282 383252 99288
rect 383212 96626 383240 99282
rect 383200 96620 383252 96626
rect 383200 96562 383252 96568
rect 383108 87032 383160 87038
rect 383108 86974 383160 86980
rect 383120 79914 383148 86974
rect 383120 79886 383240 79914
rect 383212 77178 383240 79886
rect 383200 77172 383252 77178
rect 383200 77114 383252 77120
rect 383292 67652 383344 67658
rect 383292 67594 383344 67600
rect 383304 60858 383332 67594
rect 383292 60852 383344 60858
rect 383292 60794 383344 60800
rect 383200 60716 383252 60722
rect 383200 60658 383252 60664
rect 383212 57934 383240 60658
rect 383200 57928 383252 57934
rect 383200 57870 383252 57876
rect 383292 48340 383344 48346
rect 383292 48282 383344 48288
rect 383304 43466 383332 48282
rect 383212 43438 383332 43466
rect 383212 38622 383240 43438
rect 383200 38616 383252 38622
rect 383200 38558 383252 38564
rect 383292 29028 383344 29034
rect 383292 28970 383344 28976
rect 383304 28914 383332 28970
rect 383304 28886 383424 28914
rect 383396 25294 383424 28886
rect 383384 25288 383436 25294
rect 383384 25230 383436 25236
rect 383384 19372 383436 19378
rect 383384 19314 383436 19320
rect 383396 19258 383424 19314
rect 383304 19230 383424 19258
rect 383304 12578 383332 19230
rect 383292 12572 383344 12578
rect 383292 12514 383344 12520
rect 383292 9716 383344 9722
rect 383292 9658 383344 9664
rect 383304 7546 383332 9658
rect 383292 7540 383344 7546
rect 383292 7482 383344 7488
rect 383488 5982 383516 119734
rect 384212 118244 384264 118250
rect 384212 118186 384264 118192
rect 384224 118130 384252 118186
rect 384224 118102 384344 118130
rect 383568 117360 383620 117366
rect 383568 117302 383620 117308
rect 383476 5976 383528 5982
rect 383476 5918 383528 5924
rect 383580 5828 383608 117302
rect 383488 5800 383608 5828
rect 382188 5772 382240 5778
rect 382188 5714 382240 5720
rect 382372 3800 382424 3806
rect 382372 3742 382424 3748
rect 382384 480 382412 3742
rect 383488 3330 383516 5800
rect 383568 4548 383620 4554
rect 383568 4490 383620 4496
rect 383476 3324 383528 3330
rect 383476 3266 383528 3272
rect 383580 480 383608 4490
rect 384316 3942 384344 118102
rect 384408 117570 384436 120006
rect 384396 117564 384448 117570
rect 384396 117506 384448 117512
rect 384960 8294 384988 120006
rect 385604 117366 385632 120006
rect 386248 118250 386276 120006
rect 386236 118244 386288 118250
rect 386236 118186 386288 118192
rect 386800 117366 386828 120006
rect 387628 118674 387656 120006
rect 387536 118646 387656 118674
rect 385592 117360 385644 117366
rect 385592 117302 385644 117308
rect 386328 117360 386380 117366
rect 386328 117302 386380 117308
rect 386788 117360 386840 117366
rect 386788 117302 386840 117308
rect 384948 8288 385000 8294
rect 384948 8230 385000 8236
rect 384672 6588 384724 6594
rect 384672 6530 384724 6536
rect 384304 3936 384356 3942
rect 384304 3878 384356 3884
rect 384684 480 384712 6530
rect 386340 5914 386368 117302
rect 387536 109070 387564 118646
rect 388088 117366 388116 120006
rect 387616 117360 387668 117366
rect 387616 117302 387668 117308
rect 388076 117360 388128 117366
rect 388076 117302 388128 117308
rect 387524 109064 387576 109070
rect 387524 109006 387576 109012
rect 387628 8226 387656 117302
rect 388732 115938 388760 120278
rect 414736 120142 414888 120170
rect 388962 119762 388990 120020
rect 389620 120006 389956 120034
rect 390172 120006 390508 120034
rect 390816 120006 391152 120034
rect 391460 120006 391888 120034
rect 392012 120006 392348 120034
rect 392656 120006 393176 120034
rect 393300 120006 393636 120034
rect 393852 120006 394372 120034
rect 394496 120006 394648 120034
rect 395140 120006 395476 120034
rect 395692 120006 395936 120034
rect 396336 120006 396672 120034
rect 396980 120006 397316 120034
rect 397532 120006 397868 120034
rect 398176 120006 398696 120034
rect 398820 120006 399156 120034
rect 399372 120006 399708 120034
rect 388962 119734 389036 119762
rect 388720 115932 388772 115938
rect 388720 115874 388772 115880
rect 388904 115932 388956 115938
rect 388904 115874 388956 115880
rect 387708 109064 387760 109070
rect 387708 109006 387760 109012
rect 387616 8220 387668 8226
rect 387616 8162 387668 8168
rect 387720 6050 387748 109006
rect 388916 106321 388944 115874
rect 388718 106312 388774 106321
rect 388902 106312 388958 106321
rect 388718 106247 388720 106256
rect 388772 106247 388774 106256
rect 388812 106276 388864 106282
rect 388720 106218 388772 106224
rect 388902 106247 388958 106256
rect 388812 106218 388864 106224
rect 388824 96642 388852 106218
rect 388732 96626 388852 96642
rect 388720 96620 388852 96626
rect 388772 96614 388852 96620
rect 388720 96562 388772 96568
rect 388732 96531 388760 96562
rect 388628 87032 388680 87038
rect 388628 86974 388680 86980
rect 388640 82090 388668 86974
rect 388640 82062 388852 82090
rect 388824 79914 388852 82062
rect 388732 79886 388852 79914
rect 388732 77178 388760 79886
rect 388720 77172 388772 77178
rect 388720 77114 388772 77120
rect 388812 67652 388864 67658
rect 388812 67594 388864 67600
rect 388824 60858 388852 67594
rect 388812 60852 388864 60858
rect 388812 60794 388864 60800
rect 388720 60716 388772 60722
rect 388720 60658 388772 60664
rect 388732 57934 388760 60658
rect 388720 57928 388772 57934
rect 388720 57870 388772 57876
rect 388812 48340 388864 48346
rect 388812 48282 388864 48288
rect 388824 43466 388852 48282
rect 388732 43438 388852 43466
rect 388732 31754 388760 43438
rect 388720 31748 388772 31754
rect 388720 31690 388772 31696
rect 388904 31748 388956 31754
rect 388904 31690 388956 31696
rect 388916 28830 388944 31690
rect 388720 28824 388772 28830
rect 388720 28766 388772 28772
rect 388904 28824 388956 28830
rect 388904 28766 388956 28772
rect 388732 12458 388760 28766
rect 388732 12430 388944 12458
rect 388916 8158 388944 12430
rect 388904 8152 388956 8158
rect 388904 8094 388956 8100
rect 388260 6452 388312 6458
rect 388260 6394 388312 6400
rect 387708 6044 387760 6050
rect 387708 5986 387760 5992
rect 386328 5908 386380 5914
rect 386328 5850 386380 5856
rect 387064 4684 387116 4690
rect 387064 4626 387116 4632
rect 385868 3732 385920 3738
rect 385868 3674 385920 3680
rect 385880 480 385908 3674
rect 387076 480 387104 4626
rect 388272 480 388300 6394
rect 389008 6118 389036 119734
rect 389824 118448 389876 118454
rect 389824 118390 389876 118396
rect 389088 117360 389140 117366
rect 389088 117302 389140 117308
rect 388996 6112 389048 6118
rect 388996 6054 389048 6060
rect 389100 3398 389128 117302
rect 389836 3806 389864 118390
rect 389928 118250 389956 120006
rect 389916 118244 389968 118250
rect 389916 118186 389968 118192
rect 390480 8090 390508 120006
rect 391124 117366 391152 120006
rect 391112 117360 391164 117366
rect 391112 117302 391164 117308
rect 391756 117360 391808 117366
rect 391756 117302 391808 117308
rect 390468 8084 390520 8090
rect 390468 8026 390520 8032
rect 391768 6866 391796 117302
rect 391756 6860 391808 6866
rect 391756 6802 391808 6808
rect 391860 6746 391888 120006
rect 392320 117366 392348 120006
rect 393148 118674 393176 120006
rect 393056 118646 393176 118674
rect 392308 117360 392360 117366
rect 392308 117302 392360 117308
rect 393056 109070 393084 118646
rect 393608 118522 393636 120006
rect 393596 118516 393648 118522
rect 393596 118458 393648 118464
rect 393964 117700 394016 117706
rect 393964 117642 394016 117648
rect 393136 117360 393188 117366
rect 393136 117302 393188 117308
rect 393044 109064 393096 109070
rect 393044 109006 393096 109012
rect 393148 8022 393176 117302
rect 393228 109064 393280 109070
rect 393228 109006 393280 109012
rect 393136 8016 393188 8022
rect 393136 7958 393188 7964
rect 393240 6798 393268 109006
rect 391768 6718 391888 6746
rect 393228 6792 393280 6798
rect 393228 6734 393280 6740
rect 390652 5500 390704 5506
rect 390652 5442 390704 5448
rect 389824 3800 389876 3806
rect 389824 3742 389876 3748
rect 389456 3664 389508 3670
rect 389456 3606 389508 3612
rect 389088 3392 389140 3398
rect 389088 3334 389140 3340
rect 389468 480 389496 3606
rect 390664 480 390692 5442
rect 391768 4146 391796 6718
rect 391848 6520 391900 6526
rect 391848 6462 391900 6468
rect 391756 4140 391808 4146
rect 391756 4082 391808 4088
rect 391860 480 391888 6462
rect 393044 3868 393096 3874
rect 393044 3810 393096 3816
rect 393056 480 393084 3810
rect 393976 3670 394004 117642
rect 394344 111058 394372 120006
rect 394344 111030 394464 111058
rect 394436 106282 394464 111030
rect 394424 106276 394476 106282
rect 394424 106218 394476 106224
rect 394424 99340 394476 99346
rect 394424 99282 394476 99288
rect 394436 96642 394464 99282
rect 394436 96614 394556 96642
rect 394528 89758 394556 96614
rect 394332 89752 394384 89758
rect 394516 89752 394568 89758
rect 394384 89700 394464 89706
rect 394332 89694 394464 89700
rect 394516 89694 394568 89700
rect 394344 89678 394464 89694
rect 394436 86970 394464 89678
rect 394424 86964 394476 86970
rect 394424 86906 394476 86912
rect 394516 77308 394568 77314
rect 394516 77250 394568 77256
rect 394528 67658 394556 77250
rect 394424 67652 394476 67658
rect 394424 67594 394476 67600
rect 394516 67652 394568 67658
rect 394516 67594 394568 67600
rect 394436 60738 394464 67594
rect 394436 60710 394556 60738
rect 394528 48346 394556 60710
rect 394424 48340 394476 48346
rect 394424 48282 394476 48288
rect 394516 48340 394568 48346
rect 394516 48282 394568 48288
rect 394436 41426 394464 48282
rect 394436 41398 394556 41426
rect 394528 29034 394556 41398
rect 394424 29028 394476 29034
rect 394424 28970 394476 28976
rect 394516 29028 394568 29034
rect 394516 28970 394568 28976
rect 394436 28914 394464 28970
rect 394436 28886 394556 28914
rect 394528 22302 394556 28886
rect 394516 22296 394568 22302
rect 394516 22238 394568 22244
rect 394424 22228 394476 22234
rect 394424 22170 394476 22176
rect 394436 19394 394464 22170
rect 394344 19366 394464 19394
rect 394344 19310 394372 19366
rect 394332 19304 394384 19310
rect 394332 19246 394384 19252
rect 394424 9716 394476 9722
rect 394424 9658 394476 9664
rect 394436 9602 394464 9658
rect 394344 9574 394464 9602
rect 394344 7954 394372 9574
rect 394332 7948 394384 7954
rect 394332 7890 394384 7896
rect 394620 6730 394648 120006
rect 395448 117366 395476 120006
rect 395436 117360 395488 117366
rect 395436 117302 395488 117308
rect 395908 7886 395936 120006
rect 396644 117366 396672 120006
rect 396724 118652 396776 118658
rect 396724 118594 396776 118600
rect 395988 117360 396040 117366
rect 395988 117302 396040 117308
rect 396632 117360 396684 117366
rect 396632 117302 396684 117308
rect 395896 7880 395948 7886
rect 395896 7822 395948 7828
rect 394608 6724 394660 6730
rect 394608 6666 394660 6672
rect 395436 6384 395488 6390
rect 395436 6326 395488 6332
rect 394240 4752 394292 4758
rect 394240 4694 394292 4700
rect 393964 3664 394016 3670
rect 393964 3606 394016 3612
rect 394252 480 394280 4694
rect 395448 480 395476 6326
rect 396000 4078 396028 117302
rect 395988 4072 396040 4078
rect 395988 4014 396040 4020
rect 396632 3936 396684 3942
rect 396632 3878 396684 3884
rect 396644 480 396672 3878
rect 396736 3738 396764 118594
rect 397288 118454 397316 120006
rect 397276 118448 397328 118454
rect 397276 118390 397328 118396
rect 397840 117366 397868 120006
rect 398104 117632 398156 117638
rect 398104 117574 398156 117580
rect 397368 117360 397420 117366
rect 397368 117302 397420 117308
rect 397828 117360 397880 117366
rect 397828 117302 397880 117308
rect 397380 6662 397408 117302
rect 397368 6656 397420 6662
rect 397368 6598 397420 6604
rect 397828 5432 397880 5438
rect 397828 5374 397880 5380
rect 396724 3732 396776 3738
rect 396724 3674 396776 3680
rect 397840 480 397868 5374
rect 398116 3602 398144 117574
rect 398668 6594 398696 120006
rect 399128 117366 399156 120006
rect 399680 117502 399708 120006
rect 400002 119762 400030 120020
rect 400568 120006 400904 120034
rect 401212 120006 401548 120034
rect 401856 120006 402192 120034
rect 402408 120006 402928 120034
rect 403052 120006 403388 120034
rect 399956 119734 400030 119762
rect 399668 117496 399720 117502
rect 399668 117438 399720 117444
rect 398748 117360 398800 117366
rect 398748 117302 398800 117308
rect 399116 117360 399168 117366
rect 399116 117302 399168 117308
rect 398656 6588 398708 6594
rect 398656 6530 398708 6536
rect 398760 4214 398788 117302
rect 399956 6526 399984 119734
rect 400876 118658 400904 120006
rect 400864 118652 400916 118658
rect 400864 118594 400916 118600
rect 400036 117496 400088 117502
rect 400036 117438 400088 117444
rect 399944 6520 399996 6526
rect 399944 6462 399996 6468
rect 399024 6248 399076 6254
rect 399024 6190 399076 6196
rect 398748 4208 398800 4214
rect 398748 4150 398800 4156
rect 398104 3596 398156 3602
rect 398104 3538 398156 3544
rect 399036 480 399064 6190
rect 400048 4282 400076 117438
rect 400128 117360 400180 117366
rect 400128 117302 400180 117308
rect 400036 4276 400088 4282
rect 400036 4218 400088 4224
rect 400140 4010 400168 117302
rect 401324 5364 401376 5370
rect 401324 5306 401376 5312
rect 400128 4004 400180 4010
rect 400128 3946 400180 3952
rect 400220 2848 400272 2854
rect 400220 2790 400272 2796
rect 400232 480 400260 2790
rect 401336 480 401364 5306
rect 401520 4418 401548 120006
rect 402164 117366 402192 120006
rect 402244 117768 402296 117774
rect 402244 117710 402296 117716
rect 402152 117360 402204 117366
rect 402152 117302 402204 117308
rect 401508 4412 401560 4418
rect 401508 4354 401560 4360
rect 402256 2854 402284 117710
rect 402796 117360 402848 117366
rect 402796 117302 402848 117308
rect 402808 6458 402836 117302
rect 402796 6452 402848 6458
rect 402796 6394 402848 6400
rect 402520 6316 402572 6322
rect 402520 6258 402572 6264
rect 402244 2848 402296 2854
rect 402244 2790 402296 2796
rect 402532 480 402560 6258
rect 402900 3942 402928 120006
rect 403360 117366 403388 120006
rect 403682 119762 403710 120020
rect 404234 119762 404262 120020
rect 404892 120006 405228 120034
rect 403682 119734 403756 119762
rect 404234 119734 404308 119762
rect 403348 117360 403400 117366
rect 403348 117302 403400 117308
rect 403728 116074 403756 119734
rect 404280 117706 404308 119734
rect 404268 117700 404320 117706
rect 404268 117642 404320 117648
rect 405200 117434 405228 120006
rect 405522 119762 405550 120020
rect 406088 120006 406424 120034
rect 406732 120006 406976 120034
rect 407376 120006 407712 120034
rect 407928 120006 408264 120034
rect 408572 120006 408908 120034
rect 409216 120006 409644 120034
rect 405522 119734 405596 119762
rect 405188 117428 405240 117434
rect 405188 117370 405240 117376
rect 404268 117360 404320 117366
rect 404268 117302 404320 117308
rect 403716 116068 403768 116074
rect 403716 116010 403768 116016
rect 403992 116068 404044 116074
rect 403992 116010 404044 116016
rect 404004 115938 404032 116010
rect 403992 115932 404044 115938
rect 403992 115874 404044 115880
rect 403900 106344 403952 106350
rect 403900 106286 403952 106292
rect 403912 99414 403940 106286
rect 403900 99408 403952 99414
rect 403900 99350 403952 99356
rect 403992 99340 404044 99346
rect 403992 99282 404044 99288
rect 404004 96626 404032 99282
rect 403992 96620 404044 96626
rect 403992 96562 404044 96568
rect 403900 87032 403952 87038
rect 403900 86974 403952 86980
rect 403912 79914 403940 86974
rect 403912 79886 404032 79914
rect 404004 77178 404032 79886
rect 403992 77172 404044 77178
rect 403992 77114 404044 77120
rect 404084 67652 404136 67658
rect 404084 67594 404136 67600
rect 404096 60858 404124 67594
rect 404084 60852 404136 60858
rect 404084 60794 404136 60800
rect 403992 60716 404044 60722
rect 403992 60658 404044 60664
rect 404004 57934 404032 60658
rect 403992 57928 404044 57934
rect 403992 57870 404044 57876
rect 404084 48340 404136 48346
rect 404084 48282 404136 48288
rect 404096 43466 404124 48282
rect 404004 43438 404124 43466
rect 404004 38622 404032 43438
rect 403992 38616 404044 38622
rect 403992 38558 404044 38564
rect 404084 29028 404136 29034
rect 404084 28970 404136 28976
rect 404096 22166 404124 28970
rect 404084 22160 404136 22166
rect 404084 22102 404136 22108
rect 403992 22092 404044 22098
rect 403992 22034 404044 22040
rect 404004 12458 404032 22034
rect 404004 12430 404216 12458
rect 404188 6390 404216 12430
rect 404176 6384 404228 6390
rect 404176 6326 404228 6332
rect 404280 4350 404308 117302
rect 405568 6254 405596 119734
rect 405648 117428 405700 117434
rect 405648 117370 405700 117376
rect 405556 6248 405608 6254
rect 405556 6190 405608 6196
rect 404912 5296 404964 5302
rect 404912 5238 404964 5244
rect 404268 4344 404320 4350
rect 404268 4286 404320 4292
rect 402888 3936 402940 3942
rect 402888 3878 402940 3884
rect 403716 3800 403768 3806
rect 403716 3742 403768 3748
rect 403728 480 403756 3742
rect 404924 480 404952 5238
rect 405660 4486 405688 117370
rect 406396 117366 406424 120006
rect 406384 117360 406436 117366
rect 406384 117302 406436 117308
rect 406108 6180 406160 6186
rect 406108 6122 406160 6128
rect 405648 4480 405700 4486
rect 405648 4422 405700 4428
rect 406120 480 406148 6122
rect 406948 4554 406976 120006
rect 407684 117366 407712 120006
rect 408236 117638 408264 120006
rect 408224 117632 408276 117638
rect 408224 117574 408276 117580
rect 408880 117502 408908 120006
rect 408868 117496 408920 117502
rect 408868 117438 408920 117444
rect 407028 117360 407080 117366
rect 407028 117302 407080 117308
rect 407672 117360 407724 117366
rect 407672 117302 407724 117308
rect 408408 117360 408460 117366
rect 408408 117302 408460 117308
rect 406936 4548 406988 4554
rect 406936 4490 406988 4496
rect 407040 3874 407068 117302
rect 408420 6322 408448 117302
rect 409512 9240 409564 9246
rect 409512 9182 409564 9188
rect 408408 6316 408460 6322
rect 408408 6258 408460 6264
rect 408684 5228 408736 5234
rect 408684 5170 408736 5176
rect 407028 3868 407080 3874
rect 407028 3810 407080 3816
rect 408314 3768 408370 3777
rect 408314 3703 408370 3712
rect 408498 3768 408554 3777
rect 408498 3703 408554 3712
rect 408328 3602 408356 3703
rect 408512 3602 408540 3703
rect 408316 3596 408368 3602
rect 408316 3538 408368 3544
rect 408500 3596 408552 3602
rect 408500 3538 408552 3544
rect 407304 3528 407356 3534
rect 408696 3482 408724 5170
rect 409524 3806 409552 9182
rect 409616 6186 409644 120006
rect 409754 119762 409782 120020
rect 410412 120006 410748 120034
rect 409754 119734 409828 119762
rect 409696 117496 409748 117502
rect 409696 117438 409748 117444
rect 409708 8514 409736 117438
rect 409800 9246 409828 119734
rect 410720 117434 410748 120006
rect 411042 119762 411070 120020
rect 411608 120006 411944 120034
rect 412252 120006 412588 120034
rect 412896 120006 413232 120034
rect 413448 120006 413784 120034
rect 414092 120006 414428 120034
rect 411042 119734 411116 119762
rect 410708 117428 410760 117434
rect 410708 117370 410760 117376
rect 409788 9240 409840 9246
rect 409788 9182 409840 9188
rect 409708 8486 409828 8514
rect 409696 7744 409748 7750
rect 409696 7686 409748 7692
rect 409604 6180 409656 6186
rect 409604 6122 409656 6128
rect 409512 3800 409564 3806
rect 409512 3742 409564 3748
rect 407304 3470 407356 3476
rect 407316 480 407344 3470
rect 408512 3454 408724 3482
rect 408512 480 408540 3454
rect 409708 480 409736 7686
rect 409800 4622 409828 8486
rect 411088 6225 411116 119734
rect 411916 117774 411944 120006
rect 411904 117768 411956 117774
rect 411904 117710 411956 117716
rect 411168 117428 411220 117434
rect 411168 117370 411220 117376
rect 411074 6216 411130 6225
rect 411074 6151 411130 6160
rect 411180 4690 411208 117370
rect 412088 5160 412140 5166
rect 412088 5102 412140 5108
rect 411168 4684 411220 4690
rect 411168 4626 411220 4632
rect 409788 4616 409840 4622
rect 409788 4558 409840 4564
rect 410892 3732 410944 3738
rect 410892 3674 410944 3680
rect 410904 480 410932 3674
rect 412100 480 412128 5102
rect 412560 4758 412588 120006
rect 413204 117366 413232 120006
rect 413284 117564 413336 117570
rect 413284 117506 413336 117512
rect 413192 117360 413244 117366
rect 413192 117302 413244 117308
rect 413296 10690 413324 117506
rect 413756 117434 413784 120006
rect 413744 117428 413796 117434
rect 413744 117370 413796 117376
rect 414400 117366 414428 120006
rect 413928 117360 413980 117366
rect 413928 117302 413980 117308
rect 414388 117360 414440 117366
rect 414388 117302 414440 117308
rect 413204 10662 413324 10690
rect 412548 4752 412600 4758
rect 412548 4694 412600 4700
rect 413204 3670 413232 10662
rect 413940 7818 413968 117302
rect 414860 115938 414888 120142
rect 415274 119762 415302 120020
rect 415932 120006 416268 120034
rect 415274 119734 415348 119762
rect 415320 117774 415348 119734
rect 415308 117768 415360 117774
rect 415308 117710 415360 117716
rect 416240 117434 416268 120006
rect 416562 119762 416590 120020
rect 417128 120006 417464 120034
rect 417772 120006 418108 120034
rect 418324 120006 418660 120034
rect 418968 120006 419304 120034
rect 419612 120006 419948 120034
rect 420164 120006 420316 120034
rect 416562 119734 416636 119762
rect 416044 117428 416096 117434
rect 416044 117370 416096 117376
rect 416228 117428 416280 117434
rect 416228 117370 416280 117376
rect 415308 117360 415360 117366
rect 415308 117302 415360 117308
rect 414848 115932 414900 115938
rect 414848 115874 414900 115880
rect 414940 115932 414992 115938
rect 414940 115874 414992 115880
rect 414952 108882 414980 115874
rect 414952 108854 415072 108882
rect 415044 104854 415072 108854
rect 415032 104848 415084 104854
rect 415032 104790 415084 104796
rect 415216 95260 415268 95266
rect 415216 95202 415268 95208
rect 415228 89826 415256 95202
rect 415216 89820 415268 89826
rect 415216 89762 415268 89768
rect 415124 89684 415176 89690
rect 415124 89626 415176 89632
rect 415136 75954 415164 89626
rect 415032 75948 415084 75954
rect 415032 75890 415084 75896
rect 415124 75948 415176 75954
rect 415124 75890 415176 75896
rect 415044 66230 415072 75890
rect 415032 66224 415084 66230
rect 415032 66166 415084 66172
rect 415032 56636 415084 56642
rect 415032 56578 415084 56584
rect 415044 51338 415072 56578
rect 415032 51332 415084 51338
rect 415032 51274 415084 51280
rect 415216 51332 415268 51338
rect 415216 51274 415268 51280
rect 415228 48385 415256 51274
rect 415030 48376 415086 48385
rect 414952 48334 415030 48362
rect 414952 45558 414980 48334
rect 415030 48311 415086 48320
rect 415214 48376 415270 48385
rect 415214 48311 415270 48320
rect 414940 45552 414992 45558
rect 414940 45494 414992 45500
rect 415032 35964 415084 35970
rect 415032 35906 415084 35912
rect 415044 26246 415072 35906
rect 415032 26240 415084 26246
rect 415032 26182 415084 26188
rect 415032 16652 415084 16658
rect 415032 16594 415084 16600
rect 415044 12510 415072 16594
rect 415032 12504 415084 12510
rect 415032 12446 415084 12452
rect 414940 12436 414992 12442
rect 414940 12378 414992 12384
rect 413928 7812 413980 7818
rect 413928 7754 413980 7760
rect 414952 7750 414980 12378
rect 414940 7744 414992 7750
rect 414940 7686 414992 7692
rect 413284 7676 413336 7682
rect 413284 7618 413336 7624
rect 413192 3664 413244 3670
rect 413192 3606 413244 3612
rect 413296 480 413324 7618
rect 415320 5506 415348 117302
rect 415308 5500 415360 5506
rect 415308 5442 415360 5448
rect 415676 5092 415728 5098
rect 415676 5034 415728 5040
rect 414480 2984 414532 2990
rect 414480 2926 414532 2932
rect 414492 480 414520 2926
rect 415688 480 415716 5034
rect 416056 2990 416084 117370
rect 416608 7682 416636 119734
rect 416780 117836 416832 117842
rect 416780 117778 416832 117784
rect 416688 117428 416740 117434
rect 416688 117370 416740 117376
rect 416596 7676 416648 7682
rect 416596 7618 416648 7624
rect 416700 5438 416728 117370
rect 416792 7614 416820 117778
rect 417436 117570 417464 120006
rect 417424 117564 417476 117570
rect 417424 117506 417476 117512
rect 416780 7608 416832 7614
rect 416780 7550 416832 7556
rect 417976 7608 418028 7614
rect 417976 7550 418028 7556
rect 416872 7064 416924 7070
rect 416872 7006 416924 7012
rect 416688 5432 416740 5438
rect 416688 5374 416740 5380
rect 416044 2984 416096 2990
rect 416044 2926 416096 2932
rect 416884 480 416912 7006
rect 417882 3632 417938 3641
rect 417882 3567 417938 3576
rect 417896 3534 417924 3567
rect 417884 3528 417936 3534
rect 417884 3470 417936 3476
rect 417988 480 418016 7550
rect 418080 5370 418108 120006
rect 418632 117434 418660 120006
rect 419276 117842 419304 120006
rect 419264 117836 419316 117842
rect 419264 117778 419316 117784
rect 419920 117434 419948 120006
rect 420184 117836 420236 117842
rect 420184 117778 420236 117784
rect 418620 117428 418672 117434
rect 418620 117370 418672 117376
rect 419448 117428 419500 117434
rect 419448 117370 419500 117376
rect 419908 117428 419960 117434
rect 419908 117370 419960 117376
rect 419460 9450 419488 117370
rect 419448 9444 419500 9450
rect 419448 9386 419500 9392
rect 418068 5364 418120 5370
rect 418068 5306 418120 5312
rect 419172 5024 419224 5030
rect 419172 4966 419224 4972
rect 418160 3732 418212 3738
rect 418160 3674 418212 3680
rect 418172 2990 418200 3674
rect 418342 3632 418398 3641
rect 418342 3567 418398 3576
rect 418356 3466 418384 3567
rect 418344 3460 418396 3466
rect 418344 3402 418396 3408
rect 418160 2984 418212 2990
rect 418160 2926 418212 2932
rect 419184 480 419212 4966
rect 420196 3670 420224 117778
rect 420288 116006 420316 120006
rect 420794 119762 420822 120020
rect 421452 120006 421788 120034
rect 422004 120006 422156 120034
rect 422648 120006 422984 120034
rect 423292 120006 423628 120034
rect 423844 120006 424180 120034
rect 424488 120006 425008 120034
rect 425132 120006 425468 120034
rect 425684 120006 425928 120034
rect 420794 119734 420868 119762
rect 420840 117570 420868 119734
rect 420828 117564 420880 117570
rect 420828 117506 420880 117512
rect 421760 117434 421788 120006
rect 420828 117428 420880 117434
rect 420828 117370 420880 117376
rect 421748 117428 421800 117434
rect 421748 117370 421800 117376
rect 420276 116000 420328 116006
rect 420276 115942 420328 115948
rect 420460 116000 420512 116006
rect 420460 115942 420512 115948
rect 420472 115870 420500 115942
rect 420460 115864 420512 115870
rect 420460 115806 420512 115812
rect 420644 108996 420696 109002
rect 420644 108938 420696 108944
rect 420656 104854 420684 108938
rect 420644 104848 420696 104854
rect 420644 104790 420696 104796
rect 420644 95260 420696 95266
rect 420644 95202 420696 95208
rect 420656 89758 420684 95202
rect 420644 89752 420696 89758
rect 420644 89694 420696 89700
rect 420644 89616 420696 89622
rect 420644 89558 420696 89564
rect 420656 82142 420684 89558
rect 420276 82136 420328 82142
rect 420276 82078 420328 82084
rect 420644 82136 420696 82142
rect 420644 82078 420696 82084
rect 420288 77353 420316 82078
rect 420274 77344 420330 77353
rect 420274 77279 420330 77288
rect 420458 77344 420514 77353
rect 420514 77302 420592 77330
rect 420458 77279 420514 77288
rect 420564 66298 420592 77302
rect 420460 66292 420512 66298
rect 420460 66234 420512 66240
rect 420552 66292 420604 66298
rect 420552 66234 420604 66240
rect 420472 66162 420500 66234
rect 420460 66156 420512 66162
rect 420460 66098 420512 66104
rect 420644 66156 420696 66162
rect 420644 66098 420696 66104
rect 420656 61441 420684 66098
rect 420642 61432 420698 61441
rect 420642 61367 420698 61376
rect 420550 48376 420606 48385
rect 420472 48334 420550 48362
rect 420472 46918 420500 48334
rect 420550 48311 420606 48320
rect 420460 46912 420512 46918
rect 420460 46854 420512 46860
rect 420644 46912 420696 46918
rect 420644 46854 420696 46860
rect 420656 42129 420684 46854
rect 420642 42120 420698 42129
rect 420642 42055 420698 42064
rect 420550 29064 420606 29073
rect 420472 29022 420550 29050
rect 420472 27606 420500 29022
rect 420550 28999 420606 29008
rect 420460 27600 420512 27606
rect 420460 27542 420512 27548
rect 420552 18012 420604 18018
rect 420552 17954 420604 17960
rect 420564 12510 420592 17954
rect 420552 12504 420604 12510
rect 420552 12446 420604 12452
rect 420460 12436 420512 12442
rect 420460 12378 420512 12384
rect 420472 9382 420500 12378
rect 420460 9376 420512 9382
rect 420460 9318 420512 9324
rect 420368 9172 420420 9178
rect 420368 9114 420420 9120
rect 420184 3664 420236 3670
rect 420184 3606 420236 3612
rect 420380 480 420408 9114
rect 420840 5302 420868 117370
rect 422128 9314 422156 120006
rect 422956 117774 422984 120006
rect 422944 117768 422996 117774
rect 422944 117710 422996 117716
rect 422208 117428 422260 117434
rect 422208 117370 422260 117376
rect 422116 9308 422168 9314
rect 422116 9250 422168 9256
rect 420828 5296 420880 5302
rect 420828 5238 420880 5244
rect 422220 5234 422248 117370
rect 422208 5228 422260 5234
rect 422208 5170 422260 5176
rect 423600 5166 423628 120006
rect 424152 117434 424180 120006
rect 424980 117994 425008 120006
rect 424980 117966 425192 117994
rect 425164 117910 425192 117966
rect 425060 117904 425112 117910
rect 425060 117846 425112 117852
rect 425152 117904 425204 117910
rect 425152 117846 425204 117852
rect 424324 117768 424376 117774
rect 424324 117710 424376 117716
rect 424140 117428 424192 117434
rect 424140 117370 424192 117376
rect 423956 9104 424008 9110
rect 423956 9046 424008 9052
rect 423588 5160 423640 5166
rect 423588 5102 423640 5108
rect 422760 4888 422812 4894
rect 422760 4830 422812 4836
rect 421564 3528 421616 3534
rect 421564 3470 421616 3476
rect 421576 480 421604 3470
rect 422772 480 422800 4830
rect 423968 480 423996 9046
rect 424336 3602 424364 117710
rect 424968 117428 425020 117434
rect 424968 117370 425020 117376
rect 424980 9246 425008 117370
rect 424968 9240 425020 9246
rect 424968 9182 425020 9188
rect 424324 3596 424376 3602
rect 424324 3538 424376 3544
rect 425072 626 425100 117846
rect 425440 117434 425468 120006
rect 425428 117428 425480 117434
rect 425428 117370 425480 117376
rect 425900 116006 425928 120006
rect 426314 119762 426342 120020
rect 426972 120006 427308 120034
rect 427524 120006 427676 120034
rect 428168 120006 428504 120034
rect 428812 120006 429148 120034
rect 429364 120006 429700 120034
rect 430008 120006 430344 120034
rect 430652 120006 430988 120034
rect 431204 120006 431356 120034
rect 426314 119734 426388 119762
rect 426360 117774 426388 119734
rect 426348 117768 426400 117774
rect 426348 117710 426400 117716
rect 427280 117570 427308 120006
rect 427268 117564 427320 117570
rect 427268 117506 427320 117512
rect 426348 117428 426400 117434
rect 426348 117370 426400 117376
rect 425888 116000 425940 116006
rect 425888 115942 425940 115948
rect 425980 116000 426032 116006
rect 425980 115942 426032 115948
rect 425992 109018 426020 115942
rect 425992 108990 426204 109018
rect 426176 96642 426204 108990
rect 426176 96614 426296 96642
rect 426268 95198 426296 96614
rect 426256 95192 426308 95198
rect 426256 95134 426308 95140
rect 426164 85604 426216 85610
rect 426164 85546 426216 85552
rect 426176 84182 426204 85546
rect 426164 84176 426216 84182
rect 426164 84118 426216 84124
rect 426072 69692 426124 69698
rect 426072 69634 426124 69640
rect 426084 53174 426112 69634
rect 426072 53168 426124 53174
rect 426072 53110 426124 53116
rect 426256 53168 426308 53174
rect 426256 53110 426308 53116
rect 426268 48385 426296 53110
rect 426070 48376 426126 48385
rect 425992 48334 426070 48362
rect 425992 46918 426020 48334
rect 426070 48311 426126 48320
rect 426254 48376 426310 48385
rect 426254 48311 426310 48320
rect 425980 46912 426032 46918
rect 425980 46854 426032 46860
rect 426072 37324 426124 37330
rect 426072 37266 426124 37272
rect 426084 19310 426112 37266
rect 425980 19304 426032 19310
rect 425980 19246 426032 19252
rect 426072 19304 426124 19310
rect 426072 19246 426124 19252
rect 425992 9178 426020 19246
rect 425980 9172 426032 9178
rect 425980 9114 426032 9120
rect 426360 5098 426388 117370
rect 427648 9110 427676 120006
rect 428476 118726 428504 120006
rect 428464 118720 428516 118726
rect 428464 118662 428516 118668
rect 427728 117564 427780 117570
rect 427728 117506 427780 117512
rect 427636 9104 427688 9110
rect 427636 9046 427688 9052
rect 427544 9036 427596 9042
rect 427544 8978 427596 8984
rect 426348 5092 426400 5098
rect 426348 5034 426400 5040
rect 426348 4956 426400 4962
rect 426348 4898 426400 4904
rect 425072 598 425192 626
rect 425164 480 425192 598
rect 426360 480 426388 4898
rect 427556 480 427584 8978
rect 427740 5030 427768 117506
rect 427728 5024 427780 5030
rect 427728 4966 427780 4972
rect 429120 4962 429148 120006
rect 429672 117502 429700 120006
rect 430316 117570 430344 120006
rect 429844 117564 429896 117570
rect 429844 117506 429896 117512
rect 430304 117564 430356 117570
rect 430304 117506 430356 117512
rect 429660 117496 429712 117502
rect 429660 117438 429712 117444
rect 429108 4956 429160 4962
rect 429108 4898 429160 4904
rect 429856 2922 429884 117506
rect 430960 117502 430988 120006
rect 431224 117564 431276 117570
rect 431224 117506 431276 117512
rect 430488 117496 430540 117502
rect 430488 117438 430540 117444
rect 430948 117496 431000 117502
rect 430948 117438 431000 117444
rect 430500 7614 430528 117438
rect 431132 8968 431184 8974
rect 431132 8910 431184 8916
rect 430488 7608 430540 7614
rect 430488 7550 430540 7556
rect 429936 4820 429988 4826
rect 429936 4762 429988 4768
rect 428740 2916 428792 2922
rect 428740 2858 428792 2864
rect 429844 2916 429896 2922
rect 429844 2858 429896 2864
rect 428752 480 428780 2858
rect 429948 480 429976 4762
rect 431144 480 431172 8910
rect 431236 3369 431264 117506
rect 431328 116006 431356 120006
rect 431834 119762 431862 120020
rect 432492 120006 432828 120034
rect 433044 120006 433196 120034
rect 433688 120006 434024 120034
rect 431788 119734 431862 119762
rect 431788 117570 431816 119734
rect 431776 117564 431828 117570
rect 431776 117506 431828 117512
rect 432800 117502 432828 120006
rect 431868 117496 431920 117502
rect 431868 117438 431920 117444
rect 432788 117496 432840 117502
rect 432788 117438 432840 117444
rect 431316 116000 431368 116006
rect 431316 115942 431368 115948
rect 431500 116000 431552 116006
rect 431500 115942 431552 115948
rect 431512 109018 431540 115942
rect 431512 108990 431724 109018
rect 431696 106282 431724 108990
rect 431684 106276 431736 106282
rect 431684 106218 431736 106224
rect 431684 99340 431736 99346
rect 431684 99282 431736 99288
rect 431696 96642 431724 99282
rect 431696 96614 431816 96642
rect 431788 87009 431816 96614
rect 431590 87000 431646 87009
rect 431590 86935 431646 86944
rect 431774 87000 431830 87009
rect 431774 86935 431830 86944
rect 431604 80102 431632 86935
rect 431788 80102 431816 80133
rect 431592 80096 431644 80102
rect 431776 80096 431828 80102
rect 431644 80044 431776 80050
rect 431592 80038 431828 80044
rect 431604 80022 431816 80038
rect 431604 75886 431632 80022
rect 431592 75880 431644 75886
rect 431592 75822 431644 75828
rect 431592 66292 431644 66298
rect 431592 66234 431644 66240
rect 431604 56574 431632 66234
rect 431592 56568 431644 56574
rect 431592 56510 431644 56516
rect 431776 56568 431828 56574
rect 431776 56510 431828 56516
rect 431788 47025 431816 56510
rect 431590 47016 431646 47025
rect 431590 46951 431646 46960
rect 431774 47016 431830 47025
rect 431774 46951 431830 46960
rect 431604 46918 431632 46951
rect 431592 46912 431644 46918
rect 431592 46854 431644 46860
rect 431592 37324 431644 37330
rect 431592 37266 431644 37272
rect 431604 37194 431632 37266
rect 431592 37188 431644 37194
rect 431592 37130 431644 37136
rect 431684 31680 431736 31686
rect 431684 31622 431736 31628
rect 431696 26246 431724 31622
rect 431684 26240 431736 26246
rect 431684 26182 431736 26188
rect 431500 16652 431552 16658
rect 431500 16594 431552 16600
rect 431512 9042 431540 16594
rect 431500 9036 431552 9042
rect 431500 8978 431552 8984
rect 431880 4894 431908 117438
rect 433168 8974 433196 120006
rect 433996 118017 434024 120006
rect 433982 118008 434038 118017
rect 433982 117943 434038 117952
rect 433248 117496 433300 117502
rect 433248 117438 433300 117444
rect 433156 8968 433208 8974
rect 433156 8910 433208 8916
rect 431868 4888 431920 4894
rect 431868 4830 431920 4836
rect 433260 4826 433288 117438
rect 435008 80034 435036 196143
rect 435100 188873 435128 251194
rect 435180 207052 435232 207058
rect 435180 206994 435232 207000
rect 435192 190233 435220 206994
rect 435178 190224 435234 190233
rect 435178 190159 435234 190168
rect 435086 188864 435142 188873
rect 435086 188799 435142 188808
rect 436112 180305 436140 355302
rect 436560 201136 436612 201142
rect 436560 201078 436612 201084
rect 436468 201068 436520 201074
rect 436468 201010 436520 201016
rect 436376 201000 436428 201006
rect 436376 200942 436428 200948
rect 436190 198928 436246 198937
rect 436190 198863 436246 198872
rect 436098 180296 436154 180305
rect 436098 180231 436154 180240
rect 436100 155236 436152 155242
rect 436100 155178 436152 155184
rect 436112 155145 436140 155178
rect 436098 155136 436154 155145
rect 436098 155071 436154 155080
rect 436100 149048 436152 149054
rect 436100 148990 436152 148996
rect 436112 148753 436140 148990
rect 436098 148744 436154 148753
rect 436098 148679 436154 148688
rect 436100 142112 436152 142118
rect 436098 142080 436100 142089
rect 436152 142080 436154 142089
rect 436098 142015 436154 142024
rect 434996 80028 435048 80034
rect 434996 79970 435048 79976
rect 436204 35902 436232 198863
rect 436282 194032 436338 194041
rect 436282 193967 436338 193976
rect 436296 121038 436324 193967
rect 436388 176225 436416 200942
rect 436480 177993 436508 201010
rect 436572 182073 436600 201078
rect 436652 200184 436704 200190
rect 436652 200126 436704 200132
rect 436664 193089 436692 200126
rect 436650 193080 436706 193089
rect 436650 193015 436706 193024
rect 436558 182064 436614 182073
rect 436558 181999 436614 182008
rect 436466 177984 436522 177993
rect 436466 177919 436522 177928
rect 436374 176216 436430 176225
rect 436374 176151 436430 176160
rect 436756 140457 436784 438874
rect 436836 157412 436888 157418
rect 436836 157354 436888 157360
rect 436742 140448 436798 140457
rect 436742 140383 436798 140392
rect 436848 127809 436876 157354
rect 438136 155242 438164 700402
rect 462332 700398 462360 703520
rect 478524 700505 478552 703520
rect 478510 700496 478566 700505
rect 494808 700466 494836 703520
rect 478510 700431 478566 700440
rect 494796 700460 494848 700466
rect 494796 700402 494848 700408
rect 462320 700392 462372 700398
rect 462320 700334 462372 700340
rect 447784 700324 447836 700330
rect 447784 700266 447836 700272
rect 446404 673532 446456 673538
rect 446404 673474 446456 673480
rect 445024 626612 445076 626618
rect 445024 626554 445076 626560
rect 442264 579692 442316 579698
rect 442264 579634 442316 579640
rect 438216 485852 438268 485858
rect 438216 485794 438268 485800
rect 438124 155236 438176 155242
rect 438124 155178 438176 155184
rect 437388 153196 437440 153202
rect 437388 153138 437440 153144
rect 437400 152833 437428 153138
rect 437386 152824 437442 152833
rect 437386 152759 437442 152768
rect 437388 150408 437440 150414
rect 437388 150350 437440 150356
rect 437400 150249 437428 150350
rect 437386 150240 437442 150249
rect 437386 150175 437442 150184
rect 437386 146296 437442 146305
rect 437386 146231 437442 146240
rect 437400 146198 437428 146231
rect 437388 146192 437440 146198
rect 437388 146134 437440 146140
rect 437020 144900 437072 144906
rect 437020 144842 437072 144848
rect 437032 144537 437060 144842
rect 437018 144528 437074 144537
rect 437018 144463 437074 144472
rect 438228 142118 438256 485794
rect 442276 146198 442304 579634
rect 445036 149054 445064 626554
rect 446416 150414 446444 673474
rect 447796 153202 447824 700266
rect 484400 556300 484452 556306
rect 484400 556242 484452 556248
rect 484412 554676 484440 556242
rect 511264 556232 511316 556238
rect 511264 556174 511316 556180
rect 511276 554676 511304 556174
rect 514024 532772 514076 532778
rect 514024 532714 514076 532720
rect 479996 518294 480024 520132
rect 479984 518288 480036 518294
rect 479984 518230 480036 518236
rect 506860 518226 506888 520132
rect 506848 518220 506900 518226
rect 506848 518162 506900 518168
rect 464252 389428 464304 389434
rect 464252 389370 464304 389376
rect 464264 387532 464292 389370
rect 487436 389360 487488 389366
rect 487436 389302 487488 389308
rect 475844 389292 475896 389298
rect 475844 389234 475896 389240
rect 475856 387532 475884 389234
rect 487448 387532 487476 389302
rect 499028 389224 499080 389230
rect 499028 389166 499080 389172
rect 499040 387532 499068 389166
rect 504730 378448 504786 378457
rect 503732 378406 504730 378434
rect 456798 375184 456854 375193
rect 456798 375119 456854 375128
rect 456812 374066 456840 375119
rect 456800 374060 456852 374066
rect 456800 374002 456852 374008
rect 503732 361434 503760 378406
rect 504730 378383 504786 378392
rect 503640 361406 503760 361434
rect 503640 360074 503668 361406
rect 504730 360496 504786 360505
rect 504376 360454 504730 360482
rect 503640 360046 503760 360074
rect 503732 359938 503760 360046
rect 503732 359910 503852 359938
rect 456798 358048 456854 358057
rect 456798 357983 456854 357992
rect 456812 357474 456840 357983
rect 456800 357468 456852 357474
rect 456800 357410 456852 357416
rect 503824 350554 503852 359910
rect 504376 351914 504404 360454
rect 504730 360431 504786 360440
rect 504100 351886 504404 351914
rect 504100 350554 504128 351886
rect 503824 350526 504036 350554
rect 504100 350526 504220 350554
rect 504008 344978 504036 350526
rect 503916 344950 504036 344978
rect 503812 342032 503864 342038
rect 503812 341974 503864 341980
rect 503718 340912 503774 340921
rect 503718 340847 503774 340856
rect 460584 337618 460612 340068
rect 460572 337612 460624 337618
rect 460572 337554 460624 337560
rect 472176 337550 472204 340068
rect 472164 337544 472216 337550
rect 472164 337486 472216 337492
rect 483768 337482 483796 340068
rect 483756 337476 483808 337482
rect 483756 337418 483808 337424
rect 495360 337414 495388 340068
rect 495348 337408 495400 337414
rect 495348 337350 495400 337356
rect 503536 333328 503588 333334
rect 503536 333270 503588 333276
rect 503548 328522 503576 333270
rect 503732 331378 503760 340847
rect 503824 333334 503852 341974
rect 503916 340921 503944 344950
rect 504192 342038 504220 350526
rect 504824 345092 504876 345098
rect 504824 345034 504876 345040
rect 504730 343632 504786 343641
rect 504730 343567 504786 343576
rect 504180 342032 504232 342038
rect 504180 341974 504232 341980
rect 503902 340912 503958 340921
rect 504744 340882 504772 343567
rect 503902 340847 503958 340856
rect 504732 340876 504784 340882
rect 504732 340818 504784 340824
rect 503904 340808 503956 340814
rect 503904 340750 503956 340756
rect 503812 333328 503864 333334
rect 503812 333270 503864 333276
rect 503640 331350 503760 331378
rect 503640 331226 503668 331350
rect 503628 331220 503680 331226
rect 503628 331162 503680 331168
rect 503548 328494 503760 328522
rect 503732 321858 503760 328494
rect 503640 321830 503760 321858
rect 503640 318866 503668 321830
rect 503916 321774 503944 340750
rect 504836 333334 504864 345034
rect 504364 333328 504416 333334
rect 504364 333270 504416 333276
rect 504824 333328 504876 333334
rect 504824 333270 504876 333276
rect 503996 331220 504048 331226
rect 503996 331162 504048 331168
rect 503904 321768 503956 321774
rect 503904 321710 503956 321716
rect 504008 321706 504036 331162
rect 503996 321700 504048 321706
rect 503996 321642 504048 321648
rect 503904 321564 503956 321570
rect 503904 321506 503956 321512
rect 503640 318838 503760 318866
rect 503732 318782 503760 318838
rect 503720 318776 503772 318782
rect 503720 318718 503772 318724
rect 503628 311908 503680 311914
rect 503628 311850 503680 311856
rect 503640 311778 503668 311850
rect 503628 311772 503680 311778
rect 503628 311714 503680 311720
rect 503812 309188 503864 309194
rect 503812 309130 503864 309136
rect 503824 292482 503852 309130
rect 503732 292454 503852 292482
rect 503732 283082 503760 292454
rect 503720 283076 503772 283082
rect 503720 283018 503772 283024
rect 503812 283008 503864 283014
rect 503812 282950 503864 282956
rect 503628 273352 503680 273358
rect 503628 273294 503680 273300
rect 503640 273222 503668 273294
rect 503628 273216 503680 273222
rect 503628 273158 503680 273164
rect 503720 263696 503772 263702
rect 503720 263638 503772 263644
rect 503732 263566 503760 263638
rect 503720 263560 503772 263566
rect 503720 263502 503772 263508
rect 503628 254040 503680 254046
rect 503628 253982 503680 253988
rect 503640 253910 503668 253982
rect 503628 253904 503680 253910
rect 503824 253858 503852 282950
rect 503628 253846 503680 253852
rect 503732 253830 503852 253858
rect 503732 244458 503760 253830
rect 503720 244452 503772 244458
rect 503720 244394 503772 244400
rect 503812 244384 503864 244390
rect 503812 244326 503864 244332
rect 503628 234728 503680 234734
rect 503628 234670 503680 234676
rect 503640 234598 503668 234670
rect 503628 234592 503680 234598
rect 503824 234546 503852 244326
rect 503628 234534 503680 234540
rect 503732 234518 503852 234546
rect 503732 225146 503760 234518
rect 503720 225140 503772 225146
rect 503720 225082 503772 225088
rect 503812 225072 503864 225078
rect 503812 225014 503864 225020
rect 503628 215416 503680 215422
rect 503628 215358 503680 215364
rect 503640 215286 503668 215358
rect 503628 215280 503680 215286
rect 503824 215234 503852 225014
rect 503628 215222 503680 215228
rect 503732 215206 503852 215234
rect 503732 205834 503760 215206
rect 503720 205828 503772 205834
rect 503720 205770 503772 205776
rect 503812 205760 503864 205766
rect 503812 205702 503864 205708
rect 503720 205692 503772 205698
rect 503720 205634 503772 205640
rect 503732 202162 503760 205634
rect 503824 202230 503852 205702
rect 503916 202298 503944 321506
rect 503996 318844 504048 318850
rect 503996 318786 504048 318792
rect 504008 311914 504036 318786
rect 503996 311908 504048 311914
rect 503996 311850 504048 311856
rect 503996 311772 504048 311778
rect 503996 311714 504048 311720
rect 504008 273358 504036 311714
rect 504376 309346 504404 333270
rect 504376 309318 504496 309346
rect 504468 309210 504496 309318
rect 504376 309182 504496 309210
rect 504376 309126 504404 309182
rect 504364 309120 504416 309126
rect 504364 309062 504416 309068
rect 504456 299532 504508 299538
rect 504456 299474 504508 299480
rect 504468 292602 504496 299474
rect 504272 292596 504324 292602
rect 504272 292538 504324 292544
rect 504456 292596 504508 292602
rect 504456 292538 504508 292544
rect 504284 288454 504312 292538
rect 504272 288448 504324 288454
rect 504272 288390 504324 288396
rect 504456 280288 504508 280294
rect 504456 280230 504508 280236
rect 504468 278730 504496 280230
rect 504456 278724 504508 278730
rect 504456 278666 504508 278672
rect 503996 273352 504048 273358
rect 503996 273294 504048 273300
rect 503996 273216 504048 273222
rect 503996 273158 504048 273164
rect 504008 263702 504036 273158
rect 504640 269136 504692 269142
rect 504640 269078 504692 269084
rect 503996 263696 504048 263702
rect 503996 263638 504048 263644
rect 503996 263560 504048 263566
rect 503996 263502 504048 263508
rect 504008 254046 504036 263502
rect 504652 260953 504680 269078
rect 504270 260944 504326 260953
rect 504270 260879 504326 260888
rect 504638 260944 504694 260953
rect 504638 260879 504694 260888
rect 504284 260846 504312 260879
rect 504272 260840 504324 260846
rect 504272 260782 504324 260788
rect 503996 254040 504048 254046
rect 503996 253982 504048 253988
rect 503996 253904 504048 253910
rect 503996 253846 504048 253852
rect 504008 234734 504036 253846
rect 504272 253836 504324 253842
rect 504272 253778 504324 253784
rect 504284 251190 504312 253778
rect 504272 251184 504324 251190
rect 504272 251126 504324 251132
rect 504456 241528 504508 241534
rect 504456 241470 504508 241476
rect 504468 234734 504496 241470
rect 503996 234728 504048 234734
rect 503996 234670 504048 234676
rect 504456 234728 504508 234734
rect 504456 234670 504508 234676
rect 503996 234592 504048 234598
rect 503996 234534 504048 234540
rect 504364 234592 504416 234598
rect 504364 234534 504416 234540
rect 504008 215422 504036 234534
rect 504376 231810 504404 234534
rect 504364 231804 504416 231810
rect 504364 231746 504416 231752
rect 504456 222216 504508 222222
rect 504456 222158 504508 222164
rect 504468 215422 504496 222158
rect 503996 215416 504048 215422
rect 503996 215358 504048 215364
rect 504456 215416 504508 215422
rect 504456 215358 504508 215364
rect 503996 215280 504048 215286
rect 503996 215222 504048 215228
rect 504272 215280 504324 215286
rect 504272 215222 504324 215228
rect 504008 205698 504036 215222
rect 504284 212514 504312 215222
rect 504192 212486 504312 212514
rect 504192 205698 504220 212486
rect 503996 205692 504048 205698
rect 503996 205634 504048 205640
rect 504180 205692 504232 205698
rect 504180 205634 504232 205640
rect 504180 202904 504232 202910
rect 504180 202846 504232 202852
rect 504192 202774 504220 202846
rect 504180 202768 504232 202774
rect 504180 202710 504232 202716
rect 504456 202768 504508 202774
rect 504456 202710 504508 202716
rect 503904 202292 503956 202298
rect 503904 202234 503956 202240
rect 503812 202224 503864 202230
rect 503812 202166 503864 202172
rect 503720 202156 503772 202162
rect 503720 202098 503772 202104
rect 504468 186266 504496 202710
rect 504376 186238 504496 186266
rect 504376 183569 504404 186238
rect 504362 183560 504418 183569
rect 504362 183495 504418 183504
rect 504638 183560 504694 183569
rect 504638 183495 504694 183504
rect 504652 173942 504680 183495
rect 504456 173936 504508 173942
rect 504456 173878 504508 173884
rect 504640 173936 504692 173942
rect 504640 173878 504692 173884
rect 504468 166954 504496 173878
rect 504376 166926 504496 166954
rect 504376 164218 504404 166926
rect 504180 164212 504232 164218
rect 504180 164154 504232 164160
rect 504364 164212 504416 164218
rect 504364 164154 504416 164160
rect 504192 154601 504220 164154
rect 504178 154592 504234 154601
rect 504178 154527 504234 154536
rect 504454 154592 504510 154601
rect 504454 154527 504510 154536
rect 447784 153196 447836 153202
rect 447784 153138 447836 153144
rect 446404 150408 446456 150414
rect 446404 150350 446456 150356
rect 445024 149048 445076 149054
rect 445024 148990 445076 148996
rect 442264 146192 442316 146198
rect 442264 146134 442316 146140
rect 438216 142112 438268 142118
rect 438216 142054 438268 142060
rect 437388 137964 437440 137970
rect 437388 137906 437440 137912
rect 437400 137873 437428 137906
rect 437386 137864 437442 137873
rect 437386 137799 437442 137808
rect 504468 136610 504496 154527
rect 514036 144906 514064 532714
rect 527192 200705 527220 703520
rect 543476 700369 543504 703520
rect 543462 700360 543518 700369
rect 559668 700330 559696 703520
rect 543462 700295 543518 700304
rect 559656 700324 559708 700330
rect 559656 700266 559708 700272
rect 580170 674656 580226 674665
rect 580170 674591 580226 674600
rect 580184 673538 580212 674591
rect 580172 673532 580224 673538
rect 580172 673474 580224 673480
rect 580170 627736 580226 627745
rect 580170 627671 580226 627680
rect 580184 626618 580212 627671
rect 580172 626612 580224 626618
rect 580172 626554 580224 626560
rect 580170 580816 580226 580825
rect 580170 580751 580226 580760
rect 580184 579698 580212 580751
rect 580172 579692 580224 579698
rect 580172 579634 580224 579640
rect 580262 557288 580318 557297
rect 580262 557223 580318 557232
rect 580170 533896 580226 533905
rect 580170 533831 580226 533840
rect 580184 532778 580212 533831
rect 580172 532772 580224 532778
rect 580172 532714 580224 532720
rect 580170 498672 580226 498681
rect 580170 498607 580226 498616
rect 580184 498234 580212 498607
rect 580172 498228 580224 498234
rect 580172 498170 580224 498176
rect 580170 486840 580226 486849
rect 580170 486775 580226 486784
rect 580184 485858 580212 486775
rect 580172 485852 580224 485858
rect 580172 485794 580224 485800
rect 579802 463448 579858 463457
rect 579802 463383 579858 463392
rect 579816 462398 579844 463383
rect 579804 462392 579856 462398
rect 579804 462334 579856 462340
rect 580170 451752 580226 451761
rect 580170 451687 580226 451696
rect 580184 451314 580212 451687
rect 580172 451308 580224 451314
rect 580172 451250 580224 451256
rect 580170 439920 580226 439929
rect 580170 439855 580226 439864
rect 580184 438938 580212 439855
rect 580172 438932 580224 438938
rect 580172 438874 580224 438880
rect 579802 416528 579858 416537
rect 579802 416463 579858 416472
rect 579816 415478 579844 416463
rect 579804 415472 579856 415478
rect 579804 415414 579856 415420
rect 579986 346080 580042 346089
rect 579986 346015 580042 346024
rect 580000 345098 580028 346015
rect 579988 345092 580040 345098
rect 579988 345034 580040 345040
rect 579618 322688 579674 322697
rect 579618 322623 579674 322632
rect 579632 321638 579660 322623
rect 579620 321632 579672 321638
rect 579620 321574 579672 321580
rect 579710 310856 579766 310865
rect 579710 310791 579766 310800
rect 579724 310554 579752 310791
rect 579712 310548 579764 310554
rect 579712 310490 579764 310496
rect 579618 275768 579674 275777
rect 579618 275703 579674 275712
rect 579632 274718 579660 275703
rect 579620 274712 579672 274718
rect 579620 274654 579672 274660
rect 580170 263936 580226 263945
rect 580170 263871 580226 263880
rect 580184 263634 580212 263871
rect 580172 263628 580224 263634
rect 580172 263570 580224 263576
rect 580170 228848 580226 228857
rect 580170 228783 580226 228792
rect 580184 227798 580212 228783
rect 580172 227792 580224 227798
rect 580172 227734 580224 227740
rect 579618 217016 579674 217025
rect 579618 216951 579674 216960
rect 579632 216714 579660 216951
rect 579620 216708 579672 216714
rect 579620 216650 579672 216656
rect 580276 200938 580304 557223
rect 580354 545592 580410 545601
rect 580354 545527 580410 545536
rect 580264 200932 580316 200938
rect 580264 200874 580316 200880
rect 580368 200802 580396 545527
rect 580446 510368 580502 510377
rect 580446 510303 580502 510312
rect 580460 200870 580488 510303
rect 580630 404832 580686 404841
rect 580630 404767 580686 404776
rect 580538 393000 580594 393009
rect 580538 392935 580594 392944
rect 580448 200864 580500 200870
rect 580448 200806 580500 200812
rect 580356 200796 580408 200802
rect 580356 200738 580408 200744
rect 527178 200696 527234 200705
rect 527178 200631 527234 200640
rect 580264 199844 580316 199850
rect 580264 199786 580316 199792
rect 580276 181937 580304 199786
rect 580262 181928 580318 181937
rect 580262 181863 580318 181872
rect 580262 170096 580318 170105
rect 580262 170031 580318 170040
rect 580170 158400 580226 158409
rect 580170 158335 580226 158344
rect 580184 157418 580212 158335
rect 580172 157412 580224 157418
rect 580172 157354 580224 157360
rect 514024 144900 514076 144906
rect 514024 144842 514076 144848
rect 437020 136604 437072 136610
rect 437020 136546 437072 136552
rect 504456 136604 504508 136610
rect 504456 136546 504508 136552
rect 437032 136105 437060 136546
rect 437018 136096 437074 136105
rect 437018 136031 437074 136040
rect 437388 133884 437440 133890
rect 437388 133826 437440 133832
rect 437400 133657 437428 133826
rect 437386 133648 437442 133657
rect 437386 133583 437442 133592
rect 437388 132456 437440 132462
rect 437388 132398 437440 132404
rect 437400 132025 437428 132398
rect 437386 132016 437442 132025
rect 437386 131951 437442 131960
rect 437388 129736 437440 129742
rect 437388 129678 437440 129684
rect 437400 129577 437428 129678
rect 437386 129568 437442 129577
rect 437386 129503 437442 129512
rect 436834 127800 436890 127809
rect 436834 127735 436890 127744
rect 436926 124536 436982 124545
rect 436926 124471 436982 124480
rect 436834 122904 436890 122913
rect 436834 122839 436890 122848
rect 436284 121032 436336 121038
rect 436284 120974 436336 120980
rect 436742 120456 436798 120465
rect 436742 120391 436798 120400
rect 436192 35896 436244 35902
rect 436192 35838 436244 35844
rect 436756 17950 436784 120391
rect 436848 64870 436876 122839
rect 436940 111790 436968 124471
rect 580276 121106 580304 170031
rect 580552 137970 580580 392935
rect 580644 341698 580672 404767
rect 580722 369608 580778 369617
rect 580722 369543 580778 369552
rect 580632 341692 580684 341698
rect 580632 341634 580684 341640
rect 580736 341562 580764 369543
rect 580814 357912 580870 357921
rect 580814 357847 580870 357856
rect 580828 341630 580856 357847
rect 580816 341624 580868 341630
rect 580816 341566 580868 341572
rect 580724 341556 580776 341562
rect 580724 341498 580776 341504
rect 580630 299160 580686 299169
rect 580630 299095 580686 299104
rect 580540 137964 580592 137970
rect 580540 137906 580592 137912
rect 580354 134872 580410 134881
rect 580354 134807 580410 134816
rect 580368 121174 580396 134807
rect 580644 133890 580672 299095
rect 580722 252240 580778 252249
rect 580722 252175 580778 252184
rect 580632 133884 580684 133890
rect 580632 133826 580684 133832
rect 580736 132462 580764 252175
rect 580814 205320 580870 205329
rect 580814 205255 580870 205264
rect 580724 132456 580776 132462
rect 580724 132398 580776 132404
rect 580828 129742 580856 205255
rect 580816 129736 580868 129742
rect 580816 129678 580868 129684
rect 580538 123176 580594 123185
rect 580538 123111 580594 123120
rect 580552 121242 580580 123111
rect 580540 121236 580592 121242
rect 580540 121178 580592 121184
rect 580356 121168 580408 121174
rect 580356 121110 580408 121116
rect 580264 121100 580316 121106
rect 580264 121042 580316 121048
rect 480904 118652 480956 118658
rect 480904 118594 480956 118600
rect 443000 118584 443052 118590
rect 443000 118526 443052 118532
rect 442262 118008 442318 118017
rect 442262 117943 442318 117952
rect 436928 111784 436980 111790
rect 436928 111726 436980 111732
rect 436836 64864 436888 64870
rect 436836 64806 436888 64812
rect 436744 17944 436796 17950
rect 436744 17886 436796 17892
rect 441804 8696 441856 8702
rect 441804 8638 441856 8644
rect 438216 8560 438268 8566
rect 438216 8502 438268 8508
rect 434628 8492 434680 8498
rect 434628 8434 434680 8440
rect 433522 4856 433578 4865
rect 433248 4820 433300 4826
rect 433522 4791 433578 4800
rect 433248 4762 433300 4768
rect 432328 3460 432380 3466
rect 432328 3402 432380 3408
rect 431222 3360 431278 3369
rect 431222 3295 431278 3304
rect 432340 480 432368 3402
rect 433536 480 433564 4791
rect 434640 480 434668 8434
rect 435824 7200 435876 7206
rect 435824 7142 435876 7148
rect 435836 480 435864 7142
rect 437020 7132 437072 7138
rect 437020 7074 437072 7080
rect 437032 480 437060 7074
rect 438228 480 438256 8502
rect 440608 7268 440660 7274
rect 440608 7210 440660 7216
rect 439412 3528 439464 3534
rect 439412 3470 439464 3476
rect 439424 480 439452 3470
rect 440620 480 440648 7210
rect 441816 480 441844 8638
rect 442276 7970 442304 117943
rect 442184 7942 442304 7970
rect 442184 3466 442212 7942
rect 442172 3460 442224 3466
rect 442172 3402 442224 3408
rect 443012 480 443040 118526
rect 475384 118516 475436 118522
rect 475384 118458 475436 118464
rect 449900 118380 449952 118386
rect 449900 118322 449952 118328
rect 448980 8764 449032 8770
rect 448980 8706 449032 8712
rect 445392 8628 445444 8634
rect 445392 8570 445444 8576
rect 444196 7336 444248 7342
rect 444196 7278 444248 7284
rect 444208 480 444236 7278
rect 445404 480 445432 8570
rect 447784 7404 447836 7410
rect 447784 7346 447836 7352
rect 446588 2848 446640 2854
rect 446588 2790 446640 2796
rect 446600 480 446628 2790
rect 447796 480 447824 7346
rect 448992 480 449020 8706
rect 449912 626 449940 118322
rect 469864 118312 469916 118318
rect 469864 118254 469916 118260
rect 456800 118176 456852 118182
rect 456800 118118 456852 118124
rect 454868 9648 454920 9654
rect 454868 9590 454920 9596
rect 452476 8832 452528 8838
rect 452476 8774 452528 8780
rect 451280 7472 451332 7478
rect 451280 7414 451332 7420
rect 449912 598 450216 626
rect 450188 480 450216 598
rect 451292 480 451320 7414
rect 452488 480 452516 8774
rect 453672 3052 453724 3058
rect 453672 2994 453724 3000
rect 453684 480 453712 2994
rect 454880 480 454908 9590
rect 456064 8900 456116 8906
rect 456064 8842 456116 8848
rect 456076 480 456104 8842
rect 456812 610 456840 118118
rect 463700 118108 463752 118114
rect 463700 118050 463752 118056
rect 463712 12442 463740 118050
rect 463700 12436 463752 12442
rect 463700 12378 463752 12384
rect 464344 12436 464396 12442
rect 464344 12378 464396 12384
rect 464356 12322 464384 12378
rect 464356 12294 464476 12322
rect 459652 10736 459704 10742
rect 459652 10678 459704 10684
rect 458456 9580 458508 9586
rect 458456 9522 458508 9528
rect 456800 604 456852 610
rect 456800 546 456852 552
rect 457260 604 457312 610
rect 457260 546 457312 552
rect 457272 480 457300 546
rect 458468 480 458496 9522
rect 459664 480 459692 10678
rect 463240 10668 463292 10674
rect 463240 10610 463292 10616
rect 462044 9512 462096 9518
rect 462044 9454 462096 9460
rect 460848 3120 460900 3126
rect 460848 3062 460900 3068
rect 460860 480 460888 3062
rect 462056 480 462084 9454
rect 463252 480 463280 10610
rect 464448 480 464476 12294
rect 466828 10600 466880 10606
rect 466828 10542 466880 10548
rect 465632 5636 465684 5642
rect 465632 5578 465684 5584
rect 465644 480 465672 5578
rect 466840 480 466868 10542
rect 469128 5568 469180 5574
rect 469128 5510 469180 5516
rect 467932 3188 467984 3194
rect 467932 3130 467984 3136
rect 467944 480 467972 3130
rect 469140 480 469168 5510
rect 469876 3126 469904 118254
rect 474004 118244 474056 118250
rect 474004 118186 474056 118192
rect 470600 118040 470652 118046
rect 470600 117982 470652 117988
rect 470324 10532 470376 10538
rect 470324 10474 470376 10480
rect 469864 3120 469916 3126
rect 469864 3062 469916 3068
rect 470336 480 470364 10474
rect 470612 610 470640 117982
rect 473360 10464 473412 10470
rect 473360 10406 473412 10412
rect 472716 5704 472768 5710
rect 472716 5646 472768 5652
rect 470600 604 470652 610
rect 470600 546 470652 552
rect 471520 604 471572 610
rect 471520 546 471572 552
rect 471532 480 471560 546
rect 472728 480 472756 5646
rect 473372 610 473400 10406
rect 474016 3194 474044 118186
rect 475108 3256 475160 3262
rect 475108 3198 475160 3204
rect 474004 3188 474056 3194
rect 474004 3130 474056 3136
rect 473360 604 473412 610
rect 473360 546 473412 552
rect 473912 604 473964 610
rect 473912 546 473964 552
rect 473924 480 473952 546
rect 475120 480 475148 3198
rect 475396 3058 475424 118458
rect 478144 118448 478196 118454
rect 478144 118390 478196 118396
rect 477500 117972 477552 117978
rect 477500 117914 477552 117920
rect 477512 7546 477540 117914
rect 477592 10396 477644 10402
rect 477592 10338 477644 10344
rect 477500 7540 477552 7546
rect 477500 7482 477552 7488
rect 477604 7426 477632 10338
rect 477512 7398 477632 7426
rect 476304 5840 476356 5846
rect 476304 5782 476356 5788
rect 475384 3052 475436 3058
rect 475384 2994 475436 3000
rect 476316 480 476344 5782
rect 477512 480 477540 7398
rect 478156 3194 478184 118390
rect 478696 7540 478748 7546
rect 478696 7482 478748 7488
rect 478144 3188 478196 3194
rect 478144 3130 478196 3136
rect 478708 480 478736 7482
rect 479892 5772 479944 5778
rect 479892 5714 479944 5720
rect 479904 480 479932 5714
rect 480916 2922 480944 118594
rect 511264 117904 511316 117910
rect 511264 117846 511316 117852
rect 500224 117836 500276 117842
rect 500224 117778 500276 117784
rect 482284 117700 482336 117706
rect 482284 117642 482336 117648
rect 482296 11370 482324 117642
rect 486424 117632 486476 117638
rect 486424 117574 486476 117580
rect 482296 11342 482416 11370
rect 481088 10328 481140 10334
rect 481088 10270 481140 10276
rect 480904 2916 480956 2922
rect 480904 2858 480956 2864
rect 481100 480 481128 10270
rect 482284 3324 482336 3330
rect 482284 3266 482336 3272
rect 482296 480 482324 3266
rect 482388 2990 482416 11342
rect 483480 7472 483532 7478
rect 483480 7414 483532 7420
rect 482376 2984 482428 2990
rect 482376 2926 482428 2932
rect 483492 480 483520 7414
rect 484584 5976 484636 5982
rect 484584 5918 484636 5924
rect 484596 480 484624 5918
rect 486436 3330 486464 117574
rect 493324 117428 493376 117434
rect 493324 117370 493376 117376
rect 489184 117360 489236 117366
rect 489184 117302 489236 117308
rect 486976 8288 487028 8294
rect 486976 8230 487028 8236
rect 486424 3324 486476 3330
rect 486424 3266 486476 3272
rect 485780 2916 485832 2922
rect 485780 2858 485832 2864
rect 485792 480 485820 2858
rect 486988 480 487016 8230
rect 488172 5908 488224 5914
rect 488172 5850 488224 5856
rect 488184 480 488212 5850
rect 489196 3058 489224 117302
rect 490564 8220 490616 8226
rect 490564 8162 490616 8168
rect 489368 3120 489420 3126
rect 489368 3062 489420 3068
rect 489184 3052 489236 3058
rect 489184 2994 489236 3000
rect 489380 480 489408 3062
rect 490576 480 490604 8162
rect 491760 6044 491812 6050
rect 491760 5986 491812 5992
rect 491772 480 491800 5986
rect 493336 3398 493364 117370
rect 496084 116952 496136 116958
rect 496084 116894 496136 116900
rect 494152 8152 494204 8158
rect 494152 8094 494204 8100
rect 492956 3392 493008 3398
rect 492956 3334 493008 3340
rect 493324 3392 493376 3398
rect 493324 3334 493376 3340
rect 492968 480 492996 3334
rect 494164 480 494192 8094
rect 495348 6112 495400 6118
rect 495348 6054 495400 6060
rect 495360 480 495388 6054
rect 496096 3398 496124 116894
rect 497740 8084 497792 8090
rect 497740 8026 497792 8032
rect 496084 3392 496136 3398
rect 496084 3334 496136 3340
rect 496544 3256 496596 3262
rect 496544 3198 496596 3204
rect 496556 480 496584 3198
rect 497752 480 497780 8026
rect 498936 6860 498988 6866
rect 498936 6802 498988 6808
rect 498948 480 498976 6802
rect 500132 4140 500184 4146
rect 500132 4082 500184 4088
rect 500144 480 500172 4082
rect 500236 3330 500264 117778
rect 507124 117768 507176 117774
rect 507124 117710 507176 117716
rect 502984 117564 503036 117570
rect 502984 117506 503036 117512
rect 501236 8016 501288 8022
rect 501236 7958 501288 7964
rect 500224 3324 500276 3330
rect 500224 3266 500276 3272
rect 501248 480 501276 7958
rect 502432 6792 502484 6798
rect 502432 6734 502484 6740
rect 502444 480 502472 6734
rect 502996 4146 503024 117506
rect 504824 7948 504876 7954
rect 504824 7890 504876 7896
rect 502984 4140 503036 4146
rect 502984 4082 503036 4088
rect 503628 3188 503680 3194
rect 503628 3130 503680 3136
rect 503640 480 503668 3130
rect 504836 480 504864 7890
rect 506020 6724 506072 6730
rect 506020 6666 506072 6672
rect 506032 480 506060 6666
rect 507136 4146 507164 117710
rect 508412 7880 508464 7886
rect 508412 7822 508464 7828
rect 507124 4140 507176 4146
rect 507124 4082 507176 4088
rect 507216 4072 507268 4078
rect 507216 4014 507268 4020
rect 507228 480 507256 4014
rect 508424 480 508452 7822
rect 509608 6656 509660 6662
rect 509608 6598 509660 6604
rect 509620 480 509648 6598
rect 511276 3398 511304 117846
rect 579804 111784 579856 111790
rect 579804 111726 579856 111732
rect 579816 111489 579844 111726
rect 579802 111480 579858 111489
rect 579802 111415 579858 111424
rect 580172 88324 580224 88330
rect 580172 88266 580224 88272
rect 580184 87961 580212 88266
rect 580170 87952 580226 87961
rect 580170 87887 580226 87896
rect 580172 77240 580224 77246
rect 580172 77182 580224 77188
rect 580184 76265 580212 77182
rect 580170 76256 580226 76265
rect 580170 76191 580226 76200
rect 579804 64864 579856 64870
rect 579804 64806 579856 64812
rect 579816 64569 579844 64806
rect 579802 64560 579858 64569
rect 579802 64495 579858 64504
rect 580172 41404 580224 41410
rect 580172 41346 580224 41352
rect 580184 41041 580212 41346
rect 580170 41032 580226 41041
rect 580170 40967 580226 40976
rect 580172 30320 580224 30326
rect 580172 30262 580224 30268
rect 580184 29345 580212 30262
rect 580170 29336 580226 29345
rect 580170 29271 580226 29280
rect 579804 17944 579856 17950
rect 579804 17886 579856 17892
rect 579816 17649 579844 17886
rect 579802 17640 579858 17649
rect 579802 17575 579858 17584
rect 552388 9444 552440 9450
rect 552388 9386 552440 9392
rect 541716 7812 541768 7818
rect 541716 7754 541768 7760
rect 513196 6588 513248 6594
rect 513196 6530 513248 6536
rect 512000 4208 512052 4214
rect 512000 4150 512052 4156
rect 510804 3392 510856 3398
rect 510804 3334 510856 3340
rect 511264 3392 511316 3398
rect 511264 3334 511316 3340
rect 510816 480 510844 3334
rect 512012 480 512040 4150
rect 513208 480 513236 6530
rect 516784 6520 516836 6526
rect 516784 6462 516836 6468
rect 515588 4276 515640 4282
rect 515588 4218 515640 4224
rect 514392 4004 514444 4010
rect 514392 3946 514444 3952
rect 514404 480 514432 3946
rect 515600 480 515628 4218
rect 516796 480 516824 6462
rect 520280 6452 520332 6458
rect 520280 6394 520332 6400
rect 519084 4412 519136 4418
rect 519084 4354 519136 4360
rect 517888 2848 517940 2854
rect 517888 2790 517940 2796
rect 517900 480 517928 2790
rect 519096 480 519124 4354
rect 520292 480 520320 6394
rect 523868 6384 523920 6390
rect 523868 6326 523920 6332
rect 522672 4344 522724 4350
rect 522672 4286 522724 4292
rect 521476 3936 521528 3942
rect 521476 3878 521528 3884
rect 521488 480 521516 3878
rect 522684 480 522712 4286
rect 523880 480 523908 6326
rect 531044 6316 531096 6322
rect 531044 6258 531096 6264
rect 527456 6248 527508 6254
rect 527456 6190 527508 6196
rect 526260 4480 526312 4486
rect 526260 4422 526312 4428
rect 525064 2916 525116 2922
rect 525064 2858 525116 2864
rect 525076 480 525104 2858
rect 526272 480 526300 4422
rect 527468 480 527496 6190
rect 529848 4548 529900 4554
rect 529848 4490 529900 4496
rect 528652 3868 528704 3874
rect 528652 3810 528704 3816
rect 528664 480 528692 3810
rect 529860 480 529888 4490
rect 531056 480 531084 6258
rect 538126 6216 538182 6225
rect 534540 6180 534592 6186
rect 538126 6151 538182 6160
rect 534540 6122 534592 6128
rect 533436 4616 533488 4622
rect 533436 4558 533488 4564
rect 532240 3052 532292 3058
rect 532240 2994 532292 3000
rect 532252 480 532280 2994
rect 533448 480 533476 4558
rect 534552 480 534580 6122
rect 536932 4684 536984 4690
rect 536932 4626 536984 4632
rect 535736 3800 535788 3806
rect 535736 3742 535788 3748
rect 535748 480 535776 3742
rect 536944 480 536972 4626
rect 538140 480 538168 6151
rect 540520 4752 540572 4758
rect 540520 4694 540572 4700
rect 539324 3120 539376 3126
rect 539324 3062 539376 3068
rect 539336 480 539364 3062
rect 540532 480 540560 4694
rect 541728 480 541756 7754
rect 545304 7744 545356 7750
rect 545304 7686 545356 7692
rect 544108 5500 544160 5506
rect 544108 5442 544160 5448
rect 542912 3732 542964 3738
rect 542912 3674 542964 3680
rect 542924 480 542952 3674
rect 544120 480 544148 5442
rect 545316 480 545344 7686
rect 548892 7676 548944 7682
rect 548892 7618 548944 7624
rect 547696 5432 547748 5438
rect 547696 5374 547748 5380
rect 546500 3256 546552 3262
rect 546500 3198 546552 3204
rect 546512 480 546540 3198
rect 547708 480 547736 5374
rect 548904 480 548932 7618
rect 551192 5364 551244 5370
rect 551192 5306 551244 5312
rect 550088 3188 550140 3194
rect 550088 3130 550140 3136
rect 550100 480 550128 3130
rect 551204 480 551232 5306
rect 552400 480 552428 9386
rect 555976 9376 556028 9382
rect 555976 9318 556028 9324
rect 554780 5296 554832 5302
rect 554780 5238 554832 5244
rect 553584 3664 553636 3670
rect 553584 3606 553636 3612
rect 553596 480 553624 3606
rect 554792 480 554820 5238
rect 555988 480 556016 9318
rect 559564 9308 559616 9314
rect 559564 9250 559616 9256
rect 558368 5228 558420 5234
rect 558368 5170 558420 5176
rect 557172 3324 557224 3330
rect 557172 3266 557224 3272
rect 557184 480 557212 3266
rect 558380 480 558408 5170
rect 559576 480 559604 9250
rect 563152 9240 563204 9246
rect 563152 9182 563204 9188
rect 561956 5160 562008 5166
rect 561956 5102 562008 5108
rect 560760 3596 560812 3602
rect 560760 3538 560812 3544
rect 560772 480 560800 3538
rect 561968 480 561996 5102
rect 563164 480 563192 9182
rect 566740 9172 566792 9178
rect 566740 9114 566792 9120
rect 565544 5092 565596 5098
rect 565544 5034 565596 5040
rect 564348 3392 564400 3398
rect 564348 3334 564400 3340
rect 564360 480 564388 3334
rect 565556 480 565584 5034
rect 566752 480 566780 9114
rect 570236 9104 570288 9110
rect 570236 9046 570288 9052
rect 569040 5024 569092 5030
rect 569040 4966 569092 4972
rect 567844 3528 567896 3534
rect 567844 3470 567896 3476
rect 567856 480 567884 3470
rect 569052 480 569080 4966
rect 570248 480 570276 9046
rect 577412 9036 577464 9042
rect 577412 8978 577464 8984
rect 573824 7608 573876 7614
rect 573824 7550 573876 7556
rect 572628 4956 572680 4962
rect 572628 4898 572680 4904
rect 571432 4140 571484 4146
rect 571432 4082 571484 4088
rect 571444 480 571472 4082
rect 572640 480 572668 4898
rect 573836 480 573864 7550
rect 576216 4888 576268 4894
rect 576216 4830 576268 4836
rect 575018 3360 575074 3369
rect 575018 3295 575074 3304
rect 575032 480 575060 3295
rect 576228 480 576256 4830
rect 577424 480 577452 8978
rect 581000 8968 581052 8974
rect 581000 8910 581052 8916
rect 579804 4820 579856 4826
rect 579804 4762 579856 4768
rect 578608 4072 578660 4078
rect 578608 4014 578660 4020
rect 578620 480 578648 4014
rect 579816 480 579844 4762
rect 581012 480 581040 8910
rect 582196 3460 582248 3466
rect 582196 3402 582248 3408
rect 582208 480 582236 3402
rect 542 -960 654 480
rect 1646 -960 1758 480
rect 2842 -960 2954 480
rect 4038 -960 4150 480
rect 5234 -960 5346 480
rect 6430 -960 6542 480
rect 7626 -960 7738 480
rect 8822 -960 8934 480
rect 10018 -960 10130 480
rect 11214 -960 11326 480
rect 12410 -960 12522 480
rect 13606 -960 13718 480
rect 14802 -960 14914 480
rect 15998 -960 16110 480
rect 17194 -960 17306 480
rect 18298 -960 18410 480
rect 19494 -960 19606 480
rect 20690 -960 20802 480
rect 21886 -960 21998 480
rect 23082 -960 23194 480
rect 24278 -960 24390 480
rect 25474 -960 25586 480
rect 26670 -960 26782 480
rect 27866 -960 27978 480
rect 29062 -960 29174 480
rect 30258 -960 30370 480
rect 31454 -960 31566 480
rect 32650 -960 32762 480
rect 33846 -960 33958 480
rect 34950 -960 35062 480
rect 36146 -960 36258 480
rect 37342 -960 37454 480
rect 38538 -960 38650 480
rect 39734 -960 39846 480
rect 40930 -960 41042 480
rect 42126 -960 42238 480
rect 43322 -960 43434 480
rect 44518 -960 44630 480
rect 45714 -960 45826 480
rect 46910 -960 47022 480
rect 48106 -960 48218 480
rect 49302 -960 49414 480
rect 50498 -960 50610 480
rect 51602 -960 51714 480
rect 52798 -960 52910 480
rect 53994 -960 54106 480
rect 55190 -960 55302 480
rect 56386 -960 56498 480
rect 57582 -960 57694 480
rect 58778 -960 58890 480
rect 59974 -960 60086 480
rect 61170 -960 61282 480
rect 62366 -960 62478 480
rect 63562 -960 63674 480
rect 64758 -960 64870 480
rect 65954 -960 66066 480
rect 67150 -960 67262 480
rect 68254 -960 68366 480
rect 69450 -960 69562 480
rect 70646 -960 70758 480
rect 71842 -960 71954 480
rect 73038 -960 73150 480
rect 74234 -960 74346 480
rect 75430 -960 75542 480
rect 76626 -960 76738 480
rect 77822 -960 77934 480
rect 79018 -960 79130 480
rect 80214 -960 80326 480
rect 81410 -960 81522 480
rect 82606 -960 82718 480
rect 83802 -960 83914 480
rect 84906 -960 85018 480
rect 86102 -960 86214 480
rect 87298 -960 87410 480
rect 88494 -960 88606 480
rect 89690 -960 89802 480
rect 90886 -960 90998 480
rect 92082 -960 92194 480
rect 93278 -960 93390 480
rect 94474 -960 94586 480
rect 95670 -960 95782 480
rect 96866 -960 96978 480
rect 98062 -960 98174 480
rect 99258 -960 99370 480
rect 100454 -960 100566 480
rect 101558 -960 101670 480
rect 102754 -960 102866 480
rect 103950 -960 104062 480
rect 105146 -960 105258 480
rect 106342 -960 106454 480
rect 107538 -960 107650 480
rect 108734 -960 108846 480
rect 109930 -960 110042 480
rect 111126 -960 111238 480
rect 112322 -960 112434 480
rect 113518 -960 113630 480
rect 114714 -960 114826 480
rect 115910 -960 116022 480
rect 117106 -960 117218 480
rect 118210 -960 118322 480
rect 119406 -960 119518 480
rect 120602 -960 120714 480
rect 121798 -960 121910 480
rect 122994 -960 123106 480
rect 124190 -960 124302 480
rect 125386 -960 125498 480
rect 126582 -960 126694 480
rect 127778 -960 127890 480
rect 128974 -960 129086 480
rect 130170 -960 130282 480
rect 131366 -960 131478 480
rect 132562 -960 132674 480
rect 133758 -960 133870 480
rect 134862 -960 134974 480
rect 136058 -960 136170 480
rect 137254 -960 137366 480
rect 138450 -960 138562 480
rect 139646 -960 139758 480
rect 140842 -960 140954 480
rect 142038 -960 142150 480
rect 143234 -960 143346 480
rect 144430 -960 144542 480
rect 145626 -960 145738 480
rect 146822 -960 146934 480
rect 148018 -960 148130 480
rect 149214 -960 149326 480
rect 150410 -960 150522 480
rect 151514 -960 151626 480
rect 152710 -960 152822 480
rect 153906 -960 154018 480
rect 155102 -960 155214 480
rect 156298 -960 156410 480
rect 157494 -960 157606 480
rect 158690 -960 158802 480
rect 159886 -960 159998 480
rect 161082 -960 161194 480
rect 162278 -960 162390 480
rect 163474 -960 163586 480
rect 164670 -960 164782 480
rect 165866 -960 165978 480
rect 167062 -960 167174 480
rect 168166 -960 168278 480
rect 169362 -960 169474 480
rect 170558 -960 170670 480
rect 171754 -960 171866 480
rect 172950 -960 173062 480
rect 174146 -960 174258 480
rect 175342 -960 175454 480
rect 176538 -960 176650 480
rect 177734 -960 177846 480
rect 178930 -960 179042 480
rect 180126 -960 180238 480
rect 181322 -960 181434 480
rect 182518 -960 182630 480
rect 183714 -960 183826 480
rect 184818 -960 184930 480
rect 186014 -960 186126 480
rect 187210 -960 187322 480
rect 188406 -960 188518 480
rect 189602 -960 189714 480
rect 190798 -960 190910 480
rect 191994 -960 192106 480
rect 193190 -960 193302 480
rect 194386 -960 194498 480
rect 195582 -960 195694 480
rect 196778 -960 196890 480
rect 197974 -960 198086 480
rect 199170 -960 199282 480
rect 200366 -960 200478 480
rect 201470 -960 201582 480
rect 202666 -960 202778 480
rect 203862 -960 203974 480
rect 205058 -960 205170 480
rect 206254 -960 206366 480
rect 207450 -960 207562 480
rect 208646 -960 208758 480
rect 209842 -960 209954 480
rect 211038 -960 211150 480
rect 212234 -960 212346 480
rect 213430 -960 213542 480
rect 214626 -960 214738 480
rect 215822 -960 215934 480
rect 217018 -960 217130 480
rect 218122 -960 218234 480
rect 219318 -960 219430 480
rect 220514 -960 220626 480
rect 221710 -960 221822 480
rect 222906 -960 223018 480
rect 224102 -960 224214 480
rect 225298 -960 225410 480
rect 226494 -960 226606 480
rect 227690 -960 227802 480
rect 228886 -960 228998 480
rect 230082 -960 230194 480
rect 231278 -960 231390 480
rect 232474 -960 232586 480
rect 233670 -960 233782 480
rect 234774 -960 234886 480
rect 235970 -960 236082 480
rect 237166 -960 237278 480
rect 238362 -960 238474 480
rect 239558 -960 239670 480
rect 240754 -960 240866 480
rect 241950 -960 242062 480
rect 243146 -960 243258 480
rect 244342 -960 244454 480
rect 245538 -960 245650 480
rect 246734 -960 246846 480
rect 247930 -960 248042 480
rect 249126 -960 249238 480
rect 250322 -960 250434 480
rect 251426 -960 251538 480
rect 252622 -960 252734 480
rect 253818 -960 253930 480
rect 255014 -960 255126 480
rect 256210 -960 256322 480
rect 257406 -960 257518 480
rect 258602 -960 258714 480
rect 259798 -960 259910 480
rect 260994 -960 261106 480
rect 262190 -960 262302 480
rect 263386 -960 263498 480
rect 264582 -960 264694 480
rect 265778 -960 265890 480
rect 266974 -960 267086 480
rect 268078 -960 268190 480
rect 269274 -960 269386 480
rect 270470 -960 270582 480
rect 271666 -960 271778 480
rect 272862 -960 272974 480
rect 274058 -960 274170 480
rect 275254 -960 275366 480
rect 276450 -960 276562 480
rect 277646 -960 277758 480
rect 278842 -960 278954 480
rect 280038 -960 280150 480
rect 281234 -960 281346 480
rect 282430 -960 282542 480
rect 283626 -960 283738 480
rect 284730 -960 284842 480
rect 285926 -960 286038 480
rect 287122 -960 287234 480
rect 288318 -960 288430 480
rect 289514 -960 289626 480
rect 290710 -960 290822 480
rect 291906 -960 292018 480
rect 293102 -960 293214 480
rect 294298 -960 294410 480
rect 295494 -960 295606 480
rect 296690 -960 296802 480
rect 297886 -960 297998 480
rect 299082 -960 299194 480
rect 300278 -960 300390 480
rect 301382 -960 301494 480
rect 302578 -960 302690 480
rect 303774 -960 303886 480
rect 304970 -960 305082 480
rect 306166 -960 306278 480
rect 307362 -960 307474 480
rect 308558 -960 308670 480
rect 309754 -960 309866 480
rect 310950 -960 311062 480
rect 312146 -960 312258 480
rect 313342 -960 313454 480
rect 314538 -960 314650 480
rect 315734 -960 315846 480
rect 316930 -960 317042 480
rect 318034 -960 318146 480
rect 319230 -960 319342 480
rect 320426 -960 320538 480
rect 321622 -960 321734 480
rect 322818 -960 322930 480
rect 324014 -960 324126 480
rect 325210 -960 325322 480
rect 326406 -960 326518 480
rect 327602 -960 327714 480
rect 328798 -960 328910 480
rect 329994 -960 330106 480
rect 331190 -960 331302 480
rect 332386 -960 332498 480
rect 333582 -960 333694 480
rect 334686 -960 334798 480
rect 335882 -960 335994 480
rect 337078 -960 337190 480
rect 338274 -960 338386 480
rect 339470 -960 339582 480
rect 340666 -960 340778 480
rect 341862 -960 341974 480
rect 343058 -960 343170 480
rect 344254 -960 344366 480
rect 345450 -960 345562 480
rect 346646 -960 346758 480
rect 347842 -960 347954 480
rect 349038 -960 349150 480
rect 350234 -960 350346 480
rect 351338 -960 351450 480
rect 352534 -960 352646 480
rect 353730 -960 353842 480
rect 354926 -960 355038 480
rect 356122 -960 356234 480
rect 357318 -960 357430 480
rect 358514 -960 358626 480
rect 359710 -960 359822 480
rect 360906 -960 361018 480
rect 362102 -960 362214 480
rect 363298 -960 363410 480
rect 364494 -960 364606 480
rect 365690 -960 365802 480
rect 366886 -960 366998 480
rect 367990 -960 368102 480
rect 369186 -960 369298 480
rect 370382 -960 370494 480
rect 371578 -960 371690 480
rect 372774 -960 372886 480
rect 373970 -960 374082 480
rect 375166 -960 375278 480
rect 376362 -960 376474 480
rect 377558 -960 377670 480
rect 378754 -960 378866 480
rect 379950 -960 380062 480
rect 381146 -960 381258 480
rect 382342 -960 382454 480
rect 383538 -960 383650 480
rect 384642 -960 384754 480
rect 385838 -960 385950 480
rect 387034 -960 387146 480
rect 388230 -960 388342 480
rect 389426 -960 389538 480
rect 390622 -960 390734 480
rect 391818 -960 391930 480
rect 393014 -960 393126 480
rect 394210 -960 394322 480
rect 395406 -960 395518 480
rect 396602 -960 396714 480
rect 397798 -960 397910 480
rect 398994 -960 399106 480
rect 400190 -960 400302 480
rect 401294 -960 401406 480
rect 402490 -960 402602 480
rect 403686 -960 403798 480
rect 404882 -960 404994 480
rect 406078 -960 406190 480
rect 407274 -960 407386 480
rect 408470 -960 408582 480
rect 409666 -960 409778 480
rect 410862 -960 410974 480
rect 412058 -960 412170 480
rect 413254 -960 413366 480
rect 414450 -960 414562 480
rect 415646 -960 415758 480
rect 416842 -960 416954 480
rect 417946 -960 418058 480
rect 419142 -960 419254 480
rect 420338 -960 420450 480
rect 421534 -960 421646 480
rect 422730 -960 422842 480
rect 423926 -960 424038 480
rect 425122 -960 425234 480
rect 426318 -960 426430 480
rect 427514 -960 427626 480
rect 428710 -960 428822 480
rect 429906 -960 430018 480
rect 431102 -960 431214 480
rect 432298 -960 432410 480
rect 433494 -960 433606 480
rect 434598 -960 434710 480
rect 435794 -960 435906 480
rect 436990 -960 437102 480
rect 438186 -960 438298 480
rect 439382 -960 439494 480
rect 440578 -960 440690 480
rect 441774 -960 441886 480
rect 442970 -960 443082 480
rect 444166 -960 444278 480
rect 445362 -960 445474 480
rect 446558 -960 446670 480
rect 447754 -960 447866 480
rect 448950 -960 449062 480
rect 450146 -960 450258 480
rect 451250 -960 451362 480
rect 452446 -960 452558 480
rect 453642 -960 453754 480
rect 454838 -960 454950 480
rect 456034 -960 456146 480
rect 457230 -960 457342 480
rect 458426 -960 458538 480
rect 459622 -960 459734 480
rect 460818 -960 460930 480
rect 462014 -960 462126 480
rect 463210 -960 463322 480
rect 464406 -960 464518 480
rect 465602 -960 465714 480
rect 466798 -960 466910 480
rect 467902 -960 468014 480
rect 469098 -960 469210 480
rect 470294 -960 470406 480
rect 471490 -960 471602 480
rect 472686 -960 472798 480
rect 473882 -960 473994 480
rect 475078 -960 475190 480
rect 476274 -960 476386 480
rect 477470 -960 477582 480
rect 478666 -960 478778 480
rect 479862 -960 479974 480
rect 481058 -960 481170 480
rect 482254 -960 482366 480
rect 483450 -960 483562 480
rect 484554 -960 484666 480
rect 485750 -960 485862 480
rect 486946 -960 487058 480
rect 488142 -960 488254 480
rect 489338 -960 489450 480
rect 490534 -960 490646 480
rect 491730 -960 491842 480
rect 492926 -960 493038 480
rect 494122 -960 494234 480
rect 495318 -960 495430 480
rect 496514 -960 496626 480
rect 497710 -960 497822 480
rect 498906 -960 499018 480
rect 500102 -960 500214 480
rect 501206 -960 501318 480
rect 502402 -960 502514 480
rect 503598 -960 503710 480
rect 504794 -960 504906 480
rect 505990 -960 506102 480
rect 507186 -960 507298 480
rect 508382 -960 508494 480
rect 509578 -960 509690 480
rect 510774 -960 510886 480
rect 511970 -960 512082 480
rect 513166 -960 513278 480
rect 514362 -960 514474 480
rect 515558 -960 515670 480
rect 516754 -960 516866 480
rect 517858 -960 517970 480
rect 519054 -960 519166 480
rect 520250 -960 520362 480
rect 521446 -960 521558 480
rect 522642 -960 522754 480
rect 523838 -960 523950 480
rect 525034 -960 525146 480
rect 526230 -960 526342 480
rect 527426 -960 527538 480
rect 528622 -960 528734 480
rect 529818 -960 529930 480
rect 531014 -960 531126 480
rect 532210 -960 532322 480
rect 533406 -960 533518 480
rect 534510 -960 534622 480
rect 535706 -960 535818 480
rect 536902 -960 537014 480
rect 538098 -960 538210 480
rect 539294 -960 539406 480
rect 540490 -960 540602 480
rect 541686 -960 541798 480
rect 542882 -960 542994 480
rect 544078 -960 544190 480
rect 545274 -960 545386 480
rect 546470 -960 546582 480
rect 547666 -960 547778 480
rect 548862 -960 548974 480
rect 550058 -960 550170 480
rect 551162 -960 551274 480
rect 552358 -960 552470 480
rect 553554 -960 553666 480
rect 554750 -960 554862 480
rect 555946 -960 556058 480
rect 557142 -960 557254 480
rect 558338 -960 558450 480
rect 559534 -960 559646 480
rect 560730 -960 560842 480
rect 561926 -960 562038 480
rect 563122 -960 563234 480
rect 564318 -960 564430 480
rect 565514 -960 565626 480
rect 566710 -960 566822 480
rect 567814 -960 567926 480
rect 569010 -960 569122 480
rect 570206 -960 570318 480
rect 571402 -960 571514 480
rect 572598 -960 572710 480
rect 573794 -960 573906 480
rect 574990 -960 575102 480
rect 576186 -960 576298 480
rect 577382 -960 577494 480
rect 578578 -960 578690 480
rect 579774 -960 579886 480
rect 580970 -960 581082 480
rect 582166 -960 582278 480
rect 583362 -960 583474 480
<< via2 >>
rect 3514 682216 3570 682272
rect 3422 667956 3478 667992
rect 3422 667936 3424 667956
rect 3424 667936 3476 667956
rect 3476 667936 3478 667956
rect 4802 653520 4858 653576
rect 3422 624824 3478 624880
rect 3422 610408 3478 610464
rect 4066 595992 4122 596048
rect 3422 567296 3478 567352
rect 3146 553016 3202 553072
rect 3330 495508 3386 495544
rect 3330 495488 3332 495508
rect 3332 495488 3384 495508
rect 3384 495488 3386 495508
rect 3054 452376 3110 452432
rect 2778 366152 2834 366208
rect 2962 337456 3018 337512
rect 3330 294344 3386 294400
rect 2778 265648 2834 265704
rect 3330 251252 3386 251288
rect 3330 251232 3332 251252
rect 3332 251232 3384 251252
rect 3384 251232 3386 251252
rect 3330 236952 3386 237008
rect 2962 222536 3018 222592
rect 2962 208120 3018 208176
rect 2870 179424 2926 179480
rect 3238 165008 3294 165064
rect 3514 538600 3570 538656
rect 3238 150728 3294 150784
rect 3330 136312 3386 136368
rect 3054 122032 3110 122088
rect 2778 93200 2834 93256
rect 3238 78920 3294 78976
rect 3330 64504 3386 64560
rect 3606 509904 3662 509960
rect 4066 481072 4122 481128
rect 3698 437960 3754 438016
rect 3606 193840 3662 193896
rect 4066 423700 4122 423736
rect 4066 423680 4068 423700
rect 4068 423680 4120 423700
rect 4120 423680 4122 423700
rect 3882 394984 3938 395040
rect 3790 380568 3846 380624
rect 3974 323040 4030 323096
rect 4066 308760 4122 308816
rect 4066 280064 4122 280120
rect 3514 107616 3570 107672
rect 69938 385192 69994 385248
rect 69846 377848 69902 377904
rect 70030 362888 70086 362944
rect 70030 355544 70086 355600
rect 70306 392536 70362 392592
rect 71594 392536 71650 392592
rect 70306 377848 70362 377904
rect 70214 370232 70270 370288
rect 70122 348200 70178 348256
rect 70030 341400 70086 341456
rect 3422 50088 3478 50144
rect 3422 35844 3424 35864
rect 3424 35844 3476 35864
rect 3476 35844 3478 35864
rect 3422 35808 3478 35844
rect 3146 21392 3202 21448
rect 3422 7112 3478 7168
rect 30286 4800 30342 4856
rect 71502 348200 71558 348256
rect 84106 545808 84162 545864
rect 84014 541456 84070 541512
rect 83922 528672 83978 528728
rect 82818 524864 82874 524920
rect 85302 537104 85358 537160
rect 85210 533024 85266 533080
rect 86406 549908 86462 549944
rect 86406 549888 86408 549908
rect 86408 549888 86460 549908
rect 86460 549888 86462 549908
rect 85394 525544 85450 525600
rect 115294 498072 115350 498128
rect 118054 546488 118110 546544
rect 117778 537376 117834 537432
rect 117778 533296 117834 533352
rect 117962 529624 118018 529680
rect 117318 521056 117374 521112
rect 118606 542428 118662 542464
rect 118606 542408 118608 542428
rect 118608 542408 118660 542428
rect 118660 542408 118662 542428
rect 124862 582528 124918 582584
rect 118606 525136 118662 525192
rect 125966 495488 126022 495544
rect 125874 492632 125930 492688
rect 125874 415384 125930 415440
rect 126150 415404 126206 415440
rect 126150 415384 126152 415404
rect 126152 415384 126204 415404
rect 126204 415384 126206 415404
rect 125690 395664 125746 395720
rect 75918 118532 75920 118552
rect 75920 118532 75972 118552
rect 75972 118532 75974 118552
rect 75918 118496 75974 118532
rect 85394 118496 85450 118552
rect 71594 117952 71650 118008
rect 76010 117952 76066 118008
rect 70214 117408 70270 117464
rect 73986 48456 74042 48512
rect 73618 48320 73674 48376
rect 73618 34448 73674 34504
rect 73802 34448 73858 34504
rect 103426 118496 103482 118552
rect 100666 117544 100722 117600
rect 100022 117272 100078 117328
rect 100666 117272 100722 117328
rect 102138 117272 102194 117328
rect 103426 117272 103482 117328
rect 110326 117816 110382 117872
rect 117226 118360 117282 118416
rect 126058 395664 126114 395720
rect 126426 417424 126482 417480
rect 126886 395664 126942 395720
rect 128174 144472 128230 144528
rect 125782 118224 125838 118280
rect 115938 117272 115994 117328
rect 117226 117272 117282 117328
rect 113546 6160 113602 6216
rect 129554 500112 129610 500168
rect 128634 481616 128690 481672
rect 128818 481616 128874 481672
rect 128542 463664 128598 463720
rect 128818 463664 128874 463720
rect 128542 444352 128598 444408
rect 128818 444352 128874 444408
rect 128542 425040 128598 425096
rect 128818 425040 128874 425096
rect 128634 388184 128690 388240
rect 129094 380568 129150 380624
rect 128910 376896 128966 376952
rect 128818 376760 128874 376816
rect 128450 373224 128506 373280
rect 128358 358264 128414 358320
rect 128818 343576 128874 343632
rect 129002 350956 129004 350976
rect 129004 350956 129056 350976
rect 129056 350956 129058 350976
rect 129002 350920 129058 350956
rect 128818 182164 128874 182200
rect 128818 182144 128820 182164
rect 128820 182144 128872 182164
rect 128872 182144 128874 182164
rect 129002 182144 129058 182200
rect 128910 153312 128966 153368
rect 128818 153176 128874 153232
rect 128910 135360 128966 135416
rect 128818 135224 128874 135280
rect 128818 118632 128874 118688
rect 127622 117680 127678 117736
rect 128266 117680 128322 117736
rect 129186 373224 129242 373280
rect 129370 365880 129426 365936
rect 129278 358264 129334 358320
rect 128726 86944 128782 87000
rect 129002 86944 129058 87000
rect 131026 582392 131082 582448
rect 130934 500248 130990 500304
rect 130842 196152 130898 196208
rect 130842 194676 130898 194712
rect 130842 194656 130844 194676
rect 130844 194656 130896 194676
rect 130896 194656 130898 194676
rect 130842 194384 130898 194440
rect 130842 193060 130844 193080
rect 130844 193060 130896 193080
rect 130896 193060 130898 193080
rect 130842 193024 130898 193060
rect 130750 192480 130806 192536
rect 130842 191392 130898 191448
rect 130842 190304 130898 190360
rect 130842 188964 130898 189000
rect 130842 188944 130844 188964
rect 130844 188944 130896 188964
rect 130896 188944 130898 188964
rect 130750 188264 130806 188320
rect 130842 187176 130898 187232
rect 131210 185544 131266 185600
rect 131210 184456 131266 184512
rect 131210 183524 131266 183560
rect 131210 183504 131212 183524
rect 131212 183504 131264 183524
rect 131264 183504 131266 183524
rect 131210 178200 131266 178256
rect 131394 198192 131450 198248
rect 131394 197104 131450 197160
rect 131302 164464 131358 164520
rect 131302 157120 131358 157176
rect 131118 156168 131174 156224
rect 131118 155080 131174 155136
rect 131118 153992 131174 154048
rect 131118 152904 131174 152960
rect 131118 150864 131174 150920
rect 131118 149776 131174 149832
rect 131118 148688 131174 148744
rect 131118 147736 131174 147792
rect 131302 151952 131358 152008
rect 131210 146648 131266 146704
rect 131118 145560 131174 145616
rect 131118 143520 131174 143576
rect 131302 139304 131358 139360
rect 131394 131960 131450 132016
rect 131762 199280 131818 199336
rect 131670 167728 131726 167784
rect 131670 158208 131726 158264
rect 131578 125568 131634 125624
rect 131486 124480 131542 124536
rect 131946 128696 132002 128752
rect 132222 170856 132278 170912
rect 132222 159296 132278 159352
rect 132130 130872 132186 130928
rect 132038 127744 132094 127800
rect 131854 126656 131910 126712
rect 132130 121352 132186 121408
rect 132498 179288 132554 179344
rect 132590 177112 132646 177168
rect 132406 171944 132462 172000
rect 132774 166640 132830 166696
rect 132682 165552 132738 165608
rect 132406 162424 132462 162480
rect 132314 138216 132370 138272
rect 132682 161336 132738 161392
rect 132406 120400 132462 120456
rect 133142 169768 133198 169824
rect 133050 168680 133106 168736
rect 133326 182416 133382 182472
rect 133418 181328 133474 181384
rect 133602 163512 133658 163568
rect 133602 160384 133658 160440
rect 133510 142432 133566 142488
rect 133234 129784 133290 129840
rect 133050 106392 133106 106448
rect 133510 106256 133566 106312
rect 133694 141344 133750 141400
rect 147586 697076 147588 697096
rect 147588 697076 147640 697096
rect 147640 697076 147642 697096
rect 147586 697040 147642 697076
rect 154486 697176 154542 697232
rect 173806 697176 173862 697232
rect 193126 697176 193182 697232
rect 212446 697176 212502 697232
rect 231766 697176 231822 697232
rect 251086 697176 251142 697232
rect 270406 697176 270462 697232
rect 289726 697176 289782 697232
rect 309046 697176 309102 697232
rect 328366 697176 328422 697232
rect 166906 697076 166908 697096
rect 166908 697076 166960 697096
rect 166960 697076 166962 697096
rect 166906 697040 166962 697076
rect 186226 697076 186228 697096
rect 186228 697076 186280 697096
rect 186280 697076 186282 697096
rect 186226 697040 186282 697076
rect 205546 697076 205548 697096
rect 205548 697076 205600 697096
rect 205600 697076 205602 697096
rect 205546 697040 205602 697076
rect 224866 697076 224868 697096
rect 224868 697076 224920 697096
rect 224920 697076 224922 697096
rect 224866 697040 224922 697076
rect 244186 697076 244188 697096
rect 244188 697076 244240 697096
rect 244240 697076 244242 697096
rect 244186 697040 244242 697076
rect 263506 697076 263508 697096
rect 263508 697076 263560 697096
rect 263560 697076 263562 697096
rect 263506 697040 263562 697076
rect 282826 697076 282828 697096
rect 282828 697076 282880 697096
rect 282880 697076 282882 697096
rect 282826 697040 282882 697076
rect 302146 697076 302148 697096
rect 302148 697076 302200 697096
rect 302200 697076 302202 697096
rect 302146 697040 302202 697076
rect 321466 697076 321468 697096
rect 321468 697076 321520 697096
rect 321520 697076 321522 697096
rect 321466 697040 321522 697076
rect 135258 686180 135314 686216
rect 135258 686160 135260 686180
rect 135260 686160 135312 686180
rect 135312 686160 135314 686180
rect 147770 686296 147826 686352
rect 147586 686024 147642 686080
rect 169022 686432 169078 686488
rect 154578 686316 154634 686352
rect 154578 686296 154580 686316
rect 154580 686296 154632 686316
rect 154632 686296 154634 686316
rect 159454 686160 159510 686216
rect 169022 686160 169078 686216
rect 142894 685888 142950 685944
rect 169022 650528 169078 650584
rect 135258 650276 135314 650312
rect 135258 650256 135260 650276
rect 135260 650256 135312 650276
rect 135312 650256 135314 650276
rect 147770 650392 147826 650448
rect 154578 650412 154634 650448
rect 154578 650392 154580 650412
rect 154580 650392 154632 650412
rect 154632 650392 154634 650412
rect 159454 650256 159510 650312
rect 169022 650256 169078 650312
rect 147586 650120 147642 650176
rect 142894 649984 142950 650040
rect 157062 639240 157118 639296
rect 157246 639240 157302 639296
rect 171046 639240 171102 639296
rect 171046 638832 171102 638888
rect 157062 603336 157118 603392
rect 157246 603336 157302 603392
rect 171046 603336 171102 603392
rect 171046 602928 171102 602984
rect 169022 592592 169078 592648
rect 135258 592340 135314 592376
rect 135258 592320 135260 592340
rect 135260 592320 135312 592340
rect 135312 592320 135314 592340
rect 147770 592456 147826 592512
rect 154578 592476 154634 592512
rect 154578 592456 154580 592476
rect 154580 592456 154632 592476
rect 154632 592456 154634 592476
rect 159454 592320 159510 592376
rect 169022 592320 169078 592376
rect 147586 592184 147642 592240
rect 142894 592048 142950 592104
rect 191102 582936 191158 582992
rect 133970 341400 134026 341456
rect 133878 180376 133934 180432
rect 134062 249736 134118 249792
rect 134246 249736 134302 249792
rect 153290 521600 153346 521656
rect 153474 521600 153530 521656
rect 153290 482976 153346 483032
rect 153474 482976 153530 483032
rect 153382 447208 153438 447264
rect 153382 444372 153438 444408
rect 153382 444352 153384 444372
rect 153384 444352 153436 444372
rect 153436 444352 153438 444372
rect 153474 425176 153530 425232
rect 153198 425040 153254 425096
rect 185582 341400 185638 341456
rect 197082 202816 197138 202872
rect 197174 202680 197230 202736
rect 211618 561720 211674 561776
rect 222198 556144 222254 556200
rect 198646 534112 198702 534168
rect 198554 524592 198610 524648
rect 198002 378664 198058 378720
rect 197910 374312 197966 374368
rect 197818 370232 197874 370288
rect 197726 361800 197782 361856
rect 197542 357448 197598 357504
rect 197450 353368 197506 353424
rect 197358 349016 197414 349072
rect 197634 344936 197690 344992
rect 197266 202408 197322 202464
rect 196990 202136 197046 202192
rect 198462 399608 198518 399664
rect 198370 387096 198426 387152
rect 198738 529216 198794 529272
rect 198830 403688 198886 403744
rect 198922 395256 198978 395312
rect 199014 391176 199070 391232
rect 199106 382744 199162 382800
rect 199198 365880 199254 365936
rect 203338 410352 203394 410408
rect 222290 552064 222346 552120
rect 222566 546896 222622 546952
rect 222474 542544 222530 542600
rect 222382 538328 222438 538384
rect 222658 533296 222714 533352
rect 222750 528944 222806 529000
rect 222842 524456 222898 524512
rect 226154 410080 226210 410136
rect 231858 410216 231914 410272
rect 263138 409944 263194 410000
rect 209778 241440 209834 241496
rect 209962 241440 210018 241496
rect 209778 222128 209834 222184
rect 209962 222128 210018 222184
rect 211158 201592 211214 201648
rect 212538 201864 212594 201920
rect 213458 201728 213514 201784
rect 218058 202000 218114 202056
rect 220358 202816 220414 202872
rect 223854 202680 223910 202736
rect 225142 202544 225198 202600
rect 226338 202408 226394 202464
rect 232134 202272 232190 202328
rect 237194 338680 237250 338736
rect 233422 202136 233478 202192
rect 257710 317328 257766 317384
rect 257802 311752 257858 311808
rect 257066 202136 257122 202192
rect 262678 201592 262734 201648
rect 266174 202816 266230 202872
rect 266910 399608 266966 399664
rect 267186 357448 267242 357504
rect 267278 353368 267334 353424
rect 267646 349016 267702 349072
rect 267922 403688 267978 403744
rect 268014 395256 268070 395312
rect 268106 391176 268162 391232
rect 268198 386824 268254 386880
rect 268290 382744 268346 382800
rect 268382 378392 268438 378448
rect 268474 374312 268530 374368
rect 268566 369960 268622 370016
rect 268658 365880 268714 365936
rect 268750 361528 268806 361584
rect 269026 344936 269082 344992
rect 274546 582800 274602 582856
rect 284022 491292 284078 491328
rect 284022 491272 284024 491292
rect 284024 491272 284076 491292
rect 284076 491272 284078 491292
rect 283838 454008 283894 454064
rect 284022 454028 284078 454064
rect 284022 454008 284024 454028
rect 284024 454008 284076 454028
rect 284076 454008 284078 454028
rect 283838 434696 283894 434752
rect 284022 434716 284078 434752
rect 284022 434696 284024 434716
rect 284024 434696 284076 434716
rect 284076 434696 284078 434716
rect 283838 415384 283894 415440
rect 284022 415404 284078 415440
rect 284022 415384 284024 415404
rect 284024 415384 284076 415404
rect 284076 415384 284078 415404
rect 284114 380160 284170 380216
rect 284114 367104 284170 367160
rect 283930 347928 283986 347984
rect 284114 347792 284170 347848
rect 284298 491272 284354 491328
rect 284114 241440 284170 241496
rect 283654 212472 283710 212528
rect 283930 212472 283986 212528
rect 284298 241440 284354 241496
rect 298006 575728 298062 575784
rect 297454 572736 297510 572792
rect 296626 565800 296682 565856
rect 296534 531392 296590 531448
rect 296902 563352 296958 563408
rect 297270 556824 297326 556880
rect 297362 541048 297418 541104
rect 297178 522144 297234 522200
rect 297270 519152 297326 519208
rect 298006 570016 298062 570072
rect 298006 544040 298062 544096
rect 297638 538328 297694 538384
rect 297914 534792 297970 534848
rect 297454 528808 297510 528864
rect 297822 516180 297878 516216
rect 297822 516160 297824 516180
rect 297824 516160 297876 516180
rect 297876 516160 297878 516180
rect 297822 513440 297878 513496
rect 297730 509632 297786 509688
rect 297730 506640 297786 506696
rect 297730 503784 297786 503840
rect 297638 298016 297694 298072
rect 297638 288496 297694 288552
rect 297362 260752 297418 260808
rect 297546 260752 297602 260808
rect 297362 240080 297418 240136
rect 297546 240080 297602 240136
rect 302790 582936 302846 582992
rect 298834 582664 298890 582720
rect 299294 560360 299350 560416
rect 299202 553560 299258 553616
rect 299110 550704 299166 550760
rect 299018 547848 299074 547904
rect 298926 525816 298982 525872
rect 324134 582528 324190 582584
rect 349526 582392 349582 582448
rect 368662 582800 368718 582856
rect 360198 582664 360254 582720
rect 313278 498072 313334 498128
rect 357438 391312 357494 391368
rect 357438 387812 357440 387832
rect 357440 387812 357492 387832
rect 357492 387812 357494 387832
rect 357438 387776 357494 387812
rect 357438 380976 357494 381032
rect 358542 384512 358598 384568
rect 358082 377712 358138 377768
rect 357438 374176 357494 374232
rect 358082 370912 358138 370968
rect 356702 364112 356758 364168
rect 358174 367376 358230 367432
rect 377402 575456 377458 575512
rect 377310 565800 377366 565856
rect 378138 557164 378194 557220
rect 377494 537512 377550 537568
rect 380714 569064 380770 569120
rect 379702 550704 379758 550760
rect 379518 519152 379574 519208
rect 379518 506504 379574 506560
rect 379518 394576 379574 394632
rect 379610 394440 379666 394496
rect 379794 547032 379850 547088
rect 379886 543768 379942 543824
rect 379978 534520 380034 534576
rect 380070 531392 380126 531448
rect 380162 525000 380218 525056
rect 380254 521736 380310 521792
rect 380346 515480 380402 515536
rect 380438 512488 380494 512544
rect 380530 509496 380586 509552
rect 380622 502968 380678 503024
rect 380806 553424 380862 553480
rect 390650 380160 390706 380216
rect 390650 366832 390706 366888
rect 390926 318688 390982 318744
rect 390926 309168 390982 309224
rect 390926 299376 390982 299432
rect 390926 289856 390982 289912
rect 390926 280064 390982 280120
rect 390926 270544 390982 270600
rect 391938 387504 391994 387560
rect 393410 390768 393466 390824
rect 393318 383968 393374 384024
rect 393318 377168 393374 377224
rect 392030 370368 392086 370424
rect 393410 373904 393466 373960
rect 393502 363568 393558 363624
rect 133786 140392 133842 140448
rect 133970 122984 134026 123040
rect 133878 121896 133934 121952
rect 434258 169632 434314 169688
rect 434534 186224 434590 186280
rect 434994 196152 435050 196208
rect 434902 184592 434958 184648
rect 434810 173848 434866 173904
rect 434718 171944 434774 172000
rect 434442 167728 434498 167784
rect 434350 165552 434406 165608
rect 434166 163512 434222 163568
rect 434074 161200 434130 161256
rect 433982 159296 434038 159352
rect 433890 157256 433946 157312
rect 133878 118088 133934 118144
rect 138202 117408 138258 117464
rect 137926 96600 137982 96656
rect 138202 96600 138258 96656
rect 140778 118632 140834 118688
rect 140778 117272 140834 117328
rect 140962 117272 141018 117328
rect 142802 118632 142858 118688
rect 142802 118088 142858 118144
rect 145562 117816 145618 117872
rect 148046 66408 148102 66464
rect 147954 66272 148010 66328
rect 149058 4800 149114 4856
rect 151818 117680 151874 117736
rect 153474 117952 153530 118008
rect 157246 118632 157302 118688
rect 157246 118088 157302 118144
rect 159086 115912 159142 115968
rect 159638 115912 159694 115968
rect 163042 115912 163098 115968
rect 163410 115912 163466 115968
rect 175646 85584 175702 85640
rect 175830 85448 175886 85504
rect 178222 52400 178278 52456
rect 178406 52400 178462 52456
rect 178130 22072 178186 22128
rect 178406 22072 178462 22128
rect 183650 106256 183706 106312
rect 183926 106256 183982 106312
rect 184754 106256 184810 106312
rect 183742 96600 183798 96656
rect 183926 96600 183982 96656
rect 184938 117544 184994 117600
rect 184938 106256 184994 106312
rect 183742 48320 183798 48376
rect 183650 38664 183706 38720
rect 186594 118496 186650 118552
rect 188434 118088 188490 118144
rect 187790 117272 187846 117328
rect 188434 117272 188490 117328
rect 192022 6160 192078 6216
rect 193954 118360 194010 118416
rect 194690 104760 194746 104816
rect 194966 104624 195022 104680
rect 194966 48320 195022 48376
rect 195150 48320 195206 48376
rect 197634 118224 197690 118280
rect 205914 91024 205970 91080
rect 206098 91024 206154 91080
rect 207294 19352 207350 19408
rect 207294 19216 207350 19272
rect 211250 100680 211306 100736
rect 211434 100544 211490 100600
rect 211158 56752 211214 56808
rect 211250 56480 211306 56536
rect 211342 45464 211398 45520
rect 211526 45464 211582 45520
rect 227994 115912 228050 115968
rect 228270 115912 228326 115968
rect 228914 19216 228970 19272
rect 229098 19216 229154 19272
rect 231122 117952 231178 118008
rect 233422 106256 233478 106312
rect 233606 106256 233662 106312
rect 240230 117952 240286 118008
rect 238942 115912 238998 115968
rect 239310 115912 239366 115968
rect 238758 96736 238814 96792
rect 238850 96620 238906 96656
rect 238850 96600 238852 96620
rect 238852 96600 238904 96620
rect 238904 96600 238906 96620
rect 243542 117272 243598 117328
rect 243450 48320 243506 48376
rect 243450 48184 243506 48240
rect 245750 117272 245806 117328
rect 248970 118088 249026 118144
rect 251546 118088 251602 118144
rect 276110 48320 276166 48376
rect 276294 48320 276350 48376
rect 279790 93880 279846 93936
rect 279974 93880 280030 93936
rect 301870 26288 301926 26344
rect 302054 26288 302110 26344
rect 325514 48320 325570 48376
rect 325698 48320 325754 48376
rect 341062 106256 341118 106312
rect 341246 106256 341302 106312
rect 341062 86944 341118 87000
rect 341246 86944 341302 87000
rect 357346 4800 357402 4856
rect 388718 106276 388774 106312
rect 388718 106256 388720 106276
rect 388720 106256 388772 106276
rect 388772 106256 388774 106276
rect 388902 106256 388958 106312
rect 408314 3712 408370 3768
rect 408498 3712 408554 3768
rect 411074 6160 411130 6216
rect 415030 48320 415086 48376
rect 415214 48320 415270 48376
rect 417882 3576 417938 3632
rect 418342 3576 418398 3632
rect 420274 77288 420330 77344
rect 420458 77288 420514 77344
rect 420642 61376 420698 61432
rect 420550 48320 420606 48376
rect 420642 42064 420698 42120
rect 420550 29008 420606 29064
rect 426070 48320 426126 48376
rect 426254 48320 426310 48376
rect 431590 86944 431646 87000
rect 431774 86944 431830 87000
rect 431590 46960 431646 47016
rect 431774 46960 431830 47016
rect 433982 117952 434038 118008
rect 435178 190168 435234 190224
rect 435086 188808 435142 188864
rect 436190 198872 436246 198928
rect 436098 180240 436154 180296
rect 436098 155080 436154 155136
rect 436098 148688 436154 148744
rect 436098 142060 436100 142080
rect 436100 142060 436152 142080
rect 436152 142060 436154 142080
rect 436098 142024 436154 142060
rect 436282 193976 436338 194032
rect 436650 193024 436706 193080
rect 436558 182008 436614 182064
rect 436466 177928 436522 177984
rect 436374 176160 436430 176216
rect 436742 140392 436798 140448
rect 478510 700440 478566 700496
rect 437386 152768 437442 152824
rect 437386 150184 437442 150240
rect 437386 146240 437442 146296
rect 437018 144472 437074 144528
rect 456798 375128 456854 375184
rect 504730 378392 504786 378448
rect 456798 357992 456854 358048
rect 504730 360440 504786 360496
rect 503718 340856 503774 340912
rect 504730 343576 504786 343632
rect 503902 340856 503958 340912
rect 504270 260888 504326 260944
rect 504638 260888 504694 260944
rect 504362 183504 504418 183560
rect 504638 183504 504694 183560
rect 504178 154536 504234 154592
rect 504454 154536 504510 154592
rect 437386 137808 437442 137864
rect 543462 700304 543518 700360
rect 580170 674600 580226 674656
rect 580170 627680 580226 627736
rect 580170 580760 580226 580816
rect 580262 557232 580318 557288
rect 580170 533840 580226 533896
rect 580170 498616 580226 498672
rect 580170 486784 580226 486840
rect 579802 463392 579858 463448
rect 580170 451696 580226 451752
rect 580170 439864 580226 439920
rect 579802 416472 579858 416528
rect 579986 346024 580042 346080
rect 579618 322632 579674 322688
rect 579710 310800 579766 310856
rect 579618 275712 579674 275768
rect 580170 263880 580226 263936
rect 580170 228792 580226 228848
rect 579618 216960 579674 217016
rect 580354 545536 580410 545592
rect 580446 510312 580502 510368
rect 580630 404776 580686 404832
rect 580538 392944 580594 393000
rect 527178 200640 527234 200696
rect 580262 181872 580318 181928
rect 580262 170040 580318 170096
rect 580170 158344 580226 158400
rect 437018 136040 437074 136096
rect 437386 133592 437442 133648
rect 437386 131960 437442 132016
rect 437386 129512 437442 129568
rect 436834 127744 436890 127800
rect 436926 124480 436982 124536
rect 436834 122848 436890 122904
rect 436742 120400 436798 120456
rect 580722 369552 580778 369608
rect 580814 357856 580870 357912
rect 580630 299104 580686 299160
rect 580354 134816 580410 134872
rect 580722 252184 580778 252240
rect 580814 205264 580870 205320
rect 580538 123120 580594 123176
rect 442262 117952 442318 118008
rect 433522 4800 433578 4856
rect 431222 3304 431278 3360
rect 579802 111424 579858 111480
rect 580170 87896 580226 87952
rect 580170 76200 580226 76256
rect 579802 64504 579858 64560
rect 580170 40976 580226 41032
rect 580170 29280 580226 29336
rect 579802 17584 579858 17640
rect 538126 6160 538182 6216
rect 575018 3304 575074 3360
<< metal3 >>
rect 132166 700436 132172 700500
rect 132236 700498 132242 700500
rect 478505 700498 478571 700501
rect 132236 700496 478571 700498
rect 132236 700440 478510 700496
rect 478566 700440 478571 700496
rect 132236 700438 478571 700440
rect 132236 700436 132242 700438
rect 478505 700435 478571 700438
rect 132350 700300 132356 700364
rect 132420 700362 132426 700364
rect 543457 700362 543523 700365
rect 132420 700360 543523 700362
rect 132420 700304 543462 700360
rect 543518 700304 543523 700360
rect 132420 700302 543523 700304
rect 132420 700300 132426 700302
rect 543457 700299 543523 700302
rect 583520 698050 584960 698140
rect 583342 697990 584960 698050
rect 133638 697172 133644 697236
rect 133708 697234 133714 697236
rect 154481 697234 154547 697237
rect 173801 697234 173867 697237
rect 193121 697234 193187 697237
rect 212441 697234 212507 697237
rect 231761 697234 231827 697237
rect 251081 697234 251147 697237
rect 270401 697234 270467 697237
rect 289721 697234 289787 697237
rect 309041 697234 309107 697237
rect 328361 697234 328427 697237
rect 133708 697174 138122 697234
rect 133708 697172 133714 697174
rect 138062 697098 138122 697174
rect 154481 697232 157442 697234
rect 154481 697176 154486 697232
rect 154542 697176 157442 697232
rect 154481 697174 157442 697176
rect 154481 697171 154547 697174
rect 147581 697098 147647 697101
rect 138062 697096 147647 697098
rect 138062 697040 147586 697096
rect 147642 697040 147647 697096
rect 138062 697038 147647 697040
rect 157382 697098 157442 697174
rect 173801 697232 176762 697234
rect 173801 697176 173806 697232
rect 173862 697176 176762 697232
rect 173801 697174 176762 697176
rect 173801 697171 173867 697174
rect 166901 697098 166967 697101
rect 157382 697096 166967 697098
rect 157382 697040 166906 697096
rect 166962 697040 166967 697096
rect 157382 697038 166967 697040
rect 176702 697098 176762 697174
rect 193121 697232 196082 697234
rect 193121 697176 193126 697232
rect 193182 697176 196082 697232
rect 193121 697174 196082 697176
rect 193121 697171 193187 697174
rect 186221 697098 186287 697101
rect 176702 697096 186287 697098
rect 176702 697040 186226 697096
rect 186282 697040 186287 697096
rect 176702 697038 186287 697040
rect 196022 697098 196082 697174
rect 212441 697232 215402 697234
rect 212441 697176 212446 697232
rect 212502 697176 215402 697232
rect 212441 697174 215402 697176
rect 212441 697171 212507 697174
rect 205541 697098 205607 697101
rect 196022 697096 205607 697098
rect 196022 697040 205546 697096
rect 205602 697040 205607 697096
rect 196022 697038 205607 697040
rect 215342 697098 215402 697174
rect 231761 697232 234722 697234
rect 231761 697176 231766 697232
rect 231822 697176 234722 697232
rect 231761 697174 234722 697176
rect 231761 697171 231827 697174
rect 224861 697098 224927 697101
rect 215342 697096 224927 697098
rect 215342 697040 224866 697096
rect 224922 697040 224927 697096
rect 215342 697038 224927 697040
rect 234662 697098 234722 697174
rect 251081 697232 254042 697234
rect 251081 697176 251086 697232
rect 251142 697176 254042 697232
rect 251081 697174 254042 697176
rect 251081 697171 251147 697174
rect 244181 697098 244247 697101
rect 234662 697096 244247 697098
rect 234662 697040 244186 697096
rect 244242 697040 244247 697096
rect 234662 697038 244247 697040
rect 253982 697098 254042 697174
rect 270401 697232 273362 697234
rect 270401 697176 270406 697232
rect 270462 697176 273362 697232
rect 270401 697174 273362 697176
rect 270401 697171 270467 697174
rect 263501 697098 263567 697101
rect 253982 697096 263567 697098
rect 253982 697040 263506 697096
rect 263562 697040 263567 697096
rect 253982 697038 263567 697040
rect 273302 697098 273362 697174
rect 289721 697232 292682 697234
rect 289721 697176 289726 697232
rect 289782 697176 292682 697232
rect 289721 697174 292682 697176
rect 289721 697171 289787 697174
rect 282821 697098 282887 697101
rect 273302 697096 282887 697098
rect 273302 697040 282826 697096
rect 282882 697040 282887 697096
rect 273302 697038 282887 697040
rect 292622 697098 292682 697174
rect 309041 697232 312002 697234
rect 309041 697176 309046 697232
rect 309102 697176 312002 697232
rect 309041 697174 312002 697176
rect 309041 697171 309107 697174
rect 302141 697098 302207 697101
rect 292622 697096 302207 697098
rect 292622 697040 302146 697096
rect 302202 697040 302207 697096
rect 292622 697038 302207 697040
rect 311942 697098 312002 697174
rect 328361 697232 340890 697234
rect 328361 697176 328366 697232
rect 328422 697176 340890 697232
rect 328361 697174 340890 697176
rect 328361 697171 328427 697174
rect 321461 697098 321527 697101
rect 311942 697096 321527 697098
rect 311942 697040 321466 697096
rect 321522 697040 321527 697096
rect 311942 697038 321527 697040
rect 340830 697098 340890 697174
rect 354630 697174 360210 697234
rect 340830 697038 350458 697098
rect 147581 697035 147647 697038
rect 166901 697035 166967 697038
rect 186221 697035 186287 697038
rect 205541 697035 205607 697038
rect 224861 697035 224927 697038
rect 244181 697035 244247 697038
rect 263501 697035 263567 697038
rect 282821 697035 282887 697038
rect 302141 697035 302207 697038
rect 321461 697035 321527 697038
rect 350398 696962 350458 697038
rect 354630 696962 354690 697174
rect 360150 697098 360210 697174
rect 373950 697174 383578 697234
rect 360150 697038 369778 697098
rect 350398 696902 354690 696962
rect 369718 696962 369778 697038
rect 373950 696962 374010 697174
rect 369718 696902 374010 696962
rect 383518 696962 383578 697174
rect 383702 697174 393330 697234
rect 383702 696962 383762 697174
rect 393270 697098 393330 697174
rect 403022 697174 412650 697234
rect 393270 697038 402898 697098
rect 383518 696902 383762 696962
rect 402838 696962 402898 697038
rect 403022 696962 403082 697174
rect 412590 697098 412650 697174
rect 422342 697174 431970 697234
rect 412590 697038 422218 697098
rect 402838 696902 403082 696962
rect 422158 696962 422218 697038
rect 422342 696962 422402 697174
rect 431910 697098 431970 697174
rect 441662 697174 451290 697234
rect 431910 697038 432154 697098
rect 422158 696902 422402 696962
rect 432094 696962 432154 697038
rect 441662 696962 441722 697174
rect 451230 697098 451290 697174
rect 460982 697174 470610 697234
rect 451230 697038 460858 697098
rect 432094 696902 441722 696962
rect 460798 696962 460858 697038
rect 460982 696962 461042 697174
rect 470550 697098 470610 697174
rect 480302 697174 489930 697234
rect 470550 697038 480178 697098
rect 460798 696902 461042 696962
rect 480118 696962 480178 697038
rect 480302 696962 480362 697174
rect 489870 697098 489930 697174
rect 499622 697174 509250 697234
rect 489870 697038 499498 697098
rect 480118 696902 480362 696962
rect 499438 696962 499498 697038
rect 499622 696962 499682 697174
rect 509190 697098 509250 697174
rect 518942 697174 528570 697234
rect 509190 697038 518818 697098
rect 499438 696902 499682 696962
rect 518758 696962 518818 697038
rect 518942 696962 519002 697174
rect 528510 697098 528570 697174
rect 538262 697174 547890 697234
rect 528510 697038 538138 697098
rect 518758 696902 519002 696962
rect 538078 696962 538138 697038
rect 538262 696962 538322 697174
rect 547830 697098 547890 697174
rect 557582 697174 567210 697234
rect 547830 697038 557458 697098
rect 538078 696902 538322 696962
rect 557398 696962 557458 697038
rect 557582 696962 557642 697174
rect 567150 697098 567210 697174
rect 583342 697098 583402 697990
rect 583520 697900 584960 697990
rect 567150 697038 576778 697098
rect 557398 696902 557642 696962
rect 576718 696962 576778 697038
rect 576902 697038 583402 697098
rect 576902 696962 576962 697038
rect 576718 696902 576962 696962
rect -960 696540 480 696780
rect 164182 686428 164188 686492
rect 164252 686490 164258 686492
rect 169017 686490 169083 686493
rect 164252 686488 169083 686490
rect 164252 686432 169022 686488
rect 169078 686432 169083 686488
rect 164252 686430 169083 686432
rect 164252 686428 164258 686430
rect 169017 686427 169083 686430
rect 147765 686354 147831 686357
rect 154573 686354 154639 686357
rect 583520 686354 584960 686444
rect 147765 686352 154639 686354
rect 147765 686296 147770 686352
rect 147826 686296 154578 686352
rect 154634 686296 154639 686352
rect 147765 686294 154639 686296
rect 147765 686291 147831 686294
rect 154573 686291 154639 686294
rect 583342 686294 584960 686354
rect 135253 686218 135319 686221
rect 132542 686216 135319 686218
rect 132542 686160 135258 686216
rect 135314 686160 135319 686216
rect 132542 686158 135319 686160
rect 131982 685884 131988 685948
rect 132052 685946 132058 685948
rect 132542 685946 132602 686158
rect 135253 686155 135319 686158
rect 159449 686218 159515 686221
rect 164182 686218 164188 686220
rect 159449 686216 164188 686218
rect 159449 686160 159454 686216
rect 159510 686160 164188 686216
rect 159449 686158 164188 686160
rect 159449 686155 159515 686158
rect 164182 686156 164188 686158
rect 164252 686156 164258 686220
rect 169017 686218 169083 686221
rect 169017 686216 180810 686218
rect 169017 686160 169022 686216
rect 169078 686160 180810 686216
rect 169017 686158 180810 686160
rect 169017 686155 169083 686158
rect 147581 686082 147647 686085
rect 144870 686080 147647 686082
rect 144870 686024 147586 686080
rect 147642 686024 147647 686080
rect 144870 686022 147647 686024
rect 180750 686082 180810 686158
rect 190502 686158 200130 686218
rect 180750 686022 190378 686082
rect 132052 685886 132602 685946
rect 142889 685946 142955 685949
rect 144870 685946 144930 686022
rect 147581 686019 147647 686022
rect 142889 685944 144930 685946
rect 142889 685888 142894 685944
rect 142950 685888 144930 685944
rect 142889 685886 144930 685888
rect 190318 685946 190378 686022
rect 190502 685946 190562 686158
rect 200070 686082 200130 686158
rect 209822 686158 219450 686218
rect 200070 686022 209698 686082
rect 190318 685886 190562 685946
rect 209638 685946 209698 686022
rect 209822 685946 209882 686158
rect 219390 686082 219450 686158
rect 229142 686158 238770 686218
rect 219390 686022 229018 686082
rect 209638 685886 209882 685946
rect 228958 685946 229018 686022
rect 229142 685946 229202 686158
rect 238710 686082 238770 686158
rect 248462 686158 258090 686218
rect 238710 686022 248338 686082
rect 228958 685886 229202 685946
rect 248278 685946 248338 686022
rect 248462 685946 248522 686158
rect 258030 686082 258090 686158
rect 267782 686158 277410 686218
rect 258030 686022 267658 686082
rect 248278 685886 248522 685946
rect 267598 685946 267658 686022
rect 267782 685946 267842 686158
rect 277350 686082 277410 686158
rect 287102 686158 296730 686218
rect 277350 686022 286978 686082
rect 267598 685886 267842 685946
rect 286918 685946 286978 686022
rect 287102 685946 287162 686158
rect 296670 686082 296730 686158
rect 306422 686158 316050 686218
rect 296670 686022 306298 686082
rect 286918 685886 287162 685946
rect 306238 685946 306298 686022
rect 306422 685946 306482 686158
rect 315990 686082 316050 686158
rect 325742 686158 335370 686218
rect 315990 686022 325618 686082
rect 306238 685886 306482 685946
rect 325558 685946 325618 686022
rect 325742 685946 325802 686158
rect 335310 686082 335370 686158
rect 345062 686158 354690 686218
rect 335310 686022 344938 686082
rect 325558 685886 325802 685946
rect 344878 685946 344938 686022
rect 345062 685946 345122 686158
rect 354630 686082 354690 686158
rect 364382 686158 374010 686218
rect 354630 686022 364258 686082
rect 344878 685886 345122 685946
rect 364198 685946 364258 686022
rect 364382 685946 364442 686158
rect 373950 686082 374010 686158
rect 383702 686158 393330 686218
rect 373950 686022 383578 686082
rect 364198 685886 364442 685946
rect 383518 685946 383578 686022
rect 383702 685946 383762 686158
rect 393270 686082 393330 686158
rect 403022 686158 412650 686218
rect 393270 686022 402898 686082
rect 383518 685886 383762 685946
rect 402838 685946 402898 686022
rect 403022 685946 403082 686158
rect 412590 686082 412650 686158
rect 422342 686158 431970 686218
rect 412590 686022 422218 686082
rect 402838 685886 403082 685946
rect 422158 685946 422218 686022
rect 422342 685946 422402 686158
rect 431910 686082 431970 686158
rect 441662 686158 451290 686218
rect 431910 686022 441538 686082
rect 422158 685886 422402 685946
rect 441478 685946 441538 686022
rect 441662 685946 441722 686158
rect 451230 686082 451290 686158
rect 460982 686158 470610 686218
rect 451230 686022 460858 686082
rect 441478 685886 441722 685946
rect 460798 685946 460858 686022
rect 460982 685946 461042 686158
rect 470550 686082 470610 686158
rect 480302 686158 489930 686218
rect 470550 686022 480178 686082
rect 460798 685886 461042 685946
rect 480118 685946 480178 686022
rect 480302 685946 480362 686158
rect 489870 686082 489930 686158
rect 499622 686158 509250 686218
rect 489870 686022 499498 686082
rect 480118 685886 480362 685946
rect 499438 685946 499498 686022
rect 499622 685946 499682 686158
rect 509190 686082 509250 686158
rect 518942 686158 528570 686218
rect 509190 686022 518818 686082
rect 499438 685886 499682 685946
rect 518758 685946 518818 686022
rect 518942 685946 519002 686158
rect 528510 686082 528570 686158
rect 538262 686158 547890 686218
rect 528510 686022 538138 686082
rect 518758 685886 519002 685946
rect 538078 685946 538138 686022
rect 538262 685946 538322 686158
rect 547830 686082 547890 686158
rect 557582 686158 567210 686218
rect 547830 686022 557458 686082
rect 538078 685886 538322 685946
rect 557398 685946 557458 686022
rect 557582 685946 557642 686158
rect 567150 686082 567210 686158
rect 583342 686082 583402 686294
rect 583520 686204 584960 686294
rect 567150 686022 576778 686082
rect 557398 685886 557642 685946
rect 576718 685946 576778 686022
rect 576902 686022 583402 686082
rect 576902 685946 576962 686022
rect 576718 685886 576962 685946
rect 132052 685884 132058 685886
rect 142889 685883 142955 685886
rect -960 682274 480 682364
rect 3509 682274 3575 682277
rect -960 682272 3575 682274
rect -960 682216 3514 682272
rect 3570 682216 3575 682272
rect -960 682214 3575 682216
rect -960 682124 480 682214
rect 3509 682211 3575 682214
rect 580165 674658 580231 674661
rect 583520 674658 584960 674748
rect 580165 674656 584960 674658
rect 580165 674600 580170 674656
rect 580226 674600 584960 674656
rect 580165 674598 584960 674600
rect 580165 674595 580231 674598
rect 583520 674508 584960 674598
rect -960 667994 480 668084
rect 3417 667994 3483 667997
rect -960 667992 3483 667994
rect -960 667936 3422 667992
rect 3478 667936 3483 667992
rect -960 667934 3483 667936
rect -960 667844 480 667934
rect 3417 667931 3483 667934
rect 583520 662676 584960 662916
rect -960 653578 480 653668
rect 4797 653578 4863 653581
rect -960 653576 4863 653578
rect -960 653520 4802 653576
rect 4858 653520 4863 653576
rect -960 653518 4863 653520
rect -960 653428 480 653518
rect 4797 653515 4863 653518
rect 583520 651130 584960 651220
rect 583342 651070 584960 651130
rect 164182 650524 164188 650588
rect 164252 650586 164258 650588
rect 169017 650586 169083 650589
rect 164252 650584 169083 650586
rect 164252 650528 169022 650584
rect 169078 650528 169083 650584
rect 164252 650526 169083 650528
rect 164252 650524 164258 650526
rect 169017 650523 169083 650526
rect 147765 650450 147831 650453
rect 154573 650450 154639 650453
rect 147765 650448 154639 650450
rect 147765 650392 147770 650448
rect 147826 650392 154578 650448
rect 154634 650392 154639 650448
rect 147765 650390 154639 650392
rect 147765 650387 147831 650390
rect 154573 650387 154639 650390
rect 133454 650252 133460 650316
rect 133524 650314 133530 650316
rect 135253 650314 135319 650317
rect 133524 650312 135319 650314
rect 133524 650256 135258 650312
rect 135314 650256 135319 650312
rect 133524 650254 135319 650256
rect 133524 650252 133530 650254
rect 135253 650251 135319 650254
rect 159449 650314 159515 650317
rect 164182 650314 164188 650316
rect 159449 650312 164188 650314
rect 159449 650256 159454 650312
rect 159510 650256 164188 650312
rect 159449 650254 164188 650256
rect 159449 650251 159515 650254
rect 164182 650252 164188 650254
rect 164252 650252 164258 650316
rect 169017 650314 169083 650317
rect 169017 650312 180810 650314
rect 169017 650256 169022 650312
rect 169078 650256 180810 650312
rect 169017 650254 180810 650256
rect 169017 650251 169083 650254
rect 147581 650178 147647 650181
rect 144870 650176 147647 650178
rect 144870 650120 147586 650176
rect 147642 650120 147647 650176
rect 144870 650118 147647 650120
rect 180750 650178 180810 650254
rect 190502 650254 200130 650314
rect 180750 650118 190378 650178
rect 142889 650042 142955 650045
rect 144870 650042 144930 650118
rect 147581 650115 147647 650118
rect 142889 650040 144930 650042
rect 142889 649984 142894 650040
rect 142950 649984 144930 650040
rect 142889 649982 144930 649984
rect 190318 650042 190378 650118
rect 190502 650042 190562 650254
rect 200070 650178 200130 650254
rect 209822 650254 219450 650314
rect 200070 650118 209698 650178
rect 190318 649982 190562 650042
rect 209638 650042 209698 650118
rect 209822 650042 209882 650254
rect 219390 650178 219450 650254
rect 229142 650254 238770 650314
rect 219390 650118 229018 650178
rect 209638 649982 209882 650042
rect 228958 650042 229018 650118
rect 229142 650042 229202 650254
rect 238710 650178 238770 650254
rect 248462 650254 258090 650314
rect 238710 650118 248338 650178
rect 228958 649982 229202 650042
rect 248278 650042 248338 650118
rect 248462 650042 248522 650254
rect 258030 650178 258090 650254
rect 267782 650254 277410 650314
rect 258030 650118 267658 650178
rect 248278 649982 248522 650042
rect 267598 650042 267658 650118
rect 267782 650042 267842 650254
rect 277350 650178 277410 650254
rect 287102 650254 296730 650314
rect 277350 650118 286978 650178
rect 267598 649982 267842 650042
rect 286918 650042 286978 650118
rect 287102 650042 287162 650254
rect 296670 650178 296730 650254
rect 306422 650254 316050 650314
rect 296670 650118 306298 650178
rect 286918 649982 287162 650042
rect 306238 650042 306298 650118
rect 306422 650042 306482 650254
rect 315990 650178 316050 650254
rect 325742 650254 335370 650314
rect 315990 650118 325618 650178
rect 306238 649982 306482 650042
rect 325558 650042 325618 650118
rect 325742 650042 325802 650254
rect 335310 650178 335370 650254
rect 345062 650254 354690 650314
rect 335310 650118 344938 650178
rect 325558 649982 325802 650042
rect 344878 650042 344938 650118
rect 345062 650042 345122 650254
rect 354630 650178 354690 650254
rect 364382 650254 374010 650314
rect 354630 650118 364258 650178
rect 344878 649982 345122 650042
rect 364198 650042 364258 650118
rect 364382 650042 364442 650254
rect 373950 650178 374010 650254
rect 383702 650254 393330 650314
rect 373950 650118 383578 650178
rect 364198 649982 364442 650042
rect 383518 650042 383578 650118
rect 383702 650042 383762 650254
rect 393270 650178 393330 650254
rect 403022 650254 412650 650314
rect 393270 650118 402898 650178
rect 383518 649982 383762 650042
rect 402838 650042 402898 650118
rect 403022 650042 403082 650254
rect 412590 650178 412650 650254
rect 422342 650254 431970 650314
rect 412590 650118 422218 650178
rect 402838 649982 403082 650042
rect 422158 650042 422218 650118
rect 422342 650042 422402 650254
rect 431910 650178 431970 650254
rect 441662 650254 451290 650314
rect 431910 650118 441538 650178
rect 422158 649982 422402 650042
rect 441478 650042 441538 650118
rect 441662 650042 441722 650254
rect 451230 650178 451290 650254
rect 460982 650254 470610 650314
rect 451230 650118 460858 650178
rect 441478 649982 441722 650042
rect 460798 650042 460858 650118
rect 460982 650042 461042 650254
rect 470550 650178 470610 650254
rect 480302 650254 489930 650314
rect 470550 650118 480178 650178
rect 460798 649982 461042 650042
rect 480118 650042 480178 650118
rect 480302 650042 480362 650254
rect 489870 650178 489930 650254
rect 499622 650254 509250 650314
rect 489870 650118 499498 650178
rect 480118 649982 480362 650042
rect 499438 650042 499498 650118
rect 499622 650042 499682 650254
rect 509190 650178 509250 650254
rect 518942 650254 528570 650314
rect 509190 650118 518818 650178
rect 499438 649982 499682 650042
rect 518758 650042 518818 650118
rect 518942 650042 519002 650254
rect 528510 650178 528570 650254
rect 538262 650254 547890 650314
rect 528510 650118 538138 650178
rect 518758 649982 519002 650042
rect 538078 650042 538138 650118
rect 538262 650042 538322 650254
rect 547830 650178 547890 650254
rect 557582 650254 567210 650314
rect 547830 650118 557458 650178
rect 538078 649982 538322 650042
rect 557398 650042 557458 650118
rect 557582 650042 557642 650254
rect 567150 650178 567210 650254
rect 583342 650178 583402 651070
rect 583520 650980 584960 651070
rect 567150 650118 576778 650178
rect 557398 649982 557642 650042
rect 576718 650042 576778 650118
rect 576902 650118 583402 650178
rect 576902 650042 576962 650118
rect 576718 649982 576962 650042
rect 142889 649979 142955 649982
rect 583520 639434 584960 639524
rect 583342 639374 584960 639434
rect 157057 639298 157123 639301
rect 132542 639296 157123 639298
rect -960 639012 480 639252
rect 132542 639240 157062 639296
rect 157118 639240 157123 639296
rect 132542 639238 157123 639240
rect 131798 638964 131804 639028
rect 131868 639026 131874 639028
rect 132542 639026 132602 639238
rect 157057 639235 157123 639238
rect 157241 639298 157307 639301
rect 171041 639298 171107 639301
rect 157241 639296 159282 639298
rect 157241 639240 157246 639296
rect 157302 639240 159282 639296
rect 157241 639238 159282 639240
rect 157241 639235 157307 639238
rect 159222 639162 159282 639238
rect 171041 639296 180810 639298
rect 171041 639240 171046 639296
rect 171102 639240 180810 639296
rect 171041 639238 180810 639240
rect 171041 639235 171107 639238
rect 164182 639162 164188 639164
rect 159222 639102 164188 639162
rect 164182 639100 164188 639102
rect 164252 639100 164258 639164
rect 180750 639162 180810 639238
rect 190502 639238 200130 639298
rect 180750 639102 190378 639162
rect 131868 638966 132602 639026
rect 190318 639026 190378 639102
rect 190502 639026 190562 639238
rect 200070 639162 200130 639238
rect 209822 639238 219450 639298
rect 200070 639102 209698 639162
rect 190318 638966 190562 639026
rect 209638 639026 209698 639102
rect 209822 639026 209882 639238
rect 219390 639162 219450 639238
rect 229142 639238 238770 639298
rect 219390 639102 229018 639162
rect 209638 638966 209882 639026
rect 228958 639026 229018 639102
rect 229142 639026 229202 639238
rect 238710 639162 238770 639238
rect 248462 639238 258090 639298
rect 238710 639102 248338 639162
rect 228958 638966 229202 639026
rect 248278 639026 248338 639102
rect 248462 639026 248522 639238
rect 258030 639162 258090 639238
rect 267782 639238 277410 639298
rect 258030 639102 267658 639162
rect 248278 638966 248522 639026
rect 267598 639026 267658 639102
rect 267782 639026 267842 639238
rect 277350 639162 277410 639238
rect 287102 639238 296730 639298
rect 277350 639102 286978 639162
rect 267598 638966 267842 639026
rect 286918 639026 286978 639102
rect 287102 639026 287162 639238
rect 296670 639162 296730 639238
rect 306422 639238 316050 639298
rect 296670 639102 306298 639162
rect 286918 638966 287162 639026
rect 306238 639026 306298 639102
rect 306422 639026 306482 639238
rect 315990 639162 316050 639238
rect 325742 639238 335370 639298
rect 315990 639102 325618 639162
rect 306238 638966 306482 639026
rect 325558 639026 325618 639102
rect 325742 639026 325802 639238
rect 335310 639162 335370 639238
rect 345062 639238 354690 639298
rect 335310 639102 344938 639162
rect 325558 638966 325802 639026
rect 344878 639026 344938 639102
rect 345062 639026 345122 639238
rect 354630 639162 354690 639238
rect 364382 639238 374010 639298
rect 354630 639102 364258 639162
rect 344878 638966 345122 639026
rect 364198 639026 364258 639102
rect 364382 639026 364442 639238
rect 373950 639162 374010 639238
rect 383702 639238 393330 639298
rect 373950 639102 383578 639162
rect 364198 638966 364442 639026
rect 383518 639026 383578 639102
rect 383702 639026 383762 639238
rect 393270 639162 393330 639238
rect 403022 639238 412650 639298
rect 393270 639102 402898 639162
rect 383518 638966 383762 639026
rect 402838 639026 402898 639102
rect 403022 639026 403082 639238
rect 412590 639162 412650 639238
rect 422342 639238 431970 639298
rect 412590 639102 422218 639162
rect 402838 638966 403082 639026
rect 422158 639026 422218 639102
rect 422342 639026 422402 639238
rect 431910 639162 431970 639238
rect 441662 639238 451290 639298
rect 431910 639102 441538 639162
rect 422158 638966 422402 639026
rect 441478 639026 441538 639102
rect 441662 639026 441722 639238
rect 451230 639162 451290 639238
rect 460982 639238 470610 639298
rect 451230 639102 460858 639162
rect 441478 638966 441722 639026
rect 460798 639026 460858 639102
rect 460982 639026 461042 639238
rect 470550 639162 470610 639238
rect 480302 639238 489930 639298
rect 470550 639102 480178 639162
rect 460798 638966 461042 639026
rect 480118 639026 480178 639102
rect 480302 639026 480362 639238
rect 489870 639162 489930 639238
rect 499622 639238 509250 639298
rect 489870 639102 499498 639162
rect 480118 638966 480362 639026
rect 499438 639026 499498 639102
rect 499622 639026 499682 639238
rect 509190 639162 509250 639238
rect 518942 639238 528570 639298
rect 509190 639102 518818 639162
rect 499438 638966 499682 639026
rect 518758 639026 518818 639102
rect 518942 639026 519002 639238
rect 528510 639162 528570 639238
rect 538262 639238 547890 639298
rect 528510 639102 538138 639162
rect 518758 638966 519002 639026
rect 538078 639026 538138 639102
rect 538262 639026 538322 639238
rect 547830 639162 547890 639238
rect 557582 639238 567210 639298
rect 547830 639102 557458 639162
rect 538078 638966 538322 639026
rect 557398 639026 557458 639102
rect 557582 639026 557642 639238
rect 567150 639162 567210 639238
rect 583342 639162 583402 639374
rect 583520 639284 584960 639374
rect 567150 639102 576778 639162
rect 557398 638966 557642 639026
rect 576718 639026 576778 639102
rect 576902 639102 583402 639162
rect 576902 639026 576962 639102
rect 576718 638966 576962 639026
rect 131868 638964 131874 638966
rect 164182 638828 164188 638892
rect 164252 638890 164258 638892
rect 171041 638890 171107 638893
rect 164252 638888 171107 638890
rect 164252 638832 171046 638888
rect 171102 638832 171107 638888
rect 164252 638830 171107 638832
rect 164252 638828 164258 638830
rect 171041 638827 171107 638830
rect 580165 627738 580231 627741
rect 583520 627738 584960 627828
rect 580165 627736 584960 627738
rect 580165 627680 580170 627736
rect 580226 627680 584960 627736
rect 580165 627678 584960 627680
rect 580165 627675 580231 627678
rect 583520 627588 584960 627678
rect -960 624882 480 624972
rect 3417 624882 3483 624885
rect -960 624880 3483 624882
rect -960 624824 3422 624880
rect 3478 624824 3483 624880
rect -960 624822 3483 624824
rect -960 624732 480 624822
rect 3417 624819 3483 624822
rect 583520 615756 584960 615996
rect -960 610466 480 610556
rect 3417 610466 3483 610469
rect -960 610464 3483 610466
rect -960 610408 3422 610464
rect 3478 610408 3483 610464
rect -960 610406 3483 610408
rect -960 610316 480 610406
rect 3417 610403 3483 610406
rect 583520 604210 584960 604300
rect 583342 604150 584960 604210
rect 133086 603332 133092 603396
rect 133156 603394 133162 603396
rect 157057 603394 157123 603397
rect 133156 603392 157123 603394
rect 133156 603336 157062 603392
rect 157118 603336 157123 603392
rect 133156 603334 157123 603336
rect 133156 603332 133162 603334
rect 157057 603331 157123 603334
rect 157241 603394 157307 603397
rect 171041 603394 171107 603397
rect 157241 603392 159466 603394
rect 157241 603336 157246 603392
rect 157302 603336 159466 603392
rect 157241 603334 159466 603336
rect 157241 603331 157307 603334
rect 159406 603258 159466 603334
rect 171041 603392 180810 603394
rect 171041 603336 171046 603392
rect 171102 603336 180810 603392
rect 171041 603334 180810 603336
rect 171041 603331 171107 603334
rect 164182 603258 164188 603260
rect 159406 603198 164188 603258
rect 164182 603196 164188 603198
rect 164252 603196 164258 603260
rect 180750 603258 180810 603334
rect 190502 603334 200130 603394
rect 180750 603198 190378 603258
rect 190318 603122 190378 603198
rect 190502 603122 190562 603334
rect 200070 603258 200130 603334
rect 209822 603334 219450 603394
rect 200070 603198 209698 603258
rect 190318 603062 190562 603122
rect 209638 603122 209698 603198
rect 209822 603122 209882 603334
rect 219390 603258 219450 603334
rect 229142 603334 238770 603394
rect 219390 603198 229018 603258
rect 209638 603062 209882 603122
rect 228958 603122 229018 603198
rect 229142 603122 229202 603334
rect 238710 603258 238770 603334
rect 248462 603334 258090 603394
rect 238710 603198 248338 603258
rect 228958 603062 229202 603122
rect 248278 603122 248338 603198
rect 248462 603122 248522 603334
rect 258030 603258 258090 603334
rect 267782 603334 277410 603394
rect 258030 603198 267658 603258
rect 248278 603062 248522 603122
rect 267598 603122 267658 603198
rect 267782 603122 267842 603334
rect 277350 603258 277410 603334
rect 287102 603334 296730 603394
rect 277350 603198 286978 603258
rect 267598 603062 267842 603122
rect 286918 603122 286978 603198
rect 287102 603122 287162 603334
rect 296670 603258 296730 603334
rect 306422 603334 316050 603394
rect 296670 603198 306298 603258
rect 286918 603062 287162 603122
rect 306238 603122 306298 603198
rect 306422 603122 306482 603334
rect 315990 603258 316050 603334
rect 325742 603334 335370 603394
rect 315990 603198 325618 603258
rect 306238 603062 306482 603122
rect 325558 603122 325618 603198
rect 325742 603122 325802 603334
rect 335310 603258 335370 603334
rect 345062 603334 354690 603394
rect 335310 603198 344938 603258
rect 325558 603062 325802 603122
rect 344878 603122 344938 603198
rect 345062 603122 345122 603334
rect 354630 603258 354690 603334
rect 364382 603334 374010 603394
rect 354630 603198 364258 603258
rect 344878 603062 345122 603122
rect 364198 603122 364258 603198
rect 364382 603122 364442 603334
rect 373950 603258 374010 603334
rect 383702 603334 393330 603394
rect 373950 603198 383578 603258
rect 364198 603062 364442 603122
rect 383518 603122 383578 603198
rect 383702 603122 383762 603334
rect 393270 603258 393330 603334
rect 403022 603334 412650 603394
rect 393270 603198 402898 603258
rect 383518 603062 383762 603122
rect 402838 603122 402898 603198
rect 403022 603122 403082 603334
rect 412590 603258 412650 603334
rect 422342 603334 431970 603394
rect 412590 603198 422218 603258
rect 402838 603062 403082 603122
rect 422158 603122 422218 603198
rect 422342 603122 422402 603334
rect 431910 603258 431970 603334
rect 441662 603334 451290 603394
rect 431910 603198 441538 603258
rect 422158 603062 422402 603122
rect 441478 603122 441538 603198
rect 441662 603122 441722 603334
rect 451230 603258 451290 603334
rect 460982 603334 470610 603394
rect 451230 603198 460858 603258
rect 441478 603062 441722 603122
rect 460798 603122 460858 603198
rect 460982 603122 461042 603334
rect 470550 603258 470610 603334
rect 480302 603334 489930 603394
rect 470550 603198 480178 603258
rect 460798 603062 461042 603122
rect 480118 603122 480178 603198
rect 480302 603122 480362 603334
rect 489870 603258 489930 603334
rect 499622 603334 509250 603394
rect 489870 603198 499498 603258
rect 480118 603062 480362 603122
rect 499438 603122 499498 603198
rect 499622 603122 499682 603334
rect 509190 603258 509250 603334
rect 518942 603334 528570 603394
rect 509190 603198 518818 603258
rect 499438 603062 499682 603122
rect 518758 603122 518818 603198
rect 518942 603122 519002 603334
rect 528510 603258 528570 603334
rect 538262 603334 547890 603394
rect 528510 603198 538138 603258
rect 518758 603062 519002 603122
rect 538078 603122 538138 603198
rect 538262 603122 538322 603334
rect 547830 603258 547890 603334
rect 557582 603334 567210 603394
rect 547830 603198 557458 603258
rect 538078 603062 538322 603122
rect 557398 603122 557458 603198
rect 557582 603122 557642 603334
rect 567150 603258 567210 603334
rect 583342 603258 583402 604150
rect 583520 604060 584960 604150
rect 567150 603198 576778 603258
rect 557398 603062 557642 603122
rect 576718 603122 576778 603198
rect 576902 603198 583402 603258
rect 576902 603122 576962 603198
rect 576718 603062 576962 603122
rect 164182 602924 164188 602988
rect 164252 602986 164258 602988
rect 171041 602986 171107 602989
rect 164252 602984 171107 602986
rect 164252 602928 171046 602984
rect 171102 602928 171107 602984
rect 164252 602926 171107 602928
rect 164252 602924 164258 602926
rect 171041 602923 171107 602926
rect -960 596050 480 596140
rect 4061 596050 4127 596053
rect -960 596048 4127 596050
rect -960 595992 4066 596048
rect 4122 595992 4127 596048
rect -960 595990 4127 595992
rect -960 595900 480 595990
rect 4061 595987 4127 595990
rect 164182 592588 164188 592652
rect 164252 592650 164258 592652
rect 169017 592650 169083 592653
rect 164252 592648 169083 592650
rect 164252 592592 169022 592648
rect 169078 592592 169083 592648
rect 164252 592590 169083 592592
rect 164252 592588 164258 592590
rect 169017 592587 169083 592590
rect 147765 592514 147831 592517
rect 154573 592514 154639 592517
rect 583520 592514 584960 592604
rect 147765 592512 154639 592514
rect 147765 592456 147770 592512
rect 147826 592456 154578 592512
rect 154634 592456 154639 592512
rect 147765 592454 154639 592456
rect 147765 592451 147831 592454
rect 154573 592451 154639 592454
rect 583342 592454 584960 592514
rect 133270 592316 133276 592380
rect 133340 592378 133346 592380
rect 135253 592378 135319 592381
rect 133340 592376 135319 592378
rect 133340 592320 135258 592376
rect 135314 592320 135319 592376
rect 133340 592318 135319 592320
rect 133340 592316 133346 592318
rect 135253 592315 135319 592318
rect 159449 592378 159515 592381
rect 164182 592378 164188 592380
rect 159449 592376 164188 592378
rect 159449 592320 159454 592376
rect 159510 592320 164188 592376
rect 159449 592318 164188 592320
rect 159449 592315 159515 592318
rect 164182 592316 164188 592318
rect 164252 592316 164258 592380
rect 169017 592378 169083 592381
rect 169017 592376 180810 592378
rect 169017 592320 169022 592376
rect 169078 592320 180810 592376
rect 169017 592318 180810 592320
rect 169017 592315 169083 592318
rect 147581 592242 147647 592245
rect 144870 592240 147647 592242
rect 144870 592184 147586 592240
rect 147642 592184 147647 592240
rect 144870 592182 147647 592184
rect 180750 592242 180810 592318
rect 190502 592318 200130 592378
rect 180750 592182 190378 592242
rect 142889 592106 142955 592109
rect 144870 592106 144930 592182
rect 147581 592179 147647 592182
rect 142889 592104 144930 592106
rect 142889 592048 142894 592104
rect 142950 592048 144930 592104
rect 142889 592046 144930 592048
rect 190318 592106 190378 592182
rect 190502 592106 190562 592318
rect 200070 592242 200130 592318
rect 209822 592318 219450 592378
rect 200070 592182 209698 592242
rect 190318 592046 190562 592106
rect 209638 592106 209698 592182
rect 209822 592106 209882 592318
rect 219390 592242 219450 592318
rect 229142 592318 238770 592378
rect 219390 592182 229018 592242
rect 209638 592046 209882 592106
rect 228958 592106 229018 592182
rect 229142 592106 229202 592318
rect 238710 592242 238770 592318
rect 248462 592318 258090 592378
rect 238710 592182 248338 592242
rect 228958 592046 229202 592106
rect 248278 592106 248338 592182
rect 248462 592106 248522 592318
rect 258030 592242 258090 592318
rect 267782 592318 277410 592378
rect 258030 592182 267658 592242
rect 248278 592046 248522 592106
rect 267598 592106 267658 592182
rect 267782 592106 267842 592318
rect 277350 592242 277410 592318
rect 287102 592318 296730 592378
rect 277350 592182 286978 592242
rect 267598 592046 267842 592106
rect 286918 592106 286978 592182
rect 287102 592106 287162 592318
rect 296670 592242 296730 592318
rect 306422 592318 316050 592378
rect 296670 592182 306298 592242
rect 286918 592046 287162 592106
rect 306238 592106 306298 592182
rect 306422 592106 306482 592318
rect 315990 592242 316050 592318
rect 325742 592318 335370 592378
rect 315990 592182 325618 592242
rect 306238 592046 306482 592106
rect 325558 592106 325618 592182
rect 325742 592106 325802 592318
rect 335310 592242 335370 592318
rect 345062 592318 354690 592378
rect 335310 592182 344938 592242
rect 325558 592046 325802 592106
rect 344878 592106 344938 592182
rect 345062 592106 345122 592318
rect 354630 592242 354690 592318
rect 364382 592318 374010 592378
rect 354630 592182 364258 592242
rect 344878 592046 345122 592106
rect 364198 592106 364258 592182
rect 364382 592106 364442 592318
rect 373950 592242 374010 592318
rect 383702 592318 393330 592378
rect 373950 592182 383578 592242
rect 364198 592046 364442 592106
rect 383518 592106 383578 592182
rect 383702 592106 383762 592318
rect 393270 592242 393330 592318
rect 403022 592318 412650 592378
rect 393270 592182 402898 592242
rect 383518 592046 383762 592106
rect 402838 592106 402898 592182
rect 403022 592106 403082 592318
rect 412590 592242 412650 592318
rect 422342 592318 431970 592378
rect 412590 592182 422218 592242
rect 402838 592046 403082 592106
rect 422158 592106 422218 592182
rect 422342 592106 422402 592318
rect 431910 592242 431970 592318
rect 441662 592318 451290 592378
rect 431910 592182 441538 592242
rect 422158 592046 422402 592106
rect 441478 592106 441538 592182
rect 441662 592106 441722 592318
rect 451230 592242 451290 592318
rect 460982 592318 470610 592378
rect 451230 592182 460858 592242
rect 441478 592046 441722 592106
rect 460798 592106 460858 592182
rect 460982 592106 461042 592318
rect 470550 592242 470610 592318
rect 480302 592318 489930 592378
rect 470550 592182 480178 592242
rect 460798 592046 461042 592106
rect 480118 592106 480178 592182
rect 480302 592106 480362 592318
rect 489870 592242 489930 592318
rect 499622 592318 509250 592378
rect 489870 592182 499498 592242
rect 480118 592046 480362 592106
rect 499438 592106 499498 592182
rect 499622 592106 499682 592318
rect 509190 592242 509250 592318
rect 518942 592318 528570 592378
rect 509190 592182 518818 592242
rect 499438 592046 499682 592106
rect 518758 592106 518818 592182
rect 518942 592106 519002 592318
rect 528510 592242 528570 592318
rect 538262 592318 547890 592378
rect 528510 592182 538138 592242
rect 518758 592046 519002 592106
rect 538078 592106 538138 592182
rect 538262 592106 538322 592318
rect 547830 592242 547890 592318
rect 557582 592318 567210 592378
rect 547830 592182 557458 592242
rect 538078 592046 538322 592106
rect 557398 592106 557458 592182
rect 557582 592106 557642 592318
rect 567150 592242 567210 592318
rect 583342 592242 583402 592454
rect 583520 592364 584960 592454
rect 567150 592182 576778 592242
rect 557398 592046 557642 592106
rect 576718 592106 576778 592182
rect 576902 592182 583402 592242
rect 576902 592106 576962 592182
rect 576718 592046 576962 592106
rect 142889 592043 142955 592046
rect 191097 582994 191163 582997
rect 302785 582994 302851 582997
rect 191097 582992 302851 582994
rect 191097 582936 191102 582992
rect 191158 582936 302790 582992
rect 302846 582936 302851 582992
rect 191097 582934 302851 582936
rect 191097 582931 191163 582934
rect 302785 582931 302851 582934
rect 274541 582858 274607 582861
rect 368657 582858 368723 582861
rect 274541 582856 368723 582858
rect 274541 582800 274546 582856
rect 274602 582800 368662 582856
rect 368718 582800 368723 582856
rect 274541 582798 368723 582800
rect 274541 582795 274607 582798
rect 368657 582795 368723 582798
rect 298829 582722 298895 582725
rect 360193 582722 360259 582725
rect 298829 582720 360259 582722
rect 298829 582664 298834 582720
rect 298890 582664 360198 582720
rect 360254 582664 360259 582720
rect 298829 582662 360259 582664
rect 298829 582659 298895 582662
rect 360193 582659 360259 582662
rect 124857 582586 124923 582589
rect 324129 582586 324195 582589
rect 124857 582584 324195 582586
rect 124857 582528 124862 582584
rect 124918 582528 324134 582584
rect 324190 582528 324195 582584
rect 124857 582526 324195 582528
rect 124857 582523 124923 582526
rect 324129 582523 324195 582526
rect 131021 582450 131087 582453
rect 349521 582450 349587 582453
rect 131021 582448 349587 582450
rect 131021 582392 131026 582448
rect 131082 582392 349526 582448
rect 349582 582392 349587 582448
rect 131021 582390 349587 582392
rect 131021 582387 131087 582390
rect 349521 582387 349587 582390
rect -960 581620 480 581860
rect 580165 580818 580231 580821
rect 583520 580818 584960 580908
rect 580165 580816 584960 580818
rect 580165 580760 580170 580816
rect 580226 580760 584960 580816
rect 580165 580758 584960 580760
rect 580165 580755 580231 580758
rect 583520 580668 584960 580758
rect 298001 575786 298067 575789
rect 299982 575786 300042 576232
rect 298001 575784 300042 575786
rect 298001 575728 298006 575784
rect 298062 575728 300042 575784
rect 298001 575726 300042 575728
rect 298001 575723 298067 575726
rect 377446 575517 377506 575960
rect 377397 575512 377506 575517
rect 377397 575456 377402 575512
rect 377458 575456 377506 575512
rect 377397 575454 377506 575456
rect 377397 575451 377463 575454
rect 297449 572794 297515 572797
rect 299982 572794 300042 572968
rect 297449 572792 300042 572794
rect 297449 572736 297454 572792
rect 297510 572736 300042 572792
rect 297449 572734 300042 572736
rect 297449 572731 297515 572734
rect 377814 572114 377874 572696
rect 380014 572114 380020 572116
rect 377814 572054 380020 572114
rect 380014 572052 380020 572054
rect 380084 572052 380090 572116
rect 298001 570074 298067 570077
rect 298001 570072 300042 570074
rect 298001 570016 298006 570072
rect 298062 570016 300042 570072
rect 298001 570014 300042 570016
rect 298001 570011 298067 570014
rect 299982 569976 300042 570014
rect 377814 569122 377874 569704
rect 380709 569122 380775 569125
rect 377814 569120 380775 569122
rect 377814 569064 380714 569120
rect 380770 569064 380775 569120
rect 377814 569062 380775 569064
rect 380709 569059 380775 569062
rect 583520 568836 584960 569076
rect -960 567354 480 567444
rect 3417 567354 3483 567357
rect -960 567352 3483 567354
rect -960 567296 3422 567352
rect 3478 567296 3483 567352
rect -960 567294 3483 567296
rect -960 567204 480 567294
rect 3417 567291 3483 567294
rect 296621 565858 296687 565861
rect 299982 565858 300042 566712
rect 296621 565856 300042 565858
rect 296621 565800 296626 565856
rect 296682 565800 300042 565856
rect 296621 565798 300042 565800
rect 377262 565861 377322 566440
rect 377262 565856 377371 565861
rect 377262 565800 377310 565856
rect 377366 565800 377371 565856
rect 377262 565798 377371 565800
rect 296621 565795 296687 565798
rect 377305 565795 377371 565798
rect 296897 563410 296963 563413
rect 299982 563410 300042 563720
rect 296897 563408 300042 563410
rect 296897 563352 296902 563408
rect 296958 563352 300042 563408
rect 296897 563350 300042 563352
rect 296897 563347 296963 563350
rect 377814 563138 377874 563448
rect 379462 563138 379468 563140
rect 377814 563078 379468 563138
rect 379462 563076 379468 563078
rect 379532 563076 379538 563140
rect 199694 561716 199700 561780
rect 199764 561778 199770 561780
rect 211613 561778 211679 561781
rect 199764 561776 211679 561778
rect 199764 561720 211618 561776
rect 211674 561720 211679 561776
rect 199764 561718 211679 561720
rect 199764 561716 199770 561718
rect 211613 561715 211679 561718
rect 299289 560418 299355 560421
rect 299982 560418 300042 560456
rect 299289 560416 300042 560418
rect 299289 560360 299294 560416
rect 299350 560360 300042 560416
rect 299289 560358 300042 560360
rect 299289 560355 299355 560358
rect 377814 559602 377874 560184
rect 379646 559602 379652 559604
rect 377814 559542 379652 559602
rect 379646 559540 379652 559542
rect 379716 559540 379722 559604
rect 198590 556684 198596 556748
rect 198660 556746 198666 556748
rect 200070 556746 200130 557328
rect 297265 556882 297331 556885
rect 299982 556882 300042 557464
rect 580257 557290 580323 557293
rect 583520 557290 584960 557380
rect 580257 557288 584960 557290
rect 580257 557232 580262 557288
rect 580318 557232 584960 557288
rect 580257 557230 584960 557232
rect 580257 557227 580323 557230
rect 378133 557222 378199 557225
rect 377844 557220 378199 557222
rect 377844 557164 378138 557220
rect 378194 557164 378199 557220
rect 377844 557162 378199 557164
rect 378133 557159 378199 557162
rect 583520 557140 584960 557230
rect 297265 556880 300042 556882
rect 297265 556824 297270 556880
rect 297326 556824 300042 556880
rect 297265 556822 300042 556824
rect 297265 556819 297331 556822
rect 198660 556686 200130 556746
rect 198660 556684 198666 556686
rect 219942 556202 220002 556784
rect 222193 556202 222259 556205
rect 219942 556200 222259 556202
rect 219942 556144 222198 556200
rect 222254 556144 222259 556200
rect 219942 556142 222259 556144
rect 222193 556139 222259 556142
rect 299197 553618 299263 553621
rect 299982 553618 300042 554200
rect 299197 553616 300042 553618
rect 299197 553560 299202 553616
rect 299258 553560 300042 553616
rect 299197 553558 300042 553560
rect 299197 553555 299263 553558
rect 377814 553482 377874 553928
rect 380801 553482 380867 553485
rect 377814 553480 380867 553482
rect 377814 553424 380806 553480
rect 380862 553424 380867 553480
rect 377814 553422 380867 553424
rect 380801 553419 380867 553422
rect -960 553074 480 553164
rect 3141 553074 3207 553077
rect -960 553072 3207 553074
rect -960 553016 3146 553072
rect 3202 553016 3207 553072
rect -960 553014 3207 553016
rect -960 552924 480 553014
rect 3141 553011 3207 553014
rect 198406 552060 198412 552124
rect 198476 552122 198482 552124
rect 200070 552122 200130 552704
rect 198476 552062 200130 552122
rect 219942 552122 220002 552160
rect 222285 552122 222351 552125
rect 219942 552120 222351 552122
rect 219942 552064 222290 552120
rect 222346 552064 222351 552120
rect 219942 552062 222351 552064
rect 198476 552060 198482 552062
rect 222285 552059 222351 552062
rect 299105 550762 299171 550765
rect 299982 550762 300042 550936
rect 379697 550762 379763 550765
rect 299105 550760 300042 550762
rect 299105 550704 299110 550760
rect 299166 550704 300042 550760
rect 299105 550702 300042 550704
rect 377814 550760 379763 550762
rect 377814 550704 379702 550760
rect 379758 550704 379763 550760
rect 377814 550702 379763 550704
rect 299105 550699 299171 550702
rect 377814 550664 377874 550702
rect 379697 550699 379763 550702
rect 86358 549949 86418 550528
rect 86358 549944 86467 549949
rect 86358 549888 86406 549944
rect 86462 549888 86467 549944
rect 86358 549886 86467 549888
rect 86401 549883 86467 549886
rect 198222 547844 198228 547908
rect 198292 547906 198298 547908
rect 200070 547906 200130 548080
rect 198292 547846 200130 547906
rect 299013 547906 299079 547909
rect 299982 547906 300042 547944
rect 299013 547904 300042 547906
rect 299013 547848 299018 547904
rect 299074 547848 300042 547904
rect 299013 547846 300042 547848
rect 198292 547844 198298 547846
rect 299013 547843 299079 547846
rect 219942 546954 220002 547536
rect 377814 547090 377874 547672
rect 379789 547090 379855 547093
rect 377814 547088 379855 547090
rect 377814 547032 379794 547088
rect 379850 547032 379855 547088
rect 377814 547030 379855 547032
rect 379789 547027 379855 547030
rect 222561 546954 222627 546957
rect 219942 546952 222627 546954
rect 219942 546896 222566 546952
rect 222622 546896 222627 546952
rect 219942 546894 222627 546896
rect 222561 546891 222627 546894
rect 115614 546546 115674 546720
rect 118049 546546 118115 546549
rect 115614 546544 118115 546546
rect 115614 546488 118054 546544
rect 118110 546488 118115 546544
rect 115614 546486 118115 546488
rect 118049 546483 118115 546486
rect 84101 545866 84167 545869
rect 85990 545866 86050 546448
rect 84101 545864 86050 545866
rect 84101 545808 84106 545864
rect 84162 545808 86050 545864
rect 84101 545806 86050 545808
rect 84101 545803 84167 545806
rect 580349 545594 580415 545597
rect 583520 545594 584960 545684
rect 580349 545592 584960 545594
rect 580349 545536 580354 545592
rect 580410 545536 584960 545592
rect 580349 545534 584960 545536
rect 580349 545531 580415 545534
rect 583520 545444 584960 545534
rect 298001 544098 298067 544101
rect 299982 544098 300042 544680
rect 298001 544096 300042 544098
rect 298001 544040 298006 544096
rect 298062 544040 300042 544096
rect 298001 544038 300042 544040
rect 298001 544035 298067 544038
rect 198038 543764 198044 543828
rect 198108 543826 198114 543828
rect 377814 543826 377874 544408
rect 379881 543826 379947 543829
rect 198108 543766 200130 543826
rect 377814 543824 379947 543826
rect 377814 543768 379886 543824
rect 379942 543768 379947 543824
rect 377814 543766 379947 543768
rect 198108 543764 198114 543766
rect 200070 543728 200130 543766
rect 379881 543763 379947 543766
rect 219942 542602 220002 543184
rect 222469 542602 222535 542605
rect 219942 542600 222535 542602
rect 219942 542544 222474 542600
rect 222530 542544 222535 542600
rect 219942 542542 222535 542544
rect 222469 542539 222535 542542
rect 118601 542466 118667 542469
rect 115614 542464 118667 542466
rect 115614 542408 118606 542464
rect 118662 542408 118667 542464
rect 115614 542406 118667 542408
rect 115614 542368 115674 542406
rect 118601 542403 118667 542406
rect 84009 541514 84075 541517
rect 85990 541514 86050 542096
rect 84009 541512 86050 541514
rect 84009 541456 84014 541512
rect 84070 541456 86050 541512
rect 84009 541454 86050 541456
rect 84009 541451 84075 541454
rect 297357 541106 297423 541109
rect 299982 541106 300042 541688
rect 297357 541104 300042 541106
rect 297357 541048 297362 541104
rect 297418 541048 300042 541104
rect 297357 541046 300042 541048
rect 377814 541106 377874 541416
rect 380198 541106 380204 541108
rect 377814 541046 380204 541106
rect 297357 541043 297423 541046
rect 380198 541044 380204 541046
rect 380268 541044 380274 541108
rect -960 538658 480 538748
rect 3509 538658 3575 538661
rect -960 538656 3575 538658
rect -960 538600 3514 538656
rect 3570 538600 3575 538656
rect -960 538598 3575 538600
rect -960 538508 480 538598
rect 3509 538595 3575 538598
rect 197854 538460 197860 538524
rect 197924 538522 197930 538524
rect 200070 538522 200130 539104
rect 197924 538462 200130 538522
rect 197924 538460 197930 538462
rect 219942 538386 220002 538560
rect 222377 538386 222443 538389
rect 219942 538384 222443 538386
rect 219942 538328 222382 538384
rect 222438 538328 222443 538384
rect 219942 538326 222443 538328
rect 222377 538323 222443 538326
rect 297633 538386 297699 538389
rect 299982 538386 300042 538424
rect 297633 538384 300042 538386
rect 297633 538328 297638 538384
rect 297694 538328 300042 538384
rect 297633 538326 300042 538328
rect 297633 538323 297699 538326
rect 85297 537162 85363 537165
rect 85990 537162 86050 537744
rect 115614 537434 115674 538016
rect 377446 537573 377506 538152
rect 377446 537568 377555 537573
rect 377446 537512 377494 537568
rect 377550 537512 377555 537568
rect 377446 537510 377555 537512
rect 377489 537507 377555 537510
rect 117773 537434 117839 537437
rect 115614 537432 117839 537434
rect 115614 537376 117778 537432
rect 117834 537376 117839 537432
rect 115614 537374 117839 537376
rect 117773 537371 117839 537374
rect 85297 537160 86050 537162
rect 85297 537104 85302 537160
rect 85358 537104 86050 537160
rect 85297 537102 86050 537104
rect 85297 537099 85363 537102
rect 297909 534850 297975 534853
rect 299982 534850 300042 535432
rect 297909 534848 300042 534850
rect 297909 534792 297914 534848
rect 297970 534792 300042 534848
rect 297909 534790 300042 534792
rect 297909 534787 297975 534790
rect 377814 534578 377874 535160
rect 379973 534578 380039 534581
rect 377814 534576 380039 534578
rect 377814 534520 379978 534576
rect 380034 534520 380039 534576
rect 377814 534518 380039 534520
rect 379973 534515 380039 534518
rect 198641 534170 198707 534173
rect 200070 534170 200130 534480
rect 198641 534168 200130 534170
rect 198641 534112 198646 534168
rect 198702 534112 200130 534168
rect 198641 534110 200130 534112
rect 198641 534107 198707 534110
rect 85205 533082 85271 533085
rect 85990 533082 86050 533664
rect 115614 533354 115674 533936
rect 117773 533354 117839 533357
rect 115614 533352 117839 533354
rect 115614 533296 117778 533352
rect 117834 533296 117839 533352
rect 115614 533294 117839 533296
rect 219942 533354 220002 533936
rect 580165 533898 580231 533901
rect 583520 533898 584960 533988
rect 580165 533896 584960 533898
rect 580165 533840 580170 533896
rect 580226 533840 584960 533896
rect 580165 533838 584960 533840
rect 580165 533835 580231 533838
rect 583520 533748 584960 533838
rect 222653 533354 222719 533357
rect 219942 533352 222719 533354
rect 219942 533296 222658 533352
rect 222714 533296 222719 533352
rect 219942 533294 222719 533296
rect 117773 533291 117839 533294
rect 222653 533291 222719 533294
rect 85205 533080 86050 533082
rect 85205 533024 85210 533080
rect 85266 533024 86050 533080
rect 85205 533022 86050 533024
rect 85205 533019 85271 533022
rect 296529 531450 296595 531453
rect 299982 531450 300042 532168
rect 296529 531448 300042 531450
rect 296529 531392 296534 531448
rect 296590 531392 300042 531448
rect 296529 531390 300042 531392
rect 377814 531450 377874 531896
rect 380065 531450 380131 531453
rect 377814 531448 380131 531450
rect 377814 531392 380070 531448
rect 380126 531392 380131 531448
rect 377814 531390 380131 531392
rect 296529 531387 296595 531390
rect 380065 531387 380131 531390
rect 117957 529682 118023 529685
rect 115614 529680 118023 529682
rect 115614 529624 117962 529680
rect 118018 529624 118023 529680
rect 115614 529622 118023 529624
rect 115614 529584 115674 529622
rect 117957 529619 118023 529622
rect 83917 528730 83983 528733
rect 85990 528730 86050 529312
rect 198733 529274 198799 529277
rect 200070 529274 200130 529856
rect 198733 529272 200130 529274
rect 198733 529216 198738 529272
rect 198794 529216 200130 529272
rect 198733 529214 200130 529216
rect 198733 529211 198799 529214
rect 219942 529002 220002 529312
rect 222745 529002 222811 529005
rect 219942 529000 222811 529002
rect 219942 528944 222750 529000
rect 222806 528944 222811 529000
rect 219942 528942 222811 528944
rect 222745 528939 222811 528942
rect 297449 528866 297515 528869
rect 299982 528866 300042 529176
rect 297449 528864 300042 528866
rect 297449 528808 297454 528864
rect 297510 528808 300042 528864
rect 297449 528806 300042 528808
rect 297449 528803 297515 528806
rect 83917 528728 86050 528730
rect 83917 528672 83922 528728
rect 83978 528672 86050 528728
rect 83917 528670 86050 528672
rect 377814 528730 377874 528904
rect 379830 528730 379836 528732
rect 377814 528670 379836 528730
rect 83917 528667 83983 528670
rect 379830 528668 379836 528670
rect 379900 528668 379906 528732
rect 298921 525874 298987 525877
rect 299982 525874 300042 525912
rect 298921 525872 300042 525874
rect 298921 525816 298926 525872
rect 298982 525816 300042 525872
rect 298921 525814 300042 525816
rect 298921 525811 298987 525814
rect 85389 525602 85455 525605
rect 85389 525600 86050 525602
rect 85389 525544 85394 525600
rect 85450 525544 86050 525600
rect 85389 525542 86050 525544
rect 85389 525539 85455 525542
rect 82813 524922 82879 524925
rect 85990 524922 86050 525542
rect 115614 525194 115674 525232
rect 118601 525194 118667 525197
rect 115614 525192 118667 525194
rect 115614 525136 118606 525192
rect 118662 525136 118667 525192
rect 115614 525134 118667 525136
rect 118601 525131 118667 525134
rect 82813 524920 86050 524922
rect 82813 524864 82818 524920
rect 82874 524864 86050 524920
rect 82813 524862 86050 524864
rect 82813 524859 82879 524862
rect 198549 524650 198615 524653
rect 200070 524650 200130 525232
rect 377814 525058 377874 525640
rect 380157 525058 380223 525061
rect 377814 525056 380223 525058
rect 377814 525000 380162 525056
rect 380218 525000 380223 525056
rect 377814 524998 380223 525000
rect 380157 524995 380223 524998
rect 198549 524648 200130 524650
rect 198549 524592 198554 524648
rect 198610 524592 200130 524648
rect 198549 524590 200130 524592
rect 198549 524587 198615 524590
rect 219942 524514 220002 524688
rect 222837 524514 222903 524517
rect 219942 524512 222903 524514
rect 219942 524456 222842 524512
rect 222898 524456 222903 524512
rect 219942 524454 222903 524456
rect 222837 524451 222903 524454
rect -960 524092 480 524332
rect 297173 522202 297239 522205
rect 299982 522202 300042 522648
rect 297173 522200 300042 522202
rect 297173 522144 297178 522200
rect 297234 522144 300042 522200
rect 297173 522142 300042 522144
rect 297173 522139 297239 522142
rect 377814 521794 377874 522376
rect 583520 521916 584960 522156
rect 380249 521794 380315 521797
rect 377814 521792 380315 521794
rect 377814 521736 380254 521792
rect 380310 521736 380315 521792
rect 377814 521734 380315 521736
rect 380249 521731 380315 521734
rect 153285 521658 153351 521661
rect 153469 521658 153535 521661
rect 153285 521656 153535 521658
rect 153285 521600 153290 521656
rect 153346 521600 153474 521656
rect 153530 521600 153535 521656
rect 153285 521598 153535 521600
rect 153285 521595 153351 521598
rect 153469 521595 153535 521598
rect 115614 521114 115674 521152
rect 117313 521114 117379 521117
rect 115614 521112 117379 521114
rect 115614 521056 117318 521112
rect 117374 521056 117379 521112
rect 115614 521054 117379 521056
rect 117313 521051 117379 521054
rect 297265 519210 297331 519213
rect 299982 519210 300042 519656
rect 297265 519208 300042 519210
rect 297265 519152 297270 519208
rect 297326 519152 300042 519208
rect 297265 519150 300042 519152
rect 377814 519210 377874 519384
rect 379513 519210 379579 519213
rect 377814 519208 379579 519210
rect 377814 519152 379518 519208
rect 379574 519152 379579 519208
rect 377814 519150 379579 519152
rect 297265 519147 297331 519150
rect 379513 519147 379579 519150
rect 297817 516218 297883 516221
rect 299982 516218 300042 516392
rect 297817 516216 300042 516218
rect 297817 516160 297822 516216
rect 297878 516160 300042 516216
rect 297817 516158 300042 516160
rect 297817 516155 297883 516158
rect 377814 515538 377874 516120
rect 380341 515538 380407 515541
rect 377814 515536 380407 515538
rect 377814 515480 380346 515536
rect 380402 515480 380407 515536
rect 377814 515478 380407 515480
rect 380341 515475 380407 515478
rect 297817 513498 297883 513501
rect 297817 513496 300042 513498
rect 297817 513440 297822 513496
rect 297878 513440 300042 513496
rect 297817 513438 300042 513440
rect 297817 513435 297883 513438
rect 299982 513400 300042 513438
rect 377814 512546 377874 513128
rect 380433 512546 380499 512549
rect 377814 512544 380499 512546
rect 377814 512488 380438 512544
rect 380494 512488 380499 512544
rect 377814 512486 380499 512488
rect 380433 512483 380499 512486
rect 580441 510370 580507 510373
rect 583520 510370 584960 510460
rect 580441 510368 584960 510370
rect 580441 510312 580446 510368
rect 580502 510312 584960 510368
rect 580441 510310 584960 510312
rect 580441 510307 580507 510310
rect 583520 510220 584960 510310
rect -960 509962 480 510052
rect 3601 509962 3667 509965
rect -960 509960 3667 509962
rect -960 509904 3606 509960
rect 3662 509904 3667 509960
rect -960 509902 3667 509904
rect -960 509812 480 509902
rect 3601 509899 3667 509902
rect 297725 509690 297791 509693
rect 299982 509690 300042 510136
rect 297725 509688 300042 509690
rect 297725 509632 297730 509688
rect 297786 509632 300042 509688
rect 297725 509630 300042 509632
rect 297725 509627 297791 509630
rect 377814 509554 377874 509864
rect 380525 509554 380591 509557
rect 377814 509552 380591 509554
rect 377814 509496 380530 509552
rect 380586 509496 380591 509552
rect 377814 509494 380591 509496
rect 380525 509491 380591 509494
rect 297725 506698 297791 506701
rect 299982 506698 300042 507144
rect 297725 506696 300042 506698
rect 297725 506640 297730 506696
rect 297786 506640 300042 506696
rect 297725 506638 300042 506640
rect 297725 506635 297791 506638
rect 377814 506562 377874 506872
rect 379513 506562 379579 506565
rect 377814 506560 379579 506562
rect 377814 506504 379518 506560
rect 379574 506504 379579 506560
rect 377814 506502 379579 506504
rect 379513 506499 379579 506502
rect 297725 503842 297791 503845
rect 299982 503842 300042 503880
rect 297725 503840 300042 503842
rect 297725 503784 297730 503840
rect 297786 503784 300042 503840
rect 297725 503782 300042 503784
rect 297725 503779 297791 503782
rect 377814 503026 377874 503608
rect 380617 503026 380683 503029
rect 377814 503024 380683 503026
rect 377814 502968 380622 503024
rect 380678 502968 380683 503024
rect 377814 502966 380683 502968
rect 380617 502963 380683 502966
rect 130929 500306 130995 500309
rect 380198 500306 380204 500308
rect 130929 500304 380204 500306
rect 130929 500248 130934 500304
rect 130990 500248 380204 500304
rect 130929 500246 380204 500248
rect 130929 500243 130995 500246
rect 380198 500244 380204 500246
rect 380268 500244 380274 500308
rect 129549 500170 129615 500173
rect 380014 500170 380020 500172
rect 129549 500168 380020 500170
rect 129549 500112 129554 500168
rect 129610 500112 380020 500168
rect 129549 500110 380020 500112
rect 129549 500107 129615 500110
rect 380014 500108 380020 500110
rect 380084 500108 380090 500172
rect 580165 498674 580231 498677
rect 583520 498674 584960 498764
rect 580165 498672 584960 498674
rect 580165 498616 580170 498672
rect 580226 498616 584960 498672
rect 580165 498614 584960 498616
rect 580165 498611 580231 498614
rect 583520 498524 584960 498614
rect 115289 498130 115355 498133
rect 313273 498130 313339 498133
rect 115289 498128 313339 498130
rect 115289 498072 115294 498128
rect 115350 498072 313278 498128
rect 313334 498072 313339 498128
rect 115289 498070 313339 498072
rect 115289 498067 115355 498070
rect 313273 498067 313339 498070
rect -960 495546 480 495636
rect 3325 495546 3391 495549
rect 125961 495548 126027 495549
rect 125910 495546 125916 495548
rect -960 495544 3391 495546
rect -960 495488 3330 495544
rect 3386 495488 3391 495544
rect -960 495486 3391 495488
rect 125870 495486 125916 495546
rect 125980 495544 126027 495548
rect 126022 495488 126027 495544
rect -960 495396 480 495486
rect 3325 495483 3391 495486
rect 125910 495484 125916 495486
rect 125980 495484 126027 495488
rect 125961 495483 126027 495484
rect 125869 492692 125935 492693
rect 125869 492688 125916 492692
rect 125980 492690 125986 492692
rect 125869 492632 125874 492688
rect 125869 492628 125916 492632
rect 125980 492630 126026 492690
rect 125980 492628 125986 492630
rect 125869 492627 125935 492628
rect 284017 491330 284083 491333
rect 284293 491330 284359 491333
rect 284017 491328 284359 491330
rect 284017 491272 284022 491328
rect 284078 491272 284298 491328
rect 284354 491272 284359 491328
rect 284017 491270 284359 491272
rect 284017 491267 284083 491270
rect 284293 491267 284359 491270
rect 580165 486842 580231 486845
rect 583520 486842 584960 486932
rect 580165 486840 584960 486842
rect 580165 486784 580170 486840
rect 580226 486784 584960 486840
rect 580165 486782 584960 486784
rect 580165 486779 580231 486782
rect 583520 486692 584960 486782
rect 153285 483034 153351 483037
rect 153469 483034 153535 483037
rect 153285 483032 153535 483034
rect 153285 482976 153290 483032
rect 153346 482976 153474 483032
rect 153530 482976 153535 483032
rect 153285 482974 153535 482976
rect 153285 482971 153351 482974
rect 153469 482971 153535 482974
rect 128629 481674 128695 481677
rect 128813 481674 128879 481677
rect 128629 481672 128879 481674
rect 128629 481616 128634 481672
rect 128690 481616 128818 481672
rect 128874 481616 128879 481672
rect 128629 481614 128879 481616
rect 128629 481611 128695 481614
rect 128813 481611 128879 481614
rect -960 481130 480 481220
rect 4061 481130 4127 481133
rect -960 481128 4127 481130
rect -960 481072 4066 481128
rect 4122 481072 4127 481128
rect -960 481070 4127 481072
rect -960 480980 480 481070
rect 4061 481067 4127 481070
rect 583520 474996 584960 475236
rect -960 466700 480 466940
rect 128537 463722 128603 463725
rect 128813 463722 128879 463725
rect 128537 463720 128879 463722
rect 128537 463664 128542 463720
rect 128598 463664 128818 463720
rect 128874 463664 128879 463720
rect 128537 463662 128879 463664
rect 128537 463659 128603 463662
rect 128813 463659 128879 463662
rect 579797 463450 579863 463453
rect 583520 463450 584960 463540
rect 579797 463448 584960 463450
rect 579797 463392 579802 463448
rect 579858 463392 584960 463448
rect 579797 463390 584960 463392
rect 579797 463387 579863 463390
rect 583520 463300 584960 463390
rect 283833 454066 283899 454069
rect 284017 454066 284083 454069
rect 283833 454064 284083 454066
rect 283833 454008 283838 454064
rect 283894 454008 284022 454064
rect 284078 454008 284083 454064
rect 283833 454006 284083 454008
rect 283833 454003 283899 454006
rect 284017 454003 284083 454006
rect -960 452434 480 452524
rect 3049 452434 3115 452437
rect -960 452432 3115 452434
rect -960 452376 3054 452432
rect 3110 452376 3115 452432
rect -960 452374 3115 452376
rect -960 452284 480 452374
rect 3049 452371 3115 452374
rect 580165 451754 580231 451757
rect 583520 451754 584960 451844
rect 580165 451752 584960 451754
rect 580165 451696 580170 451752
rect 580226 451696 584960 451752
rect 580165 451694 584960 451696
rect 580165 451691 580231 451694
rect 583520 451604 584960 451694
rect 153377 447268 153443 447269
rect 153326 447266 153332 447268
rect 153286 447206 153332 447266
rect 153396 447264 153443 447268
rect 153438 447208 153443 447264
rect 153326 447204 153332 447206
rect 153396 447204 153443 447208
rect 153377 447203 153443 447204
rect 128537 444410 128603 444413
rect 128813 444410 128879 444413
rect 153377 444412 153443 444413
rect 128537 444408 128879 444410
rect 128537 444352 128542 444408
rect 128598 444352 128818 444408
rect 128874 444352 128879 444408
rect 128537 444350 128879 444352
rect 128537 444347 128603 444350
rect 128813 444347 128879 444350
rect 153326 444348 153332 444412
rect 153396 444410 153443 444412
rect 153396 444408 153488 444410
rect 153438 444352 153488 444408
rect 153396 444350 153488 444352
rect 153396 444348 153443 444350
rect 153377 444347 153443 444348
rect 580165 439922 580231 439925
rect 583520 439922 584960 440012
rect 580165 439920 584960 439922
rect 580165 439864 580170 439920
rect 580226 439864 584960 439920
rect 580165 439862 584960 439864
rect 580165 439859 580231 439862
rect 583520 439772 584960 439862
rect -960 438018 480 438108
rect 3693 438018 3759 438021
rect -960 438016 3759 438018
rect -960 437960 3698 438016
rect 3754 437960 3759 438016
rect -960 437958 3759 437960
rect -960 437868 480 437958
rect 3693 437955 3759 437958
rect 283833 434754 283899 434757
rect 284017 434754 284083 434757
rect 283833 434752 284083 434754
rect 283833 434696 283838 434752
rect 283894 434696 284022 434752
rect 284078 434696 284083 434752
rect 283833 434694 284083 434696
rect 283833 434691 283899 434694
rect 284017 434691 284083 434694
rect 583520 428076 584960 428316
rect 153469 425234 153535 425237
rect 153150 425232 153535 425234
rect 153150 425176 153474 425232
rect 153530 425176 153535 425232
rect 153150 425174 153535 425176
rect 153150 425101 153210 425174
rect 153469 425171 153535 425174
rect 128537 425098 128603 425101
rect 128813 425098 128879 425101
rect 128537 425096 128879 425098
rect 128537 425040 128542 425096
rect 128598 425040 128818 425096
rect 128874 425040 128879 425096
rect 128537 425038 128879 425040
rect 153150 425096 153259 425101
rect 153150 425040 153198 425096
rect 153254 425040 153259 425096
rect 153150 425038 153259 425040
rect 128537 425035 128603 425038
rect 128813 425035 128879 425038
rect 153193 425035 153259 425038
rect -960 423738 480 423828
rect 4061 423738 4127 423741
rect -960 423736 4127 423738
rect -960 423680 4066 423736
rect 4122 423680 4127 423736
rect -960 423678 4127 423680
rect -960 423588 480 423678
rect 4061 423675 4127 423678
rect 126421 417482 126487 417485
rect 379830 417482 379836 417484
rect 126421 417480 379836 417482
rect 126421 417424 126426 417480
rect 126482 417424 379836 417480
rect 126421 417422 379836 417424
rect 126421 417419 126487 417422
rect 379830 417420 379836 417422
rect 379900 417420 379906 417484
rect 579797 416530 579863 416533
rect 583520 416530 584960 416620
rect 579797 416528 584960 416530
rect 579797 416472 579802 416528
rect 579858 416472 584960 416528
rect 579797 416470 584960 416472
rect 579797 416467 579863 416470
rect 583520 416380 584960 416470
rect 125869 415442 125935 415445
rect 126145 415442 126211 415445
rect 125869 415440 126211 415442
rect 125869 415384 125874 415440
rect 125930 415384 126150 415440
rect 126206 415384 126211 415440
rect 125869 415382 126211 415384
rect 125869 415379 125935 415382
rect 126145 415379 126211 415382
rect 283833 415442 283899 415445
rect 284017 415442 284083 415445
rect 283833 415440 284083 415442
rect 283833 415384 283838 415440
rect 283894 415384 284022 415440
rect 284078 415384 284083 415440
rect 283833 415382 284083 415384
rect 283833 415379 283899 415382
rect 284017 415379 284083 415382
rect 203333 410410 203399 410413
rect 266854 410410 266860 410412
rect 203333 410408 266860 410410
rect 203333 410352 203338 410408
rect 203394 410352 266860 410408
rect 203333 410350 266860 410352
rect 203333 410347 203399 410350
rect 266854 410348 266860 410350
rect 266924 410348 266930 410412
rect 231853 410274 231919 410277
rect 267774 410274 267780 410276
rect 231853 410272 267780 410274
rect 231853 410216 231858 410272
rect 231914 410216 267780 410272
rect 231853 410214 267780 410216
rect 231853 410211 231919 410214
rect 267774 410212 267780 410214
rect 267844 410212 267850 410276
rect 226149 410138 226215 410141
rect 267958 410138 267964 410140
rect 226149 410136 267964 410138
rect 226149 410080 226154 410136
rect 226210 410080 267964 410136
rect 226149 410078 267964 410080
rect 226149 410075 226215 410078
rect 267958 410076 267964 410078
rect 268028 410076 268034 410140
rect 263133 410002 263199 410005
rect 268142 410002 268148 410004
rect 263133 410000 268148 410002
rect 263133 409944 263138 410000
rect 263194 409944 268148 410000
rect 263133 409942 268148 409944
rect 263133 409939 263199 409942
rect 268142 409940 268148 409942
rect 268212 409940 268218 410004
rect -960 409172 480 409412
rect 580625 404834 580691 404837
rect 583520 404834 584960 404924
rect 580625 404832 584960 404834
rect 580625 404776 580630 404832
rect 580686 404776 584960 404832
rect 580625 404774 584960 404776
rect 580625 404771 580691 404774
rect 583520 404684 584960 404774
rect 198825 403746 198891 403749
rect 267917 403746 267983 403749
rect 198825 403744 200100 403746
rect 198825 403688 198830 403744
rect 198886 403688 200100 403744
rect 198825 403686 200100 403688
rect 266524 403744 267983 403746
rect 266524 403688 267922 403744
rect 267978 403688 267983 403744
rect 266524 403686 267983 403688
rect 198825 403683 198891 403686
rect 267917 403683 267983 403686
rect 198457 399666 198523 399669
rect 266905 399666 266971 399669
rect 198457 399664 200100 399666
rect 198457 399608 198462 399664
rect 198518 399608 200100 399664
rect 198457 399606 200100 399608
rect 266524 399664 266971 399666
rect 266524 399608 266910 399664
rect 266966 399608 266971 399664
rect 266524 399606 266971 399608
rect 198457 399603 198523 399606
rect 266905 399603 266971 399606
rect 125685 395722 125751 395725
rect 126053 395722 126119 395725
rect 126881 395722 126947 395725
rect 125685 395720 126947 395722
rect 125685 395664 125690 395720
rect 125746 395664 126058 395720
rect 126114 395664 126886 395720
rect 126942 395664 126947 395720
rect 125685 395662 126947 395664
rect 125685 395659 125751 395662
rect 126053 395659 126119 395662
rect 126881 395659 126947 395662
rect 198917 395314 198983 395317
rect 268009 395314 268075 395317
rect 198917 395312 200100 395314
rect 198917 395256 198922 395312
rect 198978 395256 200100 395312
rect 198917 395254 200100 395256
rect 266524 395312 268075 395314
rect 266524 395256 268014 395312
rect 268070 395256 268075 395312
rect 266524 395254 268075 395256
rect 198917 395251 198983 395254
rect 268009 395251 268075 395254
rect -960 395042 480 395132
rect 3877 395042 3943 395045
rect -960 395040 3943 395042
rect -960 394984 3882 395040
rect 3938 394984 3943 395040
rect -960 394982 3943 394984
rect -960 394892 480 394982
rect 3877 394979 3943 394982
rect 379513 394636 379579 394637
rect 379462 394634 379468 394636
rect 379422 394574 379468 394634
rect 379532 394632 379579 394636
rect 379574 394576 379579 394632
rect 379462 394572 379468 394574
rect 379532 394572 379579 394576
rect 379513 394571 379579 394572
rect 379605 394500 379671 394501
rect 379605 394498 379652 394500
rect 379560 394496 379652 394498
rect 379560 394440 379610 394496
rect 379560 394438 379652 394440
rect 379605 394436 379652 394438
rect 379716 394436 379722 394500
rect 379605 394435 379671 394436
rect 580533 393002 580599 393005
rect 583520 393002 584960 393092
rect 580533 393000 584960 393002
rect 580533 392944 580538 393000
rect 580594 392944 584960 393000
rect 580533 392942 584960 392944
rect 580533 392939 580599 392942
rect 583520 392852 584960 392942
rect 70301 392594 70367 392597
rect 71589 392594 71655 392597
rect 70301 392592 72036 392594
rect 70301 392536 70306 392592
rect 70362 392536 71594 392592
rect 71650 392536 72036 392592
rect 70301 392534 72036 392536
rect 70301 392531 70367 392534
rect 71589 392531 71655 392534
rect 357433 391370 357499 391373
rect 357433 391368 360180 391370
rect 357433 391312 357438 391368
rect 357494 391312 360180 391368
rect 357433 391310 360180 391312
rect 357433 391307 357499 391310
rect 199009 391234 199075 391237
rect 268101 391234 268167 391237
rect 199009 391232 200100 391234
rect 199009 391176 199014 391232
rect 199070 391176 200100 391232
rect 199009 391174 200100 391176
rect 266524 391232 268167 391234
rect 266524 391176 268106 391232
rect 268162 391176 268167 391232
rect 266524 391174 268167 391176
rect 199009 391171 199075 391174
rect 268101 391171 268167 391174
rect 393405 390826 393471 390829
rect 391092 390824 393471 390826
rect 391092 390768 393410 390824
rect 393466 390768 393471 390824
rect 391092 390766 393471 390768
rect 393405 390763 393471 390766
rect 128629 388242 128695 388245
rect 125734 388240 128695 388242
rect 125734 388184 128634 388240
rect 128690 388184 128695 388240
rect 125734 388182 128695 388184
rect 125734 387940 125794 388182
rect 128629 388179 128695 388182
rect 357433 387834 357499 387837
rect 357433 387832 360180 387834
rect 357433 387776 357438 387832
rect 357494 387776 360180 387832
rect 357433 387774 360180 387776
rect 357433 387771 357499 387774
rect 391933 387562 391999 387565
rect 391092 387560 391999 387562
rect 391092 387504 391938 387560
rect 391994 387504 391999 387560
rect 391092 387502 391999 387504
rect 391933 387499 391999 387502
rect 198365 387154 198431 387157
rect 198365 387152 200100 387154
rect 198365 387096 198370 387152
rect 198426 387096 200100 387152
rect 198365 387094 200100 387096
rect 198365 387091 198431 387094
rect 268193 386882 268259 386885
rect 266524 386880 268259 386882
rect 266524 386824 268198 386880
rect 268254 386824 268259 386880
rect 266524 386822 268259 386824
rect 268193 386819 268259 386822
rect 69933 385250 69999 385253
rect 69933 385248 72036 385250
rect 69933 385192 69938 385248
rect 69994 385192 72036 385248
rect 69933 385190 72036 385192
rect 69933 385187 69999 385190
rect 358537 384570 358603 384573
rect 358537 384568 360180 384570
rect 358537 384512 358542 384568
rect 358598 384512 360180 384568
rect 358537 384510 360180 384512
rect 358537 384507 358603 384510
rect 393313 384026 393379 384029
rect 391092 384024 393379 384026
rect 391092 383968 393318 384024
rect 393374 383968 393379 384024
rect 391092 383966 393379 383968
rect 393313 383963 393379 383966
rect 199101 382802 199167 382805
rect 268285 382802 268351 382805
rect 199101 382800 200100 382802
rect 199101 382744 199106 382800
rect 199162 382744 200100 382800
rect 199101 382742 200100 382744
rect 266524 382800 268351 382802
rect 266524 382744 268290 382800
rect 268346 382744 268351 382800
rect 266524 382742 268351 382744
rect 199101 382739 199167 382742
rect 268285 382739 268351 382742
rect 583520 381156 584960 381396
rect 357433 381034 357499 381037
rect 357433 381032 360180 381034
rect 357433 380976 357438 381032
rect 357494 380976 360180 381032
rect 357433 380974 360180 380976
rect 357433 380971 357499 380974
rect -960 380626 480 380716
rect 3785 380626 3851 380629
rect 129089 380626 129155 380629
rect -960 380624 3851 380626
rect -960 380568 3790 380624
rect 3846 380568 3851 380624
rect -960 380566 3851 380568
rect 126132 380624 129155 380626
rect 126132 380568 129094 380624
rect 129150 380568 129155 380624
rect 126132 380566 129155 380568
rect -960 380476 480 380566
rect 3785 380563 3851 380566
rect 129089 380563 129155 380566
rect 390694 380221 390754 380732
rect 283966 380156 283972 380220
rect 284036 380218 284042 380220
rect 284109 380218 284175 380221
rect 284036 380216 284175 380218
rect 284036 380160 284114 380216
rect 284170 380160 284175 380216
rect 284036 380158 284175 380160
rect 284036 380156 284042 380158
rect 284109 380155 284175 380158
rect 390645 380216 390754 380221
rect 390645 380160 390650 380216
rect 390706 380160 390754 380216
rect 390645 380158 390754 380160
rect 390645 380155 390711 380158
rect 197997 378722 198063 378725
rect 197997 378720 200100 378722
rect 197997 378664 198002 378720
rect 198058 378664 200100 378720
rect 197997 378662 200100 378664
rect 197997 378659 198063 378662
rect 268377 378450 268443 378453
rect 266524 378448 268443 378450
rect 266524 378392 268382 378448
rect 268438 378392 268443 378448
rect 266524 378390 268443 378392
rect 268377 378387 268443 378390
rect 504725 378450 504791 378453
rect 504725 378448 504834 378450
rect 504725 378392 504730 378448
rect 504786 378392 504834 378448
rect 504725 378387 504834 378392
rect 504774 378148 504834 378387
rect 69841 377906 69907 377909
rect 70301 377906 70367 377909
rect 69841 377904 72036 377906
rect 69841 377848 69846 377904
rect 69902 377848 70306 377904
rect 70362 377848 72036 377904
rect 69841 377846 72036 377848
rect 69841 377843 69907 377846
rect 70301 377843 70367 377846
rect 358077 377770 358143 377773
rect 358077 377768 360180 377770
rect 358077 377712 358082 377768
rect 358138 377712 360180 377768
rect 358077 377710 360180 377712
rect 358077 377707 358143 377710
rect 393313 377226 393379 377229
rect 391092 377224 393379 377226
rect 391092 377168 393318 377224
rect 393374 377168 393379 377224
rect 391092 377166 393379 377168
rect 393313 377163 393379 377166
rect 128905 376954 128971 376957
rect 128678 376952 128971 376954
rect 128678 376896 128910 376952
rect 128966 376896 128971 376952
rect 128678 376894 128971 376896
rect 128678 376818 128738 376894
rect 128905 376891 128971 376894
rect 128813 376818 128879 376821
rect 128678 376816 128879 376818
rect 128678 376760 128818 376816
rect 128874 376760 128879 376816
rect 128678 376758 128879 376760
rect 128813 376755 128879 376758
rect 456793 375186 456859 375189
rect 456793 375184 460092 375186
rect 456793 375128 456798 375184
rect 456854 375128 460092 375184
rect 456793 375126 460092 375128
rect 456793 375123 456859 375126
rect 197905 374370 197971 374373
rect 268469 374370 268535 374373
rect 197905 374368 200100 374370
rect 197905 374312 197910 374368
rect 197966 374312 200100 374368
rect 197905 374310 200100 374312
rect 266524 374368 268535 374370
rect 266524 374312 268474 374368
rect 268530 374312 268535 374368
rect 266524 374310 268535 374312
rect 197905 374307 197971 374310
rect 268469 374307 268535 374310
rect 357433 374234 357499 374237
rect 357433 374232 360180 374234
rect 357433 374176 357438 374232
rect 357494 374176 360180 374232
rect 357433 374174 360180 374176
rect 357433 374171 357499 374174
rect 393405 373962 393471 373965
rect 391092 373960 393471 373962
rect 391092 373904 393410 373960
rect 393466 373904 393471 373960
rect 391092 373902 393471 373904
rect 393405 373899 393471 373902
rect 128445 373282 128511 373285
rect 129181 373282 129247 373285
rect 126132 373280 129247 373282
rect 126132 373224 128450 373280
rect 128506 373224 129186 373280
rect 129242 373224 129247 373280
rect 126132 373222 129247 373224
rect 128445 373219 128511 373222
rect 129181 373219 129247 373222
rect 358077 370970 358143 370973
rect 358077 370968 360180 370970
rect 358077 370912 358082 370968
rect 358138 370912 360180 370968
rect 358077 370910 360180 370912
rect 358077 370907 358143 370910
rect 392025 370426 392091 370429
rect 391092 370424 392091 370426
rect 391092 370368 392030 370424
rect 392086 370368 392091 370424
rect 391092 370366 392091 370368
rect 392025 370363 392091 370366
rect 70209 370290 70275 370293
rect 197813 370290 197879 370293
rect 70209 370288 72036 370290
rect 70209 370232 70214 370288
rect 70270 370232 72036 370288
rect 70209 370230 72036 370232
rect 197813 370288 200100 370290
rect 197813 370232 197818 370288
rect 197874 370232 200100 370288
rect 197813 370230 200100 370232
rect 70209 370227 70275 370230
rect 197813 370227 197879 370230
rect 268561 370018 268627 370021
rect 266524 370016 268627 370018
rect 266524 369960 268566 370016
rect 268622 369960 268627 370016
rect 266524 369958 268627 369960
rect 268561 369955 268627 369958
rect 580717 369610 580783 369613
rect 583520 369610 584960 369700
rect 580717 369608 584960 369610
rect 580717 369552 580722 369608
rect 580778 369552 584960 369608
rect 580717 369550 584960 369552
rect 580717 369547 580783 369550
rect 583520 369460 584960 369550
rect 358169 367434 358235 367437
rect 358169 367432 360180 367434
rect 358169 367376 358174 367432
rect 358230 367376 360180 367432
rect 358169 367374 360180 367376
rect 358169 367371 358235 367374
rect 283966 367236 283972 367300
rect 284036 367298 284042 367300
rect 284036 367238 284218 367298
rect 284036 367236 284042 367238
rect 284158 367165 284218 367238
rect 284109 367160 284218 367165
rect 284109 367104 284114 367160
rect 284170 367104 284218 367160
rect 284109 367102 284218 367104
rect 284109 367099 284175 367102
rect 390694 366893 390754 367132
rect 390645 366888 390754 366893
rect 390645 366832 390650 366888
rect 390706 366832 390754 366888
rect 390645 366830 390754 366832
rect 390645 366827 390711 366830
rect -960 366210 480 366300
rect 2773 366210 2839 366213
rect -960 366208 2839 366210
rect -960 366152 2778 366208
rect 2834 366152 2839 366208
rect -960 366150 2839 366152
rect -960 366060 480 366150
rect 2773 366147 2839 366150
rect 129365 365938 129431 365941
rect 126132 365936 129431 365938
rect 126132 365880 129370 365936
rect 129426 365880 129431 365936
rect 126132 365878 129431 365880
rect 129365 365875 129431 365878
rect 199193 365938 199259 365941
rect 268653 365938 268719 365941
rect 199193 365936 200100 365938
rect 199193 365880 199198 365936
rect 199254 365880 200100 365936
rect 199193 365878 200100 365880
rect 266524 365936 268719 365938
rect 266524 365880 268658 365936
rect 268714 365880 268719 365936
rect 266524 365878 268719 365880
rect 199193 365875 199259 365878
rect 268653 365875 268719 365878
rect 356697 364170 356763 364173
rect 356697 364168 360180 364170
rect 356697 364112 356702 364168
rect 356758 364112 360180 364168
rect 356697 364110 360180 364112
rect 356697 364107 356763 364110
rect 393497 363626 393563 363629
rect 391092 363624 393563 363626
rect 391092 363568 393502 363624
rect 393558 363568 393563 363624
rect 391092 363566 393563 363568
rect 393497 363563 393563 363566
rect 70025 362946 70091 362949
rect 70025 362944 72036 362946
rect 70025 362888 70030 362944
rect 70086 362888 72036 362944
rect 70025 362886 72036 362888
rect 70025 362883 70091 362886
rect 197721 361858 197787 361861
rect 197721 361856 200100 361858
rect 197721 361800 197726 361856
rect 197782 361800 200100 361856
rect 197721 361798 200100 361800
rect 197721 361795 197787 361798
rect 268745 361586 268811 361589
rect 266524 361584 268811 361586
rect 266524 361528 268750 361584
rect 268806 361528 268811 361584
rect 266524 361526 268811 361528
rect 268745 361523 268811 361526
rect 504774 360501 504834 361012
rect 504725 360496 504834 360501
rect 504725 360440 504730 360496
rect 504786 360440 504834 360496
rect 504725 360438 504834 360440
rect 504725 360435 504791 360438
rect 128353 358322 128419 358325
rect 129273 358322 129339 358325
rect 126132 358320 129339 358322
rect 126132 358264 128358 358320
rect 128414 358264 129278 358320
rect 129334 358264 129339 358320
rect 126132 358262 129339 358264
rect 128353 358259 128419 358262
rect 129273 358259 129339 358262
rect 456793 358050 456859 358053
rect 456793 358048 460092 358050
rect 456793 357992 456798 358048
rect 456854 357992 460092 358048
rect 456793 357990 460092 357992
rect 456793 357987 456859 357990
rect 580809 357914 580875 357917
rect 583520 357914 584960 358004
rect 580809 357912 584960 357914
rect 580809 357856 580814 357912
rect 580870 357856 584960 357912
rect 580809 357854 584960 357856
rect 580809 357851 580875 357854
rect 583520 357764 584960 357854
rect 197537 357506 197603 357509
rect 267181 357506 267247 357509
rect 197537 357504 200100 357506
rect 197537 357448 197542 357504
rect 197598 357448 200100 357504
rect 197537 357446 200100 357448
rect 266524 357504 267247 357506
rect 266524 357448 267186 357504
rect 267242 357448 267247 357504
rect 266524 357446 267247 357448
rect 197537 357443 197603 357446
rect 267181 357443 267247 357446
rect 70025 355602 70091 355605
rect 70025 355600 72036 355602
rect 70025 355544 70030 355600
rect 70086 355544 72036 355600
rect 70025 355542 72036 355544
rect 70025 355539 70091 355542
rect 197445 353426 197511 353429
rect 267273 353426 267339 353429
rect 197445 353424 200100 353426
rect 197445 353368 197450 353424
rect 197506 353368 200100 353424
rect 197445 353366 200100 353368
rect 266524 353424 267339 353426
rect 266524 353368 267278 353424
rect 267334 353368 267339 353424
rect 266524 353366 267339 353368
rect 197445 353363 197511 353366
rect 267273 353363 267339 353366
rect -960 351780 480 352020
rect 128997 350978 129063 350981
rect 126132 350976 129063 350978
rect 126132 350920 129002 350976
rect 129058 350920 129063 350976
rect 126132 350918 129063 350920
rect 128997 350915 129063 350918
rect 197353 349074 197419 349077
rect 267641 349074 267707 349077
rect 197353 349072 200100 349074
rect 197353 349016 197358 349072
rect 197414 349016 200100 349072
rect 197353 349014 200100 349016
rect 266524 349072 267707 349074
rect 266524 349016 267646 349072
rect 267702 349016 267707 349072
rect 266524 349014 267707 349016
rect 197353 349011 197419 349014
rect 267641 349011 267707 349014
rect 70117 348258 70183 348261
rect 71497 348258 71563 348261
rect 70117 348256 72036 348258
rect 70117 348200 70122 348256
rect 70178 348200 71502 348256
rect 71558 348200 72036 348256
rect 70117 348198 72036 348200
rect 70117 348195 70183 348198
rect 71497 348195 71563 348198
rect 283925 347986 283991 347989
rect 283925 347984 284218 347986
rect 283925 347928 283930 347984
rect 283986 347928 284218 347984
rect 283925 347926 284218 347928
rect 283925 347923 283991 347926
rect 284158 347853 284218 347926
rect 284109 347848 284218 347853
rect 284109 347792 284114 347848
rect 284170 347792 284218 347848
rect 284109 347790 284218 347792
rect 284109 347787 284175 347790
rect 579981 346082 580047 346085
rect 583520 346082 584960 346172
rect 579981 346080 584960 346082
rect 579981 346024 579986 346080
rect 580042 346024 584960 346080
rect 579981 346022 584960 346024
rect 579981 346019 580047 346022
rect 583520 345932 584960 346022
rect 197629 344994 197695 344997
rect 269021 344994 269087 344997
rect 197629 344992 200100 344994
rect 197629 344936 197634 344992
rect 197690 344936 200100 344992
rect 197629 344934 200100 344936
rect 266524 344992 269087 344994
rect 266524 344936 269026 344992
rect 269082 344936 269087 344992
rect 266524 344934 269087 344936
rect 197629 344931 197695 344934
rect 269021 344931 269087 344934
rect 504774 343637 504834 343876
rect 128813 343634 128879 343637
rect 126132 343632 128879 343634
rect 126132 343576 128818 343632
rect 128874 343576 128879 343632
rect 126132 343574 128879 343576
rect 128813 343571 128879 343574
rect 504725 343632 504834 343637
rect 504725 343576 504730 343632
rect 504786 343576 504834 343632
rect 504725 343574 504834 343576
rect 504725 343571 504791 343574
rect 70025 341458 70091 341461
rect 133965 341458 134031 341461
rect 185577 341458 185643 341461
rect 70025 341456 185643 341458
rect 70025 341400 70030 341456
rect 70086 341400 133970 341456
rect 134026 341400 185582 341456
rect 185638 341400 185643 341456
rect 70025 341398 185643 341400
rect 70025 341395 70091 341398
rect 133965 341395 134031 341398
rect 185577 341395 185643 341398
rect 503713 340914 503779 340917
rect 503897 340914 503963 340917
rect 503713 340912 503963 340914
rect 503713 340856 503718 340912
rect 503774 340856 503902 340912
rect 503958 340856 503963 340912
rect 503713 340854 503963 340856
rect 503713 340851 503779 340854
rect 503897 340851 503963 340854
rect 237189 338738 237255 338741
rect 268142 338738 268148 338740
rect 237189 338736 268148 338738
rect 237189 338680 237194 338736
rect 237250 338680 268148 338736
rect 237189 338678 268148 338680
rect 237189 338675 237255 338678
rect 268142 338676 268148 338678
rect 268212 338676 268218 338740
rect -960 337514 480 337604
rect 2957 337514 3023 337517
rect -960 337512 3023 337514
rect -960 337456 2962 337512
rect 3018 337456 3023 337512
rect -960 337454 3023 337456
rect -960 337364 480 337454
rect 2957 337451 3023 337454
rect 583520 334236 584960 334476
rect -960 323098 480 323188
rect 3969 323098 4035 323101
rect -960 323096 4035 323098
rect -960 323040 3974 323096
rect 4030 323040 4035 323096
rect -960 323038 4035 323040
rect -960 322948 480 323038
rect 3969 323035 4035 323038
rect 579613 322690 579679 322693
rect 583520 322690 584960 322780
rect 579613 322688 584960 322690
rect 579613 322632 579618 322688
rect 579674 322632 584960 322688
rect 579613 322630 584960 322632
rect 579613 322627 579679 322630
rect 583520 322540 584960 322630
rect 390921 318746 390987 318749
rect 391054 318746 391060 318748
rect 390921 318744 391060 318746
rect 390921 318688 390926 318744
rect 390982 318688 391060 318744
rect 390921 318686 391060 318688
rect 390921 318683 390987 318686
rect 391054 318684 391060 318686
rect 391124 318684 391130 318748
rect 257705 317388 257771 317389
rect 257654 317324 257660 317388
rect 257724 317386 257771 317388
rect 257724 317384 257816 317386
rect 257766 317328 257816 317384
rect 257724 317326 257816 317328
rect 257724 317324 257771 317326
rect 257705 317323 257771 317324
rect 257654 311748 257660 311812
rect 257724 311810 257730 311812
rect 257797 311810 257863 311813
rect 257724 311808 257863 311810
rect 257724 311752 257802 311808
rect 257858 311752 257863 311808
rect 257724 311750 257863 311752
rect 257724 311748 257730 311750
rect 257797 311747 257863 311750
rect 579705 310858 579771 310861
rect 583520 310858 584960 310948
rect 579705 310856 584960 310858
rect 579705 310800 579710 310856
rect 579766 310800 584960 310856
rect 579705 310798 584960 310800
rect 579705 310795 579771 310798
rect 583520 310708 584960 310798
rect 390921 309226 390987 309229
rect 391054 309226 391060 309228
rect 390921 309224 391060 309226
rect 390921 309168 390926 309224
rect 390982 309168 391060 309224
rect 390921 309166 391060 309168
rect 390921 309163 390987 309166
rect 391054 309164 391060 309166
rect 391124 309164 391130 309228
rect -960 308818 480 308908
rect 4061 308818 4127 308821
rect -960 308816 4127 308818
rect -960 308760 4066 308816
rect 4122 308760 4127 308816
rect -960 308758 4127 308760
rect -960 308668 480 308758
rect 4061 308755 4127 308758
rect 390921 299434 390987 299437
rect 391054 299434 391060 299436
rect 390921 299432 391060 299434
rect 390921 299376 390926 299432
rect 390982 299376 391060 299432
rect 390921 299374 391060 299376
rect 390921 299371 390987 299374
rect 391054 299372 391060 299374
rect 391124 299372 391130 299436
rect 580625 299162 580691 299165
rect 583520 299162 584960 299252
rect 580625 299160 584960 299162
rect 580625 299104 580630 299160
rect 580686 299104 584960 299160
rect 580625 299102 584960 299104
rect 580625 299099 580691 299102
rect 583520 299012 584960 299102
rect 297633 298074 297699 298077
rect 297766 298074 297772 298076
rect 297633 298072 297772 298074
rect 297633 298016 297638 298072
rect 297694 298016 297772 298072
rect 297633 298014 297772 298016
rect 297633 298011 297699 298014
rect 297766 298012 297772 298014
rect 297836 298012 297842 298076
rect -960 294402 480 294492
rect 3325 294402 3391 294405
rect -960 294400 3391 294402
rect -960 294344 3330 294400
rect 3386 294344 3391 294400
rect -960 294342 3391 294344
rect -960 294252 480 294342
rect 3325 294339 3391 294342
rect 390921 289914 390987 289917
rect 391054 289914 391060 289916
rect 390921 289912 391060 289914
rect 390921 289856 390926 289912
rect 390982 289856 391060 289912
rect 390921 289854 391060 289856
rect 390921 289851 390987 289854
rect 391054 289852 391060 289854
rect 391124 289852 391130 289916
rect 297633 288554 297699 288557
rect 297766 288554 297772 288556
rect 297633 288552 297772 288554
rect 297633 288496 297638 288552
rect 297694 288496 297772 288552
rect 297633 288494 297772 288496
rect 297633 288491 297699 288494
rect 297766 288492 297772 288494
rect 297836 288492 297842 288556
rect 583520 287316 584960 287556
rect -960 280122 480 280212
rect 4061 280122 4127 280125
rect -960 280120 4127 280122
rect -960 280064 4066 280120
rect 4122 280064 4127 280120
rect -960 280062 4127 280064
rect -960 279972 480 280062
rect 4061 280059 4127 280062
rect 390921 280122 390987 280125
rect 391054 280122 391060 280124
rect 390921 280120 391060 280122
rect 390921 280064 390926 280120
rect 390982 280064 391060 280120
rect 390921 280062 391060 280064
rect 390921 280059 390987 280062
rect 391054 280060 391060 280062
rect 391124 280060 391130 280124
rect 579613 275770 579679 275773
rect 583520 275770 584960 275860
rect 579613 275768 584960 275770
rect 579613 275712 579618 275768
rect 579674 275712 584960 275768
rect 579613 275710 584960 275712
rect 579613 275707 579679 275710
rect 583520 275620 584960 275710
rect 390921 270602 390987 270605
rect 391054 270602 391060 270604
rect 390921 270600 391060 270602
rect 390921 270544 390926 270600
rect 390982 270544 391060 270600
rect 390921 270542 391060 270544
rect 390921 270539 390987 270542
rect 391054 270540 391060 270542
rect 391124 270540 391130 270604
rect -960 265706 480 265796
rect 2773 265706 2839 265709
rect -960 265704 2839 265706
rect -960 265648 2778 265704
rect 2834 265648 2839 265704
rect -960 265646 2839 265648
rect -960 265556 480 265646
rect 2773 265643 2839 265646
rect 580165 263938 580231 263941
rect 583520 263938 584960 264028
rect 580165 263936 584960 263938
rect 580165 263880 580170 263936
rect 580226 263880 584960 263936
rect 580165 263878 584960 263880
rect 580165 263875 580231 263878
rect 583520 263788 584960 263878
rect 504265 260946 504331 260949
rect 504633 260946 504699 260949
rect 504265 260944 504699 260946
rect 504265 260888 504270 260944
rect 504326 260888 504638 260944
rect 504694 260888 504699 260944
rect 504265 260886 504699 260888
rect 504265 260883 504331 260886
rect 504633 260883 504699 260886
rect 297357 260810 297423 260813
rect 297541 260810 297607 260813
rect 297357 260808 297607 260810
rect 297357 260752 297362 260808
rect 297418 260752 297546 260808
rect 297602 260752 297607 260808
rect 297357 260750 297607 260752
rect 297357 260747 297423 260750
rect 297541 260747 297607 260750
rect 580717 252242 580783 252245
rect 583520 252242 584960 252332
rect 580717 252240 584960 252242
rect 580717 252184 580722 252240
rect 580778 252184 584960 252240
rect 580717 252182 584960 252184
rect 580717 252179 580783 252182
rect 583520 252092 584960 252182
rect -960 251290 480 251380
rect 3325 251290 3391 251293
rect -960 251288 3391 251290
rect -960 251232 3330 251288
rect 3386 251232 3391 251288
rect -960 251230 3391 251232
rect -960 251140 480 251230
rect 3325 251227 3391 251230
rect 134057 249794 134123 249797
rect 134241 249794 134307 249797
rect 134057 249792 134307 249794
rect 134057 249736 134062 249792
rect 134118 249736 134246 249792
rect 134302 249736 134307 249792
rect 134057 249734 134307 249736
rect 134057 249731 134123 249734
rect 134241 249731 134307 249734
rect 209773 241498 209839 241501
rect 209957 241498 210023 241501
rect 209773 241496 210023 241498
rect 209773 241440 209778 241496
rect 209834 241440 209962 241496
rect 210018 241440 210023 241496
rect 209773 241438 210023 241440
rect 209773 241435 209839 241438
rect 209957 241435 210023 241438
rect 284109 241498 284175 241501
rect 284293 241498 284359 241501
rect 284109 241496 284359 241498
rect 284109 241440 284114 241496
rect 284170 241440 284298 241496
rect 284354 241440 284359 241496
rect 284109 241438 284359 241440
rect 284109 241435 284175 241438
rect 284293 241435 284359 241438
rect 583520 240396 584960 240636
rect 297357 240138 297423 240141
rect 297541 240138 297607 240141
rect 297357 240136 297607 240138
rect 297357 240080 297362 240136
rect 297418 240080 297546 240136
rect 297602 240080 297607 240136
rect 297357 240078 297607 240080
rect 297357 240075 297423 240078
rect 297541 240075 297607 240078
rect -960 237010 480 237100
rect 3325 237010 3391 237013
rect -960 237008 3391 237010
rect -960 236952 3330 237008
rect 3386 236952 3391 237008
rect -960 236950 3391 236952
rect -960 236860 480 236950
rect 3325 236947 3391 236950
rect 580165 228850 580231 228853
rect 583520 228850 584960 228940
rect 580165 228848 584960 228850
rect 580165 228792 580170 228848
rect 580226 228792 584960 228848
rect 580165 228790 584960 228792
rect 580165 228787 580231 228790
rect 583520 228700 584960 228790
rect -960 222594 480 222684
rect 2957 222594 3023 222597
rect -960 222592 3023 222594
rect -960 222536 2962 222592
rect 3018 222536 3023 222592
rect -960 222534 3023 222536
rect -960 222444 480 222534
rect 2957 222531 3023 222534
rect 209773 222186 209839 222189
rect 209957 222186 210023 222189
rect 209773 222184 210023 222186
rect 209773 222128 209778 222184
rect 209834 222128 209962 222184
rect 210018 222128 210023 222184
rect 209773 222126 210023 222128
rect 209773 222123 209839 222126
rect 209957 222123 210023 222126
rect 579613 217018 579679 217021
rect 583520 217018 584960 217108
rect 579613 217016 584960 217018
rect 579613 216960 579618 217016
rect 579674 216960 584960 217016
rect 579613 216958 584960 216960
rect 579613 216955 579679 216958
rect 583520 216868 584960 216958
rect 283649 212530 283715 212533
rect 283925 212530 283991 212533
rect 283649 212528 283991 212530
rect 283649 212472 283654 212528
rect 283710 212472 283930 212528
rect 283986 212472 283991 212528
rect 283649 212470 283991 212472
rect 283649 212467 283715 212470
rect 283925 212467 283991 212470
rect -960 208178 480 208268
rect 2957 208178 3023 208181
rect -960 208176 3023 208178
rect -960 208120 2962 208176
rect 3018 208120 3023 208176
rect -960 208118 3023 208120
rect -960 208028 480 208118
rect 2957 208115 3023 208118
rect 580809 205322 580875 205325
rect 583520 205322 584960 205412
rect 580809 205320 584960 205322
rect 580809 205264 580814 205320
rect 580870 205264 584960 205320
rect 580809 205262 584960 205264
rect 580809 205259 580875 205262
rect 583520 205172 584960 205262
rect 197077 202874 197143 202877
rect 220353 202874 220419 202877
rect 197077 202872 220419 202874
rect 197077 202816 197082 202872
rect 197138 202816 220358 202872
rect 220414 202816 220419 202872
rect 197077 202814 220419 202816
rect 197077 202811 197143 202814
rect 220353 202811 220419 202814
rect 266169 202874 266235 202877
rect 266854 202874 266860 202876
rect 266169 202872 266860 202874
rect 266169 202816 266174 202872
rect 266230 202816 266860 202872
rect 266169 202814 266860 202816
rect 266169 202811 266235 202814
rect 266854 202812 266860 202814
rect 266924 202812 266930 202876
rect 197169 202738 197235 202741
rect 223849 202738 223915 202741
rect 197169 202736 223915 202738
rect 197169 202680 197174 202736
rect 197230 202680 223854 202736
rect 223910 202680 223915 202736
rect 197169 202678 223915 202680
rect 197169 202675 197235 202678
rect 223849 202675 223915 202678
rect 197854 202540 197860 202604
rect 197924 202602 197930 202604
rect 225137 202602 225203 202605
rect 197924 202600 225203 202602
rect 197924 202544 225142 202600
rect 225198 202544 225203 202600
rect 197924 202542 225203 202544
rect 197924 202540 197930 202542
rect 225137 202539 225203 202542
rect 197261 202466 197327 202469
rect 226333 202466 226399 202469
rect 197261 202464 226399 202466
rect 197261 202408 197266 202464
rect 197322 202408 226338 202464
rect 226394 202408 226399 202464
rect 197261 202406 226399 202408
rect 197261 202403 197327 202406
rect 226333 202403 226399 202406
rect 198222 202268 198228 202332
rect 198292 202330 198298 202332
rect 232129 202330 232195 202333
rect 198292 202328 232195 202330
rect 198292 202272 232134 202328
rect 232190 202272 232195 202328
rect 198292 202270 232195 202272
rect 198292 202268 198298 202270
rect 232129 202267 232195 202270
rect 196985 202194 197051 202197
rect 233417 202194 233483 202197
rect 196985 202192 233483 202194
rect 196985 202136 196990 202192
rect 197046 202136 233422 202192
rect 233478 202136 233483 202192
rect 196985 202134 233483 202136
rect 196985 202131 197051 202134
rect 233417 202131 233483 202134
rect 257061 202194 257127 202197
rect 267774 202194 267780 202196
rect 257061 202192 267780 202194
rect 257061 202136 257066 202192
rect 257122 202136 267780 202192
rect 257061 202134 267780 202136
rect 257061 202131 257127 202134
rect 267774 202132 267780 202134
rect 267844 202132 267850 202196
rect 199694 201996 199700 202060
rect 199764 202058 199770 202060
rect 218053 202058 218119 202061
rect 199764 202056 218119 202058
rect 199764 202000 218058 202056
rect 218114 202000 218119 202056
rect 199764 201998 218119 202000
rect 199764 201996 199770 201998
rect 218053 201995 218119 201998
rect 198406 201860 198412 201924
rect 198476 201922 198482 201924
rect 212533 201922 212599 201925
rect 198476 201920 212599 201922
rect 198476 201864 212538 201920
rect 212594 201864 212599 201920
rect 198476 201862 212599 201864
rect 198476 201860 198482 201862
rect 212533 201859 212599 201862
rect 198590 201724 198596 201788
rect 198660 201786 198666 201788
rect 213453 201786 213519 201789
rect 198660 201784 213519 201786
rect 198660 201728 213458 201784
rect 213514 201728 213519 201784
rect 198660 201726 213519 201728
rect 198660 201724 198666 201726
rect 213453 201723 213519 201726
rect 198038 201588 198044 201652
rect 198108 201650 198114 201652
rect 211153 201650 211219 201653
rect 198108 201648 211219 201650
rect 198108 201592 211158 201648
rect 211214 201592 211219 201648
rect 198108 201590 211219 201592
rect 198108 201588 198114 201590
rect 211153 201587 211219 201590
rect 262673 201650 262739 201653
rect 267958 201650 267964 201652
rect 262673 201648 267964 201650
rect 262673 201592 262678 201648
rect 262734 201592 267964 201648
rect 262673 201590 267964 201592
rect 262673 201587 262739 201590
rect 267958 201588 267964 201590
rect 268028 201588 268034 201652
rect 132902 200636 132908 200700
rect 132972 200698 132978 200700
rect 527173 200698 527239 200701
rect 132972 200696 527239 200698
rect 132972 200640 527178 200696
rect 527234 200640 527239 200696
rect 132972 200638 527239 200640
rect 132972 200636 132978 200638
rect 527173 200635 527239 200638
rect 131757 199338 131823 199341
rect 131757 199336 134044 199338
rect 131757 199280 131762 199336
rect 131818 199280 134044 199336
rect 131757 199278 134044 199280
rect 131757 199275 131823 199278
rect 436185 198930 436251 198933
rect 433934 198928 436251 198930
rect 433934 198872 436190 198928
rect 436246 198872 436251 198928
rect 433934 198870 436251 198872
rect 433934 198764 433994 198870
rect 436185 198867 436251 198870
rect 131389 198250 131455 198253
rect 131389 198248 134044 198250
rect 131389 198192 131394 198248
rect 131450 198192 134044 198248
rect 131389 198190 134044 198192
rect 131389 198187 131455 198190
rect 131389 197162 131455 197165
rect 131389 197160 134044 197162
rect 131389 197104 131394 197160
rect 131450 197104 134044 197160
rect 131389 197102 134044 197104
rect 131389 197099 131455 197102
rect 130837 196210 130903 196213
rect 433934 196210 433994 196724
rect 434989 196210 435055 196213
rect 130837 196208 134044 196210
rect 130837 196152 130842 196208
rect 130898 196152 134044 196208
rect 130837 196150 134044 196152
rect 433934 196208 435055 196210
rect 433934 196152 434994 196208
rect 435050 196152 435055 196208
rect 433934 196150 435055 196152
rect 130837 196147 130903 196150
rect 434989 196147 435055 196150
rect 130837 194714 130903 194717
rect 134014 194714 134074 195092
rect 130837 194712 134074 194714
rect 130837 194656 130842 194712
rect 130898 194656 134074 194712
rect 130837 194654 134074 194656
rect 130837 194651 130903 194654
rect 130837 194442 130903 194445
rect 130837 194440 134074 194442
rect 130837 194384 130842 194440
rect 130898 194384 134074 194440
rect 130837 194382 134074 194384
rect 130837 194379 130903 194382
rect 134014 194004 134074 194382
rect 433934 194034 433994 194548
rect 436277 194034 436343 194037
rect 433934 194032 436343 194034
rect -960 193898 480 193988
rect 433934 193976 436282 194032
rect 436338 193976 436343 194032
rect 433934 193974 436343 193976
rect 436277 193971 436343 193974
rect 3601 193898 3667 193901
rect -960 193896 3667 193898
rect -960 193840 3606 193896
rect 3662 193840 3667 193896
rect -960 193838 3667 193840
rect -960 193748 480 193838
rect 3601 193835 3667 193838
rect 583520 193476 584960 193716
rect 130837 193082 130903 193085
rect 436645 193082 436711 193085
rect 130837 193080 134074 193082
rect 130837 193024 130842 193080
rect 130898 193024 134074 193080
rect 130837 193022 134074 193024
rect 130837 193019 130903 193022
rect 134014 192916 134074 193022
rect 433934 193080 436711 193082
rect 433934 193024 436650 193080
rect 436706 193024 436711 193080
rect 433934 193022 436711 193024
rect 130745 192538 130811 192541
rect 130745 192536 134074 192538
rect 130745 192480 130750 192536
rect 130806 192480 134074 192536
rect 433934 192508 433994 193022
rect 436645 193019 436711 193022
rect 130745 192478 134074 192480
rect 130745 192475 130811 192478
rect 134014 191964 134074 192478
rect 130837 191450 130903 191453
rect 130837 191448 134074 191450
rect 130837 191392 130842 191448
rect 130898 191392 134074 191448
rect 130837 191390 134074 191392
rect 130837 191387 130903 191390
rect 134014 190876 134074 191390
rect 130837 190362 130903 190365
rect 130837 190360 134074 190362
rect 130837 190304 130842 190360
rect 130898 190304 134074 190360
rect 130837 190302 134074 190304
rect 130837 190299 130903 190302
rect 134014 189788 134074 190302
rect 433934 190226 433994 190332
rect 435173 190226 435239 190229
rect 433934 190224 435239 190226
rect 433934 190168 435178 190224
rect 435234 190168 435239 190224
rect 433934 190166 435239 190168
rect 435173 190163 435239 190166
rect 130837 189002 130903 189005
rect 130837 189000 134074 189002
rect 130837 188944 130842 189000
rect 130898 188944 134074 189000
rect 130837 188942 134074 188944
rect 130837 188939 130903 188942
rect 134014 188700 134074 188942
rect 435081 188866 435147 188869
rect 433934 188864 435147 188866
rect 433934 188808 435086 188864
rect 435142 188808 435147 188864
rect 433934 188806 435147 188808
rect 130745 188322 130811 188325
rect 130745 188320 134074 188322
rect 130745 188264 130750 188320
rect 130806 188264 134074 188320
rect 433934 188292 433994 188806
rect 435081 188803 435147 188806
rect 130745 188262 134074 188264
rect 130745 188259 130811 188262
rect 134014 187748 134074 188262
rect 130837 187234 130903 187237
rect 130837 187232 134074 187234
rect 130837 187176 130842 187232
rect 130898 187176 134074 187232
rect 130837 187174 134074 187176
rect 130837 187171 130903 187174
rect 134014 186660 134074 187174
rect 434529 186282 434595 186285
rect 433934 186280 434595 186282
rect 433934 186224 434534 186280
rect 434590 186224 434595 186280
rect 433934 186222 434595 186224
rect 433934 186116 433994 186222
rect 434529 186219 434595 186222
rect 131205 185602 131271 185605
rect 131205 185600 134044 185602
rect 131205 185544 131210 185600
rect 131266 185544 134044 185600
rect 131205 185542 134044 185544
rect 131205 185539 131271 185542
rect 434897 184650 434963 184653
rect 433934 184648 434963 184650
rect 433934 184592 434902 184648
rect 434958 184592 434963 184648
rect 433934 184590 434963 184592
rect 131205 184514 131271 184517
rect 131205 184512 134044 184514
rect 131205 184456 131210 184512
rect 131266 184456 134044 184512
rect 131205 184454 134044 184456
rect 131205 184451 131271 184454
rect 433934 184076 433994 184590
rect 434897 184587 434963 184590
rect 131205 183562 131271 183565
rect 504357 183562 504423 183565
rect 504633 183562 504699 183565
rect 131205 183560 134044 183562
rect 131205 183504 131210 183560
rect 131266 183504 134044 183560
rect 131205 183502 134044 183504
rect 504357 183560 504699 183562
rect 504357 183504 504362 183560
rect 504418 183504 504638 183560
rect 504694 183504 504699 183560
rect 504357 183502 504699 183504
rect 131205 183499 131271 183502
rect 504357 183499 504423 183502
rect 504633 183499 504699 183502
rect 133321 182474 133387 182477
rect 133321 182472 134044 182474
rect 133321 182416 133326 182472
rect 133382 182416 134044 182472
rect 133321 182414 134044 182416
rect 133321 182411 133387 182414
rect 128813 182202 128879 182205
rect 128997 182202 129063 182205
rect 128813 182200 129063 182202
rect 128813 182144 128818 182200
rect 128874 182144 129002 182200
rect 129058 182144 129063 182200
rect 128813 182142 129063 182144
rect 128813 182139 128879 182142
rect 128997 182139 129063 182142
rect 436553 182066 436619 182069
rect 433934 182064 436619 182066
rect 433934 182008 436558 182064
rect 436614 182008 436619 182064
rect 433934 182006 436619 182008
rect 433934 181900 433994 182006
rect 436553 182003 436619 182006
rect 580257 181930 580323 181933
rect 583520 181930 584960 182020
rect 580257 181928 584960 181930
rect 580257 181872 580262 181928
rect 580318 181872 584960 181928
rect 580257 181870 584960 181872
rect 580257 181867 580323 181870
rect 583520 181780 584960 181870
rect 133413 181386 133479 181389
rect 133413 181384 134044 181386
rect 133413 181328 133418 181384
rect 133474 181328 134044 181384
rect 133413 181326 134044 181328
rect 133413 181323 133479 181326
rect 133873 180434 133939 180437
rect 133873 180432 134044 180434
rect 133873 180376 133878 180432
rect 133934 180376 134044 180432
rect 133873 180374 134044 180376
rect 133873 180371 133939 180374
rect 436093 180298 436159 180301
rect 433934 180296 436159 180298
rect 433934 180240 436098 180296
rect 436154 180240 436159 180296
rect 433934 180238 436159 180240
rect 433934 179860 433994 180238
rect 436093 180235 436159 180238
rect -960 179482 480 179572
rect 2865 179482 2931 179485
rect -960 179480 2931 179482
rect -960 179424 2870 179480
rect 2926 179424 2931 179480
rect -960 179422 2931 179424
rect -960 179332 480 179422
rect 2865 179419 2931 179422
rect 132493 179346 132559 179349
rect 132493 179344 134044 179346
rect 132493 179288 132498 179344
rect 132554 179288 134044 179344
rect 132493 179286 134044 179288
rect 132493 179283 132559 179286
rect 131205 178258 131271 178261
rect 131205 178256 134044 178258
rect 131205 178200 131210 178256
rect 131266 178200 134044 178256
rect 131205 178198 134044 178200
rect 131205 178195 131271 178198
rect 436461 177986 436527 177989
rect 433934 177984 436527 177986
rect 433934 177928 436466 177984
rect 436522 177928 436527 177984
rect 433934 177926 436527 177928
rect 433934 177684 433994 177926
rect 436461 177923 436527 177926
rect 132585 177170 132651 177173
rect 132585 177168 134044 177170
rect 132585 177112 132590 177168
rect 132646 177112 134044 177168
rect 132585 177110 134044 177112
rect 132585 177107 132651 177110
rect 132902 176156 132908 176220
rect 132972 176218 132978 176220
rect 436369 176218 436435 176221
rect 132972 176158 134044 176218
rect 433934 176216 436435 176218
rect 433934 176160 436374 176216
rect 436430 176160 436435 176216
rect 433934 176158 436435 176160
rect 132972 176156 132978 176158
rect 433934 175644 433994 176158
rect 436369 176155 436435 176158
rect 133638 175068 133644 175132
rect 133708 175130 133714 175132
rect 133708 175070 134044 175130
rect 133708 175068 133714 175070
rect 133454 173980 133460 174044
rect 133524 174042 133530 174044
rect 133524 173982 134044 174042
rect 133524 173980 133530 173982
rect 434805 173906 434871 173909
rect 433934 173904 434871 173906
rect 433934 173848 434810 173904
rect 434866 173848 434871 173904
rect 433934 173846 434871 173848
rect 433934 173468 433994 173846
rect 434805 173843 434871 173846
rect 133086 172892 133092 172956
rect 133156 172954 133162 172956
rect 133156 172894 134044 172954
rect 133156 172892 133162 172894
rect 132401 172002 132467 172005
rect 434713 172002 434779 172005
rect 132401 172000 134044 172002
rect 132401 171944 132406 172000
rect 132462 171944 134044 172000
rect 132401 171942 134044 171944
rect 433934 172000 434779 172002
rect 433934 171944 434718 172000
rect 434774 171944 434779 172000
rect 433934 171942 434779 171944
rect 132401 171939 132467 171942
rect 433934 171428 433994 171942
rect 434713 171939 434779 171942
rect 132217 170914 132283 170917
rect 132217 170912 134044 170914
rect 132217 170856 132222 170912
rect 132278 170856 134044 170912
rect 132217 170854 134044 170856
rect 132217 170851 132283 170854
rect 580257 170098 580323 170101
rect 583520 170098 584960 170188
rect 580257 170096 584960 170098
rect 580257 170040 580262 170096
rect 580318 170040 584960 170096
rect 580257 170038 584960 170040
rect 580257 170035 580323 170038
rect 583520 169948 584960 170038
rect 133137 169826 133203 169829
rect 133137 169824 134044 169826
rect 133137 169768 133142 169824
rect 133198 169768 134044 169824
rect 133137 169766 134044 169768
rect 133137 169763 133203 169766
rect 434253 169690 434319 169693
rect 433934 169688 434319 169690
rect 433934 169632 434258 169688
rect 434314 169632 434319 169688
rect 433934 169630 434319 169632
rect 433934 169252 433994 169630
rect 434253 169627 434319 169630
rect 133045 168738 133111 168741
rect 133045 168736 134044 168738
rect 133045 168680 133050 168736
rect 133106 168680 134044 168736
rect 133045 168678 134044 168680
rect 133045 168675 133111 168678
rect 131665 167786 131731 167789
rect 434437 167786 434503 167789
rect 131665 167784 134044 167786
rect 131665 167728 131670 167784
rect 131726 167728 134044 167784
rect 131665 167726 134044 167728
rect 433934 167784 434503 167786
rect 433934 167728 434442 167784
rect 434498 167728 434503 167784
rect 433934 167726 434503 167728
rect 131665 167723 131731 167726
rect 433934 167212 433994 167726
rect 434437 167723 434503 167726
rect 132769 166698 132835 166701
rect 132769 166696 134044 166698
rect 132769 166640 132774 166696
rect 132830 166640 134044 166696
rect 132769 166638 134044 166640
rect 132769 166635 132835 166638
rect 132677 165610 132743 165613
rect 434345 165610 434411 165613
rect 132677 165608 134044 165610
rect 132677 165552 132682 165608
rect 132738 165552 134044 165608
rect 132677 165550 134044 165552
rect 433934 165608 434411 165610
rect 433934 165552 434350 165608
rect 434406 165552 434411 165608
rect 433934 165550 434411 165552
rect 132677 165547 132743 165550
rect -960 165066 480 165156
rect 3233 165066 3299 165069
rect -960 165064 3299 165066
rect -960 165008 3238 165064
rect 3294 165008 3299 165064
rect 433934 165036 433994 165550
rect 434345 165547 434411 165550
rect -960 165006 3299 165008
rect -960 164916 480 165006
rect 3233 165003 3299 165006
rect 131297 164522 131363 164525
rect 131297 164520 134044 164522
rect 131297 164464 131302 164520
rect 131358 164464 134044 164520
rect 131297 164462 134044 164464
rect 131297 164459 131363 164462
rect 133597 163570 133663 163573
rect 434161 163570 434227 163573
rect 133597 163568 134044 163570
rect 133597 163512 133602 163568
rect 133658 163512 134044 163568
rect 133597 163510 134044 163512
rect 433934 163568 434227 163570
rect 433934 163512 434166 163568
rect 434222 163512 434227 163568
rect 433934 163510 434227 163512
rect 133597 163507 133663 163510
rect 433934 162996 433994 163510
rect 434161 163507 434227 163510
rect 132401 162482 132467 162485
rect 132401 162480 134044 162482
rect 132401 162424 132406 162480
rect 132462 162424 134044 162480
rect 132401 162422 134044 162424
rect 132401 162419 132467 162422
rect 132677 161394 132743 161397
rect 132677 161392 134044 161394
rect 132677 161336 132682 161392
rect 132738 161336 134044 161392
rect 132677 161334 134044 161336
rect 132677 161331 132743 161334
rect 434069 161258 434135 161261
rect 433934 161256 434135 161258
rect 433934 161200 434074 161256
rect 434130 161200 434135 161256
rect 433934 161198 434135 161200
rect 433934 160956 433994 161198
rect 434069 161195 434135 161198
rect 133597 160442 133663 160445
rect 133597 160440 134044 160442
rect 133597 160384 133602 160440
rect 133658 160384 134044 160440
rect 133597 160382 134044 160384
rect 133597 160379 133663 160382
rect 132217 159354 132283 159357
rect 433977 159354 434043 159357
rect 132217 159352 134044 159354
rect 132217 159296 132222 159352
rect 132278 159296 134044 159352
rect 132217 159294 134044 159296
rect 433934 159352 434043 159354
rect 433934 159296 433982 159352
rect 434038 159296 434043 159352
rect 132217 159291 132283 159294
rect 433934 159291 434043 159296
rect 433934 158780 433994 159291
rect 580165 158402 580231 158405
rect 583520 158402 584960 158492
rect 580165 158400 584960 158402
rect 580165 158344 580170 158400
rect 580226 158344 584960 158400
rect 580165 158342 584960 158344
rect 580165 158339 580231 158342
rect 131665 158266 131731 158269
rect 131665 158264 134044 158266
rect 131665 158208 131670 158264
rect 131726 158208 134044 158264
rect 583520 158252 584960 158342
rect 131665 158206 134044 158208
rect 131665 158203 131731 158206
rect 433885 157314 433951 157317
rect 433885 157312 433994 157314
rect 433885 157256 433890 157312
rect 433946 157256 433994 157312
rect 433885 157251 433994 157256
rect 131297 157178 131363 157181
rect 131297 157176 134044 157178
rect 131297 157120 131302 157176
rect 131358 157120 134044 157176
rect 131297 157118 134044 157120
rect 131297 157115 131363 157118
rect 433934 156740 433994 157251
rect 131113 156226 131179 156229
rect 131113 156224 134044 156226
rect 131113 156168 131118 156224
rect 131174 156168 134044 156224
rect 131113 156166 134044 156168
rect 131113 156163 131179 156166
rect 131113 155138 131179 155141
rect 436093 155138 436159 155141
rect 131113 155136 134044 155138
rect 131113 155080 131118 155136
rect 131174 155080 134044 155136
rect 131113 155078 134044 155080
rect 433934 155136 436159 155138
rect 433934 155080 436098 155136
rect 436154 155080 436159 155136
rect 433934 155078 436159 155080
rect 131113 155075 131179 155078
rect 433934 154564 433994 155078
rect 436093 155075 436159 155078
rect 504173 154594 504239 154597
rect 504449 154594 504515 154597
rect 504173 154592 504515 154594
rect 504173 154536 504178 154592
rect 504234 154536 504454 154592
rect 504510 154536 504515 154592
rect 504173 154534 504515 154536
rect 504173 154531 504239 154534
rect 504449 154531 504515 154534
rect 131113 154050 131179 154053
rect 131113 154048 134044 154050
rect 131113 153992 131118 154048
rect 131174 153992 134044 154048
rect 131113 153990 134044 153992
rect 131113 153987 131179 153990
rect 128905 153370 128971 153373
rect 128862 153368 128971 153370
rect 128862 153312 128910 153368
rect 128966 153312 128971 153368
rect 128862 153307 128971 153312
rect 128862 153237 128922 153307
rect 128813 153232 128922 153237
rect 128813 153176 128818 153232
rect 128874 153176 128922 153232
rect 128813 153174 128922 153176
rect 128813 153171 128879 153174
rect 131113 152962 131179 152965
rect 131113 152960 134044 152962
rect 131113 152904 131118 152960
rect 131174 152904 134044 152960
rect 131113 152902 134044 152904
rect 131113 152899 131179 152902
rect 437381 152826 437447 152829
rect 433934 152824 437447 152826
rect 433934 152768 437386 152824
rect 437442 152768 437447 152824
rect 433934 152766 437447 152768
rect 433934 152524 433994 152766
rect 437381 152763 437447 152766
rect 131297 152010 131363 152013
rect 131297 152008 134044 152010
rect 131297 151952 131302 152008
rect 131358 151952 134044 152008
rect 131297 151950 134044 151952
rect 131297 151947 131363 151950
rect 131113 150922 131179 150925
rect 131113 150920 134044 150922
rect -960 150786 480 150876
rect 131113 150864 131118 150920
rect 131174 150864 134044 150920
rect 131113 150862 134044 150864
rect 131113 150859 131179 150862
rect 3233 150786 3299 150789
rect -960 150784 3299 150786
rect -960 150728 3238 150784
rect 3294 150728 3299 150784
rect -960 150726 3299 150728
rect -960 150636 480 150726
rect 3233 150723 3299 150726
rect 433934 150242 433994 150348
rect 437381 150242 437447 150245
rect 433934 150240 437447 150242
rect 433934 150184 437386 150240
rect 437442 150184 437447 150240
rect 433934 150182 437447 150184
rect 437381 150179 437447 150182
rect 131113 149834 131179 149837
rect 131113 149832 134044 149834
rect 131113 149776 131118 149832
rect 131174 149776 134044 149832
rect 131113 149774 134044 149776
rect 131113 149771 131179 149774
rect 131113 148746 131179 148749
rect 436093 148746 436159 148749
rect 131113 148744 134044 148746
rect 131113 148688 131118 148744
rect 131174 148688 134044 148744
rect 131113 148686 134044 148688
rect 433934 148744 436159 148746
rect 433934 148688 436098 148744
rect 436154 148688 436159 148744
rect 433934 148686 436159 148688
rect 131113 148683 131179 148686
rect 433934 148308 433994 148686
rect 436093 148683 436159 148686
rect 131113 147794 131179 147797
rect 131113 147792 134044 147794
rect 131113 147736 131118 147792
rect 131174 147736 134044 147792
rect 131113 147734 134044 147736
rect 131113 147731 131179 147734
rect 131205 146706 131271 146709
rect 131205 146704 134044 146706
rect 131205 146648 131210 146704
rect 131266 146648 134044 146704
rect 131205 146646 134044 146648
rect 131205 146643 131271 146646
rect 583520 146556 584960 146796
rect 437381 146298 437447 146301
rect 433934 146296 437447 146298
rect 433934 146240 437386 146296
rect 437442 146240 437447 146296
rect 433934 146238 437447 146240
rect 433934 146132 433994 146238
rect 437381 146235 437447 146238
rect 131113 145618 131179 145621
rect 131113 145616 134044 145618
rect 131113 145560 131118 145616
rect 131174 145560 134044 145616
rect 131113 145558 134044 145560
rect 131113 145555 131179 145558
rect 128169 144530 128235 144533
rect 437013 144530 437079 144533
rect 128169 144528 134044 144530
rect 128169 144472 128174 144528
rect 128230 144472 134044 144528
rect 128169 144470 134044 144472
rect 433934 144528 437079 144530
rect 433934 144472 437018 144528
rect 437074 144472 437079 144528
rect 433934 144470 437079 144472
rect 128169 144467 128235 144470
rect 433934 144092 433994 144470
rect 437013 144467 437079 144470
rect 131113 143578 131179 143581
rect 131113 143576 134044 143578
rect 131113 143520 131118 143576
rect 131174 143520 134044 143576
rect 131113 143518 134044 143520
rect 131113 143515 131179 143518
rect 133505 142490 133571 142493
rect 133505 142488 134044 142490
rect 133505 142432 133510 142488
rect 133566 142432 134044 142488
rect 133505 142430 134044 142432
rect 133505 142427 133571 142430
rect 436093 142082 436159 142085
rect 433934 142080 436159 142082
rect 433934 142024 436098 142080
rect 436154 142024 436159 142080
rect 433934 142022 436159 142024
rect 433934 141916 433994 142022
rect 436093 142019 436159 142022
rect 133689 141402 133755 141405
rect 133689 141400 134044 141402
rect 133689 141344 133694 141400
rect 133750 141344 134044 141400
rect 133689 141342 134044 141344
rect 133689 141339 133755 141342
rect 133781 140450 133847 140453
rect 436737 140450 436803 140453
rect 133781 140448 134044 140450
rect 133781 140392 133786 140448
rect 133842 140392 134044 140448
rect 133781 140390 134044 140392
rect 433934 140448 436803 140450
rect 433934 140392 436742 140448
rect 436798 140392 436803 140448
rect 433934 140390 436803 140392
rect 133781 140387 133847 140390
rect 433934 139876 433994 140390
rect 436737 140387 436803 140390
rect 131297 139362 131363 139365
rect 131297 139360 134044 139362
rect 131297 139304 131302 139360
rect 131358 139304 134044 139360
rect 131297 139302 134044 139304
rect 131297 139299 131363 139302
rect 132309 138274 132375 138277
rect 132309 138272 134044 138274
rect 132309 138216 132314 138272
rect 132370 138216 134044 138272
rect 132309 138214 134044 138216
rect 132309 138211 132375 138214
rect 437381 137866 437447 137869
rect 433934 137864 437447 137866
rect 433934 137808 437386 137864
rect 437442 137808 437447 137864
rect 433934 137806 437447 137808
rect 433934 137700 433994 137806
rect 437381 137803 437447 137806
rect 132166 137124 132172 137188
rect 132236 137186 132242 137188
rect 132236 137126 134044 137186
rect 132236 137124 132242 137126
rect -960 136370 480 136460
rect 3325 136370 3391 136373
rect -960 136368 3391 136370
rect -960 136312 3330 136368
rect 3386 136312 3391 136368
rect -960 136310 3391 136312
rect -960 136220 480 136310
rect 3325 136307 3391 136310
rect 132350 136172 132356 136236
rect 132420 136234 132426 136236
rect 132420 136174 134044 136234
rect 132420 136172 132426 136174
rect 437013 136098 437079 136101
rect 433934 136096 437079 136098
rect 433934 136040 437018 136096
rect 437074 136040 437079 136096
rect 433934 136038 437079 136040
rect 433934 135660 433994 136038
rect 437013 136035 437079 136038
rect 128905 135418 128971 135421
rect 128862 135416 128971 135418
rect 128862 135360 128910 135416
rect 128966 135360 128971 135416
rect 128862 135355 128971 135360
rect 128862 135285 128922 135355
rect 128813 135280 128922 135285
rect 128813 135224 128818 135280
rect 128874 135224 128922 135280
rect 128813 135222 128922 135224
rect 128813 135219 128879 135222
rect 131982 135084 131988 135148
rect 132052 135146 132058 135148
rect 132052 135086 134044 135146
rect 132052 135084 132058 135086
rect 580349 134874 580415 134877
rect 583520 134874 584960 134964
rect 580349 134872 584960 134874
rect 580349 134816 580354 134872
rect 580410 134816 584960 134872
rect 580349 134814 584960 134816
rect 580349 134811 580415 134814
rect 583520 134724 584960 134814
rect 131798 133996 131804 134060
rect 131868 134058 131874 134060
rect 131868 133998 134044 134058
rect 131868 133996 131874 133998
rect 437381 133650 437447 133653
rect 433934 133648 437447 133650
rect 433934 133592 437386 133648
rect 437442 133592 437447 133648
rect 433934 133590 437447 133592
rect 433934 133484 433994 133590
rect 437381 133587 437447 133590
rect 133270 132908 133276 132972
rect 133340 132970 133346 132972
rect 133340 132910 134044 132970
rect 133340 132908 133346 132910
rect 131389 132018 131455 132021
rect 437381 132018 437447 132021
rect 131389 132016 134044 132018
rect 131389 131960 131394 132016
rect 131450 131960 134044 132016
rect 131389 131958 134044 131960
rect 433934 132016 437447 132018
rect 433934 131960 437386 132016
rect 437442 131960 437447 132016
rect 433934 131958 437447 131960
rect 131389 131955 131455 131958
rect 433934 131444 433994 131958
rect 437381 131955 437447 131958
rect 132125 130930 132191 130933
rect 132125 130928 134044 130930
rect 132125 130872 132130 130928
rect 132186 130872 134044 130928
rect 132125 130870 134044 130872
rect 132125 130867 132191 130870
rect 133229 129842 133295 129845
rect 133229 129840 134044 129842
rect 133229 129784 133234 129840
rect 133290 129784 134044 129840
rect 133229 129782 134044 129784
rect 133229 129779 133295 129782
rect 437381 129570 437447 129573
rect 433934 129568 437447 129570
rect 433934 129512 437386 129568
rect 437442 129512 437447 129568
rect 433934 129510 437447 129512
rect 433934 129268 433994 129510
rect 437381 129507 437447 129510
rect 131941 128754 132007 128757
rect 131941 128752 134044 128754
rect 131941 128696 131946 128752
rect 132002 128696 134044 128752
rect 131941 128694 134044 128696
rect 131941 128691 132007 128694
rect 132033 127802 132099 127805
rect 436829 127802 436895 127805
rect 132033 127800 134044 127802
rect 132033 127744 132038 127800
rect 132094 127744 134044 127800
rect 132033 127742 134044 127744
rect 433934 127800 436895 127802
rect 433934 127744 436834 127800
rect 436890 127744 436895 127800
rect 433934 127742 436895 127744
rect 132033 127739 132099 127742
rect 433934 127228 433994 127742
rect 436829 127739 436895 127742
rect 131849 126714 131915 126717
rect 131849 126712 134044 126714
rect 131849 126656 131854 126712
rect 131910 126656 134044 126712
rect 131849 126654 134044 126656
rect 131849 126651 131915 126654
rect 131573 125626 131639 125629
rect 131573 125624 134044 125626
rect 131573 125568 131578 125624
rect 131634 125568 134044 125624
rect 131573 125566 134044 125568
rect 131573 125563 131639 125566
rect 131481 124538 131547 124541
rect 433934 124538 433994 125052
rect 436921 124538 436987 124541
rect 131481 124536 134044 124538
rect 131481 124480 131486 124536
rect 131542 124480 134044 124536
rect 131481 124478 134044 124480
rect 433934 124536 436987 124538
rect 433934 124480 436926 124536
rect 436982 124480 436987 124536
rect 433934 124478 436987 124480
rect 131481 124475 131547 124478
rect 436921 124475 436987 124478
rect 134014 123045 134074 123556
rect 580533 123178 580599 123181
rect 583520 123178 584960 123268
rect 580533 123176 584960 123178
rect 580533 123120 580538 123176
rect 580594 123120 584960 123176
rect 580533 123118 584960 123120
rect 580533 123115 580599 123118
rect 133965 123040 134074 123045
rect 133965 122984 133970 123040
rect 134026 122984 134074 123040
rect 583520 123028 584960 123118
rect 133965 122982 134074 122984
rect 133965 122979 134031 122982
rect 433934 122906 433994 123012
rect 436829 122906 436895 122909
rect 433934 122904 436895 122906
rect 433934 122848 436834 122904
rect 436890 122848 436895 122904
rect 433934 122846 436895 122848
rect 436829 122843 436895 122846
rect -960 122090 480 122180
rect 3049 122090 3115 122093
rect -960 122088 3115 122090
rect -960 122032 3054 122088
rect 3110 122032 3115 122088
rect -960 122030 3115 122032
rect -960 121940 480 122030
rect 3049 122027 3115 122030
rect 133873 121954 133939 121957
rect 134014 121954 134074 122468
rect 133873 121952 134074 121954
rect 133873 121896 133878 121952
rect 133934 121896 134074 121952
rect 133873 121894 134074 121896
rect 133873 121891 133939 121894
rect 132125 121410 132191 121413
rect 132125 121408 134044 121410
rect 132125 121352 132130 121408
rect 132186 121352 134044 121408
rect 132125 121350 134044 121352
rect 132125 121347 132191 121350
rect 132401 120458 132467 120461
rect 433934 120458 433994 120972
rect 436737 120458 436803 120461
rect 132401 120456 134044 120458
rect 132401 120400 132406 120456
rect 132462 120400 134044 120456
rect 132401 120398 134044 120400
rect 433934 120456 436803 120458
rect 433934 120400 436742 120456
rect 436798 120400 436803 120456
rect 433934 120398 436803 120400
rect 132401 120395 132467 120398
rect 436737 120395 436803 120398
rect 128813 118690 128879 118693
rect 140773 118690 140839 118693
rect 128813 118688 140839 118690
rect 128813 118632 128818 118688
rect 128874 118632 140778 118688
rect 140834 118632 140839 118688
rect 128813 118630 140839 118632
rect 128813 118627 128879 118630
rect 140773 118627 140839 118630
rect 142797 118690 142863 118693
rect 157241 118690 157307 118693
rect 142797 118688 157307 118690
rect 142797 118632 142802 118688
rect 142858 118632 157246 118688
rect 157302 118632 157307 118688
rect 142797 118630 157307 118632
rect 142797 118627 142863 118630
rect 157241 118627 157307 118630
rect 75913 118554 75979 118557
rect 85389 118554 85455 118557
rect 75913 118552 85455 118554
rect 75913 118496 75918 118552
rect 75974 118496 85394 118552
rect 85450 118496 85455 118552
rect 75913 118494 85455 118496
rect 75913 118491 75979 118494
rect 85389 118491 85455 118494
rect 103421 118554 103487 118557
rect 186589 118554 186655 118557
rect 103421 118552 186655 118554
rect 103421 118496 103426 118552
rect 103482 118496 186594 118552
rect 186650 118496 186655 118552
rect 103421 118494 186655 118496
rect 103421 118491 103487 118494
rect 186589 118491 186655 118494
rect 117221 118418 117287 118421
rect 193949 118418 194015 118421
rect 117221 118416 194015 118418
rect 117221 118360 117226 118416
rect 117282 118360 193954 118416
rect 194010 118360 194015 118416
rect 117221 118358 194015 118360
rect 117221 118355 117287 118358
rect 193949 118355 194015 118358
rect 125777 118282 125843 118285
rect 197629 118282 197695 118285
rect 125777 118280 197695 118282
rect 125777 118224 125782 118280
rect 125838 118224 197634 118280
rect 197690 118224 197695 118280
rect 125777 118222 197695 118224
rect 125777 118219 125843 118222
rect 197629 118219 197695 118222
rect 133873 118146 133939 118149
rect 142797 118146 142863 118149
rect 133873 118144 142863 118146
rect 133873 118088 133878 118144
rect 133934 118088 142802 118144
rect 142858 118088 142863 118144
rect 133873 118086 142863 118088
rect 133873 118083 133939 118086
rect 142797 118083 142863 118086
rect 157241 118146 157307 118149
rect 188429 118146 188495 118149
rect 157241 118144 188495 118146
rect 157241 118088 157246 118144
rect 157302 118088 188434 118144
rect 188490 118088 188495 118144
rect 157241 118086 188495 118088
rect 157241 118083 157307 118086
rect 188429 118083 188495 118086
rect 248965 118146 249031 118149
rect 251541 118146 251607 118149
rect 248965 118144 251607 118146
rect 248965 118088 248970 118144
rect 249026 118088 251546 118144
rect 251602 118088 251607 118144
rect 248965 118086 251607 118088
rect 248965 118083 249031 118086
rect 251541 118083 251607 118086
rect 71589 118010 71655 118013
rect 76005 118010 76071 118013
rect 153469 118010 153535 118013
rect 71589 118008 153535 118010
rect 71589 117952 71594 118008
rect 71650 117952 76010 118008
rect 76066 117952 153474 118008
rect 153530 117952 153535 118008
rect 71589 117950 153535 117952
rect 71589 117947 71655 117950
rect 76005 117947 76071 117950
rect 153469 117947 153535 117950
rect 231117 118010 231183 118013
rect 240225 118010 240291 118013
rect 231117 118008 240291 118010
rect 231117 117952 231122 118008
rect 231178 117952 240230 118008
rect 240286 117952 240291 118008
rect 231117 117950 240291 117952
rect 231117 117947 231183 117950
rect 240225 117947 240291 117950
rect 433977 118010 434043 118013
rect 442257 118010 442323 118013
rect 433977 118008 442323 118010
rect 433977 117952 433982 118008
rect 434038 117952 442262 118008
rect 442318 117952 442323 118008
rect 433977 117950 442323 117952
rect 433977 117947 434043 117950
rect 442257 117947 442323 117950
rect 110321 117874 110387 117877
rect 145557 117874 145623 117877
rect 110321 117872 145623 117874
rect 110321 117816 110326 117872
rect 110382 117816 145562 117872
rect 145618 117816 145623 117872
rect 110321 117814 145623 117816
rect 110321 117811 110387 117814
rect 145557 117811 145623 117814
rect 127617 117738 127683 117741
rect 128261 117738 128327 117741
rect 151813 117738 151879 117741
rect 127617 117736 151879 117738
rect 127617 117680 127622 117736
rect 127678 117680 128266 117736
rect 128322 117680 151818 117736
rect 151874 117680 151879 117736
rect 127617 117678 151879 117680
rect 127617 117675 127683 117678
rect 128261 117675 128327 117678
rect 151813 117675 151879 117678
rect 100661 117602 100727 117605
rect 184933 117602 184999 117605
rect 100661 117600 184999 117602
rect 100661 117544 100666 117600
rect 100722 117544 184938 117600
rect 184994 117544 184999 117600
rect 100661 117542 184999 117544
rect 100661 117539 100727 117542
rect 184933 117539 184999 117542
rect 70209 117466 70275 117469
rect 138197 117466 138263 117469
rect 70209 117464 138263 117466
rect 70209 117408 70214 117464
rect 70270 117408 138202 117464
rect 138258 117408 138263 117464
rect 70209 117406 138263 117408
rect 70209 117403 70275 117406
rect 138197 117403 138263 117406
rect 100017 117330 100083 117333
rect 100661 117330 100727 117333
rect 100017 117328 100727 117330
rect 100017 117272 100022 117328
rect 100078 117272 100666 117328
rect 100722 117272 100727 117328
rect 100017 117270 100727 117272
rect 100017 117267 100083 117270
rect 100661 117267 100727 117270
rect 102133 117330 102199 117333
rect 103421 117330 103487 117333
rect 102133 117328 103487 117330
rect 102133 117272 102138 117328
rect 102194 117272 103426 117328
rect 103482 117272 103487 117328
rect 102133 117270 103487 117272
rect 102133 117267 102199 117270
rect 103421 117267 103487 117270
rect 115933 117330 115999 117333
rect 117221 117330 117287 117333
rect 115933 117328 117287 117330
rect 115933 117272 115938 117328
rect 115994 117272 117226 117328
rect 117282 117272 117287 117328
rect 115933 117270 117287 117272
rect 115933 117267 115999 117270
rect 117221 117267 117287 117270
rect 140773 117330 140839 117333
rect 140957 117330 141023 117333
rect 140773 117328 141023 117330
rect 140773 117272 140778 117328
rect 140834 117272 140962 117328
rect 141018 117272 141023 117328
rect 140773 117270 141023 117272
rect 140773 117267 140839 117270
rect 140957 117267 141023 117270
rect 187785 117330 187851 117333
rect 188429 117330 188495 117333
rect 187785 117328 188495 117330
rect 187785 117272 187790 117328
rect 187846 117272 188434 117328
rect 188490 117272 188495 117328
rect 187785 117270 188495 117272
rect 187785 117267 187851 117270
rect 188429 117267 188495 117270
rect 243537 117330 243603 117333
rect 245745 117330 245811 117333
rect 243537 117328 245811 117330
rect 243537 117272 243542 117328
rect 243598 117272 245750 117328
rect 245806 117272 245811 117328
rect 243537 117270 245811 117272
rect 243537 117267 243603 117270
rect 245745 117267 245811 117270
rect 159081 115970 159147 115973
rect 159633 115970 159699 115973
rect 159081 115968 159699 115970
rect 159081 115912 159086 115968
rect 159142 115912 159638 115968
rect 159694 115912 159699 115968
rect 159081 115910 159699 115912
rect 159081 115907 159147 115910
rect 159633 115907 159699 115910
rect 163037 115970 163103 115973
rect 163405 115970 163471 115973
rect 163037 115968 163471 115970
rect 163037 115912 163042 115968
rect 163098 115912 163410 115968
rect 163466 115912 163471 115968
rect 163037 115910 163471 115912
rect 163037 115907 163103 115910
rect 163405 115907 163471 115910
rect 227989 115970 228055 115973
rect 228265 115970 228331 115973
rect 227989 115968 228331 115970
rect 227989 115912 227994 115968
rect 228050 115912 228270 115968
rect 228326 115912 228331 115968
rect 227989 115910 228331 115912
rect 227989 115907 228055 115910
rect 228265 115907 228331 115910
rect 238937 115970 239003 115973
rect 239305 115970 239371 115973
rect 238937 115968 239371 115970
rect 238937 115912 238942 115968
rect 238998 115912 239310 115968
rect 239366 115912 239371 115968
rect 238937 115910 239371 115912
rect 238937 115907 239003 115910
rect 239305 115907 239371 115910
rect 579797 111482 579863 111485
rect 583520 111482 584960 111572
rect 579797 111480 584960 111482
rect 579797 111424 579802 111480
rect 579858 111424 584960 111480
rect 579797 111422 584960 111424
rect 579797 111419 579863 111422
rect 583520 111332 584960 111422
rect -960 107674 480 107764
rect 3509 107674 3575 107677
rect -960 107672 3575 107674
rect -960 107616 3514 107672
rect 3570 107616 3575 107672
rect -960 107614 3575 107616
rect -960 107524 480 107614
rect 3509 107611 3575 107614
rect 133045 106450 133111 106453
rect 133045 106448 133706 106450
rect 133045 106392 133050 106448
rect 133106 106392 133706 106448
rect 133045 106390 133706 106392
rect 133045 106387 133111 106390
rect 133505 106314 133571 106317
rect 133646 106314 133706 106390
rect 133505 106312 133706 106314
rect 133505 106256 133510 106312
rect 133566 106256 133706 106312
rect 133505 106254 133706 106256
rect 183645 106314 183711 106317
rect 183921 106314 183987 106317
rect 183645 106312 183987 106314
rect 183645 106256 183650 106312
rect 183706 106256 183926 106312
rect 183982 106256 183987 106312
rect 183645 106254 183987 106256
rect 133505 106251 133571 106254
rect 183645 106251 183711 106254
rect 183921 106251 183987 106254
rect 184749 106314 184815 106317
rect 184933 106314 184999 106317
rect 184749 106312 184999 106314
rect 184749 106256 184754 106312
rect 184810 106256 184938 106312
rect 184994 106256 184999 106312
rect 184749 106254 184999 106256
rect 184749 106251 184815 106254
rect 184933 106251 184999 106254
rect 233417 106314 233483 106317
rect 233601 106314 233667 106317
rect 233417 106312 233667 106314
rect 233417 106256 233422 106312
rect 233478 106256 233606 106312
rect 233662 106256 233667 106312
rect 233417 106254 233667 106256
rect 233417 106251 233483 106254
rect 233601 106251 233667 106254
rect 341057 106314 341123 106317
rect 341241 106314 341307 106317
rect 341057 106312 341307 106314
rect 341057 106256 341062 106312
rect 341118 106256 341246 106312
rect 341302 106256 341307 106312
rect 341057 106254 341307 106256
rect 341057 106251 341123 106254
rect 341241 106251 341307 106254
rect 388713 106314 388779 106317
rect 388897 106314 388963 106317
rect 388713 106312 388963 106314
rect 388713 106256 388718 106312
rect 388774 106256 388902 106312
rect 388958 106256 388963 106312
rect 388713 106254 388963 106256
rect 388713 106251 388779 106254
rect 388897 106251 388963 106254
rect 194685 104818 194751 104821
rect 194550 104816 194751 104818
rect 194550 104760 194690 104816
rect 194746 104760 194751 104816
rect 194550 104758 194751 104760
rect 194550 104682 194610 104758
rect 194685 104755 194751 104758
rect 194961 104682 195027 104685
rect 194550 104680 195027 104682
rect 194550 104624 194966 104680
rect 195022 104624 195027 104680
rect 194550 104622 195027 104624
rect 194961 104619 195027 104622
rect 211245 100738 211311 100741
rect 211110 100736 211311 100738
rect 211110 100680 211250 100736
rect 211306 100680 211311 100736
rect 211110 100678 211311 100680
rect 211110 100602 211170 100678
rect 211245 100675 211311 100678
rect 211429 100602 211495 100605
rect 211110 100600 211495 100602
rect 211110 100544 211434 100600
rect 211490 100544 211495 100600
rect 211110 100542 211495 100544
rect 211429 100539 211495 100542
rect 583520 99636 584960 99876
rect 238753 96794 238819 96797
rect 238710 96792 238819 96794
rect 238710 96736 238758 96792
rect 238814 96736 238819 96792
rect 238710 96731 238819 96736
rect 137921 96658 137987 96661
rect 138197 96658 138263 96661
rect 137921 96656 138263 96658
rect 137921 96600 137926 96656
rect 137982 96600 138202 96656
rect 138258 96600 138263 96656
rect 137921 96598 138263 96600
rect 137921 96595 137987 96598
rect 138197 96595 138263 96598
rect 183737 96658 183803 96661
rect 183921 96658 183987 96661
rect 183737 96656 183987 96658
rect 183737 96600 183742 96656
rect 183798 96600 183926 96656
rect 183982 96600 183987 96656
rect 183737 96598 183987 96600
rect 238710 96658 238770 96731
rect 238845 96658 238911 96661
rect 238710 96656 238911 96658
rect 238710 96600 238850 96656
rect 238906 96600 238911 96656
rect 238710 96598 238911 96600
rect 183737 96595 183803 96598
rect 183921 96595 183987 96598
rect 238845 96595 238911 96598
rect 279785 93938 279851 93941
rect 279969 93938 280035 93941
rect 279785 93936 280035 93938
rect 279785 93880 279790 93936
rect 279846 93880 279974 93936
rect 280030 93880 280035 93936
rect 279785 93878 280035 93880
rect 279785 93875 279851 93878
rect 279969 93875 280035 93878
rect -960 93258 480 93348
rect 2773 93258 2839 93261
rect -960 93256 2839 93258
rect -960 93200 2778 93256
rect 2834 93200 2839 93256
rect -960 93198 2839 93200
rect -960 93108 480 93198
rect 2773 93195 2839 93198
rect 205909 91082 205975 91085
rect 206093 91082 206159 91085
rect 205909 91080 206159 91082
rect 205909 91024 205914 91080
rect 205970 91024 206098 91080
rect 206154 91024 206159 91080
rect 205909 91022 206159 91024
rect 205909 91019 205975 91022
rect 206093 91019 206159 91022
rect 580165 87954 580231 87957
rect 583520 87954 584960 88044
rect 580165 87952 584960 87954
rect 580165 87896 580170 87952
rect 580226 87896 584960 87952
rect 580165 87894 584960 87896
rect 580165 87891 580231 87894
rect 583520 87804 584960 87894
rect 128721 87002 128787 87005
rect 128997 87002 129063 87005
rect 128721 87000 129063 87002
rect 128721 86944 128726 87000
rect 128782 86944 129002 87000
rect 129058 86944 129063 87000
rect 128721 86942 129063 86944
rect 128721 86939 128787 86942
rect 128997 86939 129063 86942
rect 341057 87002 341123 87005
rect 341241 87002 341307 87005
rect 341057 87000 341307 87002
rect 341057 86944 341062 87000
rect 341118 86944 341246 87000
rect 341302 86944 341307 87000
rect 341057 86942 341307 86944
rect 341057 86939 341123 86942
rect 341241 86939 341307 86942
rect 431585 87002 431651 87005
rect 431769 87002 431835 87005
rect 431585 87000 431835 87002
rect 431585 86944 431590 87000
rect 431646 86944 431774 87000
rect 431830 86944 431835 87000
rect 431585 86942 431835 86944
rect 431585 86939 431651 86942
rect 431769 86939 431835 86942
rect 175641 85640 175707 85645
rect 175641 85584 175646 85640
rect 175702 85584 175707 85640
rect 175641 85579 175707 85584
rect 175644 85506 175704 85579
rect 175825 85506 175891 85509
rect 175644 85504 175891 85506
rect 175644 85448 175830 85504
rect 175886 85448 175891 85504
rect 175644 85446 175891 85448
rect 175825 85443 175891 85446
rect -960 78978 480 79068
rect 3233 78978 3299 78981
rect -960 78976 3299 78978
rect -960 78920 3238 78976
rect 3294 78920 3299 78976
rect -960 78918 3299 78920
rect -960 78828 480 78918
rect 3233 78915 3299 78918
rect 420269 77346 420335 77349
rect 420453 77346 420519 77349
rect 420269 77344 420519 77346
rect 420269 77288 420274 77344
rect 420330 77288 420458 77344
rect 420514 77288 420519 77344
rect 420269 77286 420519 77288
rect 420269 77283 420335 77286
rect 420453 77283 420519 77286
rect 580165 76258 580231 76261
rect 583520 76258 584960 76348
rect 580165 76256 584960 76258
rect 580165 76200 580170 76256
rect 580226 76200 584960 76256
rect 580165 76198 584960 76200
rect 580165 76195 580231 76198
rect 583520 76108 584960 76198
rect 148041 66466 148107 66469
rect 147814 66464 148107 66466
rect 147814 66408 148046 66464
rect 148102 66408 148107 66464
rect 147814 66406 148107 66408
rect 147814 66330 147874 66406
rect 148041 66403 148107 66406
rect 147949 66330 148015 66333
rect 147814 66328 148015 66330
rect 147814 66272 147954 66328
rect 148010 66272 148015 66328
rect 147814 66270 148015 66272
rect 147949 66267 148015 66270
rect -960 64562 480 64652
rect 3325 64562 3391 64565
rect -960 64560 3391 64562
rect -960 64504 3330 64560
rect 3386 64504 3391 64560
rect -960 64502 3391 64504
rect -960 64412 480 64502
rect 3325 64499 3391 64502
rect 579797 64562 579863 64565
rect 583520 64562 584960 64652
rect 579797 64560 584960 64562
rect 579797 64504 579802 64560
rect 579858 64504 584960 64560
rect 579797 64502 584960 64504
rect 579797 64499 579863 64502
rect 583520 64412 584960 64502
rect 420637 61436 420703 61437
rect 420637 61434 420684 61436
rect 420592 61432 420684 61434
rect 420592 61376 420642 61432
rect 420592 61374 420684 61376
rect 420637 61372 420684 61374
rect 420748 61372 420754 61436
rect 420637 61371 420703 61372
rect 211153 56810 211219 56813
rect 211153 56808 211354 56810
rect 211153 56752 211158 56808
rect 211214 56752 211354 56808
rect 211153 56750 211354 56752
rect 211153 56747 211219 56750
rect 211294 56541 211354 56750
rect 211245 56536 211354 56541
rect 211245 56480 211250 56536
rect 211306 56480 211354 56536
rect 211245 56478 211354 56480
rect 211245 56475 211311 56478
rect 583520 52716 584960 52956
rect 178217 52458 178283 52461
rect 178401 52458 178467 52461
rect 178217 52456 178467 52458
rect 178217 52400 178222 52456
rect 178278 52400 178406 52456
rect 178462 52400 178467 52456
rect 178217 52398 178467 52400
rect 178217 52395 178283 52398
rect 178401 52395 178467 52398
rect -960 50146 480 50236
rect 3417 50146 3483 50149
rect -960 50144 3483 50146
rect -960 50088 3422 50144
rect 3478 50088 3483 50144
rect -960 50086 3483 50088
rect -960 49996 480 50086
rect 3417 50083 3483 50086
rect 73981 48514 74047 48517
rect 73478 48512 74047 48514
rect 73478 48456 73986 48512
rect 74042 48456 74047 48512
rect 73478 48454 74047 48456
rect 73478 48378 73538 48454
rect 73981 48451 74047 48454
rect 73613 48378 73679 48381
rect 73478 48376 73679 48378
rect 73478 48320 73618 48376
rect 73674 48320 73679 48376
rect 73478 48318 73679 48320
rect 73613 48315 73679 48318
rect 183737 48378 183803 48381
rect 194961 48378 195027 48381
rect 195145 48378 195211 48381
rect 183737 48376 183938 48378
rect 183737 48320 183742 48376
rect 183798 48320 183938 48376
rect 183737 48318 183938 48320
rect 183737 48315 183803 48318
rect 183686 48044 183692 48108
rect 183756 48106 183762 48108
rect 183878 48106 183938 48318
rect 194961 48376 195211 48378
rect 194961 48320 194966 48376
rect 195022 48320 195150 48376
rect 195206 48320 195211 48376
rect 194961 48318 195211 48320
rect 194961 48315 195027 48318
rect 195145 48315 195211 48318
rect 243445 48378 243511 48381
rect 276105 48378 276171 48381
rect 276289 48378 276355 48381
rect 243445 48376 243554 48378
rect 243445 48320 243450 48376
rect 243506 48320 243554 48376
rect 243445 48315 243554 48320
rect 276105 48376 276355 48378
rect 276105 48320 276110 48376
rect 276166 48320 276294 48376
rect 276350 48320 276355 48376
rect 276105 48318 276355 48320
rect 276105 48315 276171 48318
rect 276289 48315 276355 48318
rect 325509 48378 325575 48381
rect 325693 48378 325759 48381
rect 325509 48376 325759 48378
rect 325509 48320 325514 48376
rect 325570 48320 325698 48376
rect 325754 48320 325759 48376
rect 325509 48318 325759 48320
rect 325509 48315 325575 48318
rect 325693 48315 325759 48318
rect 415025 48378 415091 48381
rect 415209 48378 415275 48381
rect 415025 48376 415275 48378
rect 415025 48320 415030 48376
rect 415086 48320 415214 48376
rect 415270 48320 415275 48376
rect 415025 48318 415275 48320
rect 415025 48315 415091 48318
rect 415209 48315 415275 48318
rect 420545 48378 420611 48381
rect 420678 48378 420684 48380
rect 420545 48376 420684 48378
rect 420545 48320 420550 48376
rect 420606 48320 420684 48376
rect 420545 48318 420684 48320
rect 420545 48315 420611 48318
rect 420678 48316 420684 48318
rect 420748 48316 420754 48380
rect 426065 48378 426131 48381
rect 426249 48378 426315 48381
rect 426065 48376 426315 48378
rect 426065 48320 426070 48376
rect 426126 48320 426254 48376
rect 426310 48320 426315 48376
rect 426065 48318 426315 48320
rect 426065 48315 426131 48318
rect 426249 48315 426315 48318
rect 243494 48245 243554 48315
rect 243445 48240 243554 48245
rect 243445 48184 243450 48240
rect 243506 48184 243554 48240
rect 243445 48182 243554 48184
rect 243445 48179 243511 48182
rect 183756 48046 183938 48106
rect 183756 48044 183762 48046
rect 431585 47018 431651 47021
rect 431769 47018 431835 47021
rect 431585 47016 431835 47018
rect 431585 46960 431590 47016
rect 431646 46960 431774 47016
rect 431830 46960 431835 47016
rect 431585 46958 431835 46960
rect 431585 46955 431651 46958
rect 431769 46955 431835 46958
rect 211337 45522 211403 45525
rect 211521 45522 211587 45525
rect 211337 45520 211587 45522
rect 211337 45464 211342 45520
rect 211398 45464 211526 45520
rect 211582 45464 211587 45520
rect 211337 45462 211587 45464
rect 211337 45459 211403 45462
rect 211521 45459 211587 45462
rect 420637 42124 420703 42125
rect 420637 42122 420684 42124
rect 420592 42120 420684 42122
rect 420592 42064 420642 42120
rect 420592 42062 420684 42064
rect 420637 42060 420684 42062
rect 420748 42060 420754 42124
rect 420637 42059 420703 42060
rect 580165 41034 580231 41037
rect 583520 41034 584960 41124
rect 580165 41032 584960 41034
rect 580165 40976 580170 41032
rect 580226 40976 584960 41032
rect 580165 40974 584960 40976
rect 580165 40971 580231 40974
rect 583520 40884 584960 40974
rect 183645 38724 183711 38725
rect 183645 38722 183692 38724
rect 183600 38720 183692 38722
rect 183600 38664 183650 38720
rect 183600 38662 183692 38664
rect 183645 38660 183692 38662
rect 183756 38660 183762 38724
rect 183645 38659 183711 38660
rect -960 35866 480 35956
rect 3417 35866 3483 35869
rect -960 35864 3483 35866
rect -960 35808 3422 35864
rect 3478 35808 3483 35864
rect -960 35806 3483 35808
rect -960 35716 480 35806
rect 3417 35803 3483 35806
rect 73613 34506 73679 34509
rect 73797 34506 73863 34509
rect 73613 34504 73863 34506
rect 73613 34448 73618 34504
rect 73674 34448 73802 34504
rect 73858 34448 73863 34504
rect 73613 34446 73863 34448
rect 73613 34443 73679 34446
rect 73797 34443 73863 34446
rect 580165 29338 580231 29341
rect 583520 29338 584960 29428
rect 580165 29336 584960 29338
rect 580165 29280 580170 29336
rect 580226 29280 584960 29336
rect 580165 29278 584960 29280
rect 580165 29275 580231 29278
rect 583520 29188 584960 29278
rect 420545 29066 420611 29069
rect 420678 29066 420684 29068
rect 420545 29064 420684 29066
rect 420545 29008 420550 29064
rect 420606 29008 420684 29064
rect 420545 29006 420684 29008
rect 420545 29003 420611 29006
rect 420678 29004 420684 29006
rect 420748 29004 420754 29068
rect 301865 26346 301931 26349
rect 302049 26346 302115 26349
rect 301865 26344 302115 26346
rect 301865 26288 301870 26344
rect 301926 26288 302054 26344
rect 302110 26288 302115 26344
rect 301865 26286 302115 26288
rect 301865 26283 301931 26286
rect 302049 26283 302115 26286
rect 178125 22130 178191 22133
rect 178401 22130 178467 22133
rect 178125 22128 178467 22130
rect 178125 22072 178130 22128
rect 178186 22072 178406 22128
rect 178462 22072 178467 22128
rect 178125 22070 178467 22072
rect 178125 22067 178191 22070
rect 178401 22067 178467 22070
rect -960 21450 480 21540
rect 3141 21450 3207 21453
rect -960 21448 3207 21450
rect -960 21392 3146 21448
rect 3202 21392 3207 21448
rect -960 21390 3207 21392
rect -960 21300 480 21390
rect 3141 21387 3207 21390
rect 207289 19410 207355 19413
rect 207062 19408 207355 19410
rect 207062 19352 207294 19408
rect 207350 19352 207355 19408
rect 207062 19350 207355 19352
rect 207062 19274 207122 19350
rect 207289 19347 207355 19350
rect 207289 19274 207355 19277
rect 207062 19272 207355 19274
rect 207062 19216 207294 19272
rect 207350 19216 207355 19272
rect 207062 19214 207355 19216
rect 207289 19211 207355 19214
rect 228909 19274 228975 19277
rect 229093 19274 229159 19277
rect 228909 19272 229159 19274
rect 228909 19216 228914 19272
rect 228970 19216 229098 19272
rect 229154 19216 229159 19272
rect 228909 19214 229159 19216
rect 228909 19211 228975 19214
rect 229093 19211 229159 19214
rect 579797 17642 579863 17645
rect 583520 17642 584960 17732
rect 579797 17640 584960 17642
rect 579797 17584 579802 17640
rect 579858 17584 584960 17640
rect 579797 17582 584960 17584
rect 579797 17579 579863 17582
rect 583520 17492 584960 17582
rect -960 7170 480 7260
rect 3417 7170 3483 7173
rect -960 7168 3483 7170
rect -960 7112 3422 7168
rect 3478 7112 3483 7168
rect -960 7110 3483 7112
rect -960 7020 480 7110
rect 3417 7107 3483 7110
rect 113541 6218 113607 6221
rect 192017 6218 192083 6221
rect 113541 6216 192083 6218
rect 113541 6160 113546 6216
rect 113602 6160 192022 6216
rect 192078 6160 192083 6216
rect 113541 6158 192083 6160
rect 113541 6155 113607 6158
rect 192017 6155 192083 6158
rect 411069 6218 411135 6221
rect 538121 6218 538187 6221
rect 411069 6216 538187 6218
rect 411069 6160 411074 6216
rect 411130 6160 538126 6216
rect 538182 6160 538187 6216
rect 411069 6158 538187 6160
rect 411069 6155 411135 6158
rect 538121 6155 538187 6158
rect 583520 5796 584960 6036
rect 30281 4858 30347 4861
rect 149053 4858 149119 4861
rect 30281 4856 149119 4858
rect 30281 4800 30286 4856
rect 30342 4800 149058 4856
rect 149114 4800 149119 4856
rect 30281 4798 149119 4800
rect 30281 4795 30347 4798
rect 149053 4795 149119 4798
rect 357341 4858 357407 4861
rect 433517 4858 433583 4861
rect 357341 4856 433583 4858
rect 357341 4800 357346 4856
rect 357402 4800 433522 4856
rect 433578 4800 433583 4856
rect 357341 4798 433583 4800
rect 357341 4795 357407 4798
rect 433517 4795 433583 4798
rect 408309 3770 408375 3773
rect 408493 3770 408559 3773
rect 408309 3768 408559 3770
rect 408309 3712 408314 3768
rect 408370 3712 408498 3768
rect 408554 3712 408559 3768
rect 408309 3710 408559 3712
rect 408309 3707 408375 3710
rect 408493 3707 408559 3710
rect 417877 3634 417943 3637
rect 418337 3634 418403 3637
rect 417877 3632 418403 3634
rect 417877 3576 417882 3632
rect 417938 3576 418342 3632
rect 418398 3576 418403 3632
rect 417877 3574 418403 3576
rect 417877 3571 417943 3574
rect 418337 3571 418403 3574
rect 431217 3362 431283 3365
rect 575013 3362 575079 3365
rect 431217 3360 575079 3362
rect 431217 3304 431222 3360
rect 431278 3304 575018 3360
rect 575074 3304 575079 3360
rect 431217 3302 575079 3304
rect 431217 3299 431283 3302
rect 575013 3299 575079 3302
<< via3 >>
rect 132172 700436 132236 700500
rect 132356 700300 132420 700364
rect 133644 697172 133708 697236
rect 164188 686428 164252 686492
rect 131988 685884 132052 685948
rect 164188 686156 164252 686220
rect 164188 650524 164252 650588
rect 133460 650252 133524 650316
rect 164188 650252 164252 650316
rect 131804 638964 131868 639028
rect 164188 639100 164252 639164
rect 164188 638828 164252 638892
rect 133092 603332 133156 603396
rect 164188 603196 164252 603260
rect 164188 602924 164252 602988
rect 164188 592588 164252 592652
rect 133276 592316 133340 592380
rect 164188 592316 164252 592380
rect 380020 572052 380084 572116
rect 379468 563076 379532 563140
rect 199700 561716 199764 561780
rect 379652 559540 379716 559604
rect 198596 556684 198660 556748
rect 198412 552060 198476 552124
rect 198228 547844 198292 547908
rect 198044 543764 198108 543828
rect 380204 541044 380268 541108
rect 197860 538460 197924 538524
rect 379836 528668 379900 528732
rect 380204 500244 380268 500308
rect 380020 500108 380084 500172
rect 125916 495544 125980 495548
rect 125916 495488 125966 495544
rect 125966 495488 125980 495544
rect 125916 495484 125980 495488
rect 125916 492688 125980 492692
rect 125916 492632 125930 492688
rect 125930 492632 125980 492688
rect 125916 492628 125980 492632
rect 153332 447264 153396 447268
rect 153332 447208 153382 447264
rect 153382 447208 153396 447264
rect 153332 447204 153396 447208
rect 153332 444408 153396 444412
rect 153332 444352 153382 444408
rect 153382 444352 153396 444408
rect 153332 444348 153396 444352
rect 379836 417420 379900 417484
rect 266860 410348 266924 410412
rect 267780 410212 267844 410276
rect 267964 410076 268028 410140
rect 268148 409940 268212 410004
rect 379468 394632 379532 394636
rect 379468 394576 379518 394632
rect 379518 394576 379532 394632
rect 379468 394572 379532 394576
rect 379652 394496 379716 394500
rect 379652 394440 379666 394496
rect 379666 394440 379716 394496
rect 379652 394436 379716 394440
rect 283972 380156 284036 380220
rect 283972 367236 284036 367300
rect 268148 338676 268212 338740
rect 391060 318684 391124 318748
rect 257660 317384 257724 317388
rect 257660 317328 257710 317384
rect 257710 317328 257724 317384
rect 257660 317324 257724 317328
rect 257660 311748 257724 311812
rect 391060 309164 391124 309228
rect 391060 299372 391124 299436
rect 297772 298012 297836 298076
rect 391060 289852 391124 289916
rect 297772 288492 297836 288556
rect 391060 280060 391124 280124
rect 391060 270540 391124 270604
rect 266860 202812 266924 202876
rect 197860 202540 197924 202604
rect 198228 202268 198292 202332
rect 267780 202132 267844 202196
rect 199700 201996 199764 202060
rect 198412 201860 198476 201924
rect 198596 201724 198660 201788
rect 198044 201588 198108 201652
rect 267964 201588 268028 201652
rect 132908 200636 132972 200700
rect 132908 176156 132972 176220
rect 133644 175068 133708 175132
rect 133460 173980 133524 174044
rect 133092 172892 133156 172956
rect 132172 137124 132236 137188
rect 132356 136172 132420 136236
rect 131988 135084 132052 135148
rect 131804 133996 131868 134060
rect 133276 132908 133340 132972
rect 420684 61432 420748 61436
rect 420684 61376 420698 61432
rect 420698 61376 420748 61432
rect 420684 61372 420748 61376
rect 183692 48044 183756 48108
rect 420684 48316 420748 48380
rect 420684 42120 420748 42124
rect 420684 42064 420698 42120
rect 420698 42064 420748 42120
rect 420684 42060 420748 42064
rect 183692 38720 183756 38724
rect 183692 38664 183706 38720
rect 183706 38664 183756 38720
rect 183692 38660 183756 38664
rect 420684 29004 420748 29068
<< metal4 >>
rect -8576 711418 -7976 711440
rect -8576 711182 -8394 711418
rect -8158 711182 -7976 711418
rect -8576 711098 -7976 711182
rect -8576 710862 -8394 711098
rect -8158 710862 -7976 711098
rect -8576 679254 -7976 710862
rect -8576 679018 -8394 679254
rect -8158 679018 -7976 679254
rect -8576 678934 -7976 679018
rect -8576 678698 -8394 678934
rect -8158 678698 -7976 678934
rect -8576 643254 -7976 678698
rect -8576 643018 -8394 643254
rect -8158 643018 -7976 643254
rect -8576 642934 -7976 643018
rect -8576 642698 -8394 642934
rect -8158 642698 -7976 642934
rect -8576 607254 -7976 642698
rect -8576 607018 -8394 607254
rect -8158 607018 -7976 607254
rect -8576 606934 -7976 607018
rect -8576 606698 -8394 606934
rect -8158 606698 -7976 606934
rect -8576 571254 -7976 606698
rect -8576 571018 -8394 571254
rect -8158 571018 -7976 571254
rect -8576 570934 -7976 571018
rect -8576 570698 -8394 570934
rect -8158 570698 -7976 570934
rect -8576 535254 -7976 570698
rect -8576 535018 -8394 535254
rect -8158 535018 -7976 535254
rect -8576 534934 -7976 535018
rect -8576 534698 -8394 534934
rect -8158 534698 -7976 534934
rect -8576 499254 -7976 534698
rect -8576 499018 -8394 499254
rect -8158 499018 -7976 499254
rect -8576 498934 -7976 499018
rect -8576 498698 -8394 498934
rect -8158 498698 -7976 498934
rect -8576 463254 -7976 498698
rect -8576 463018 -8394 463254
rect -8158 463018 -7976 463254
rect -8576 462934 -7976 463018
rect -8576 462698 -8394 462934
rect -8158 462698 -7976 462934
rect -8576 427254 -7976 462698
rect -8576 427018 -8394 427254
rect -8158 427018 -7976 427254
rect -8576 426934 -7976 427018
rect -8576 426698 -8394 426934
rect -8158 426698 -7976 426934
rect -8576 391254 -7976 426698
rect -8576 391018 -8394 391254
rect -8158 391018 -7976 391254
rect -8576 390934 -7976 391018
rect -8576 390698 -8394 390934
rect -8158 390698 -7976 390934
rect -8576 355254 -7976 390698
rect -8576 355018 -8394 355254
rect -8158 355018 -7976 355254
rect -8576 354934 -7976 355018
rect -8576 354698 -8394 354934
rect -8158 354698 -7976 354934
rect -8576 319254 -7976 354698
rect -8576 319018 -8394 319254
rect -8158 319018 -7976 319254
rect -8576 318934 -7976 319018
rect -8576 318698 -8394 318934
rect -8158 318698 -7976 318934
rect -8576 283254 -7976 318698
rect -8576 283018 -8394 283254
rect -8158 283018 -7976 283254
rect -8576 282934 -7976 283018
rect -8576 282698 -8394 282934
rect -8158 282698 -7976 282934
rect -8576 247254 -7976 282698
rect -8576 247018 -8394 247254
rect -8158 247018 -7976 247254
rect -8576 246934 -7976 247018
rect -8576 246698 -8394 246934
rect -8158 246698 -7976 246934
rect -8576 211254 -7976 246698
rect -8576 211018 -8394 211254
rect -8158 211018 -7976 211254
rect -8576 210934 -7976 211018
rect -8576 210698 -8394 210934
rect -8158 210698 -7976 210934
rect -8576 175254 -7976 210698
rect -8576 175018 -8394 175254
rect -8158 175018 -7976 175254
rect -8576 174934 -7976 175018
rect -8576 174698 -8394 174934
rect -8158 174698 -7976 174934
rect -8576 139254 -7976 174698
rect -8576 139018 -8394 139254
rect -8158 139018 -7976 139254
rect -8576 138934 -7976 139018
rect -8576 138698 -8394 138934
rect -8158 138698 -7976 138934
rect -8576 103254 -7976 138698
rect -8576 103018 -8394 103254
rect -8158 103018 -7976 103254
rect -8576 102934 -7976 103018
rect -8576 102698 -8394 102934
rect -8158 102698 -7976 102934
rect -8576 67254 -7976 102698
rect -8576 67018 -8394 67254
rect -8158 67018 -7976 67254
rect -8576 66934 -7976 67018
rect -8576 66698 -8394 66934
rect -8158 66698 -7976 66934
rect -8576 31254 -7976 66698
rect -8576 31018 -8394 31254
rect -8158 31018 -7976 31254
rect -8576 30934 -7976 31018
rect -8576 30698 -8394 30934
rect -8158 30698 -7976 30934
rect -8576 -6926 -7976 30698
rect -7636 710478 -7036 710500
rect -7636 710242 -7454 710478
rect -7218 710242 -7036 710478
rect -7636 710158 -7036 710242
rect -7636 709922 -7454 710158
rect -7218 709922 -7036 710158
rect -7636 697254 -7036 709922
rect 11604 710478 12204 711440
rect 11604 710242 11786 710478
rect 12022 710242 12204 710478
rect 11604 710158 12204 710242
rect 11604 709922 11786 710158
rect 12022 709922 12204 710158
rect -7636 697018 -7454 697254
rect -7218 697018 -7036 697254
rect -7636 696934 -7036 697018
rect -7636 696698 -7454 696934
rect -7218 696698 -7036 696934
rect -7636 661254 -7036 696698
rect -7636 661018 -7454 661254
rect -7218 661018 -7036 661254
rect -7636 660934 -7036 661018
rect -7636 660698 -7454 660934
rect -7218 660698 -7036 660934
rect -7636 625254 -7036 660698
rect -7636 625018 -7454 625254
rect -7218 625018 -7036 625254
rect -7636 624934 -7036 625018
rect -7636 624698 -7454 624934
rect -7218 624698 -7036 624934
rect -7636 589254 -7036 624698
rect -7636 589018 -7454 589254
rect -7218 589018 -7036 589254
rect -7636 588934 -7036 589018
rect -7636 588698 -7454 588934
rect -7218 588698 -7036 588934
rect -7636 553254 -7036 588698
rect -7636 553018 -7454 553254
rect -7218 553018 -7036 553254
rect -7636 552934 -7036 553018
rect -7636 552698 -7454 552934
rect -7218 552698 -7036 552934
rect -7636 517254 -7036 552698
rect -7636 517018 -7454 517254
rect -7218 517018 -7036 517254
rect -7636 516934 -7036 517018
rect -7636 516698 -7454 516934
rect -7218 516698 -7036 516934
rect -7636 481254 -7036 516698
rect -7636 481018 -7454 481254
rect -7218 481018 -7036 481254
rect -7636 480934 -7036 481018
rect -7636 480698 -7454 480934
rect -7218 480698 -7036 480934
rect -7636 445254 -7036 480698
rect -7636 445018 -7454 445254
rect -7218 445018 -7036 445254
rect -7636 444934 -7036 445018
rect -7636 444698 -7454 444934
rect -7218 444698 -7036 444934
rect -7636 409254 -7036 444698
rect -7636 409018 -7454 409254
rect -7218 409018 -7036 409254
rect -7636 408934 -7036 409018
rect -7636 408698 -7454 408934
rect -7218 408698 -7036 408934
rect -7636 373254 -7036 408698
rect -7636 373018 -7454 373254
rect -7218 373018 -7036 373254
rect -7636 372934 -7036 373018
rect -7636 372698 -7454 372934
rect -7218 372698 -7036 372934
rect -7636 337254 -7036 372698
rect -7636 337018 -7454 337254
rect -7218 337018 -7036 337254
rect -7636 336934 -7036 337018
rect -7636 336698 -7454 336934
rect -7218 336698 -7036 336934
rect -7636 301254 -7036 336698
rect -7636 301018 -7454 301254
rect -7218 301018 -7036 301254
rect -7636 300934 -7036 301018
rect -7636 300698 -7454 300934
rect -7218 300698 -7036 300934
rect -7636 265254 -7036 300698
rect -7636 265018 -7454 265254
rect -7218 265018 -7036 265254
rect -7636 264934 -7036 265018
rect -7636 264698 -7454 264934
rect -7218 264698 -7036 264934
rect -7636 229254 -7036 264698
rect -7636 229018 -7454 229254
rect -7218 229018 -7036 229254
rect -7636 228934 -7036 229018
rect -7636 228698 -7454 228934
rect -7218 228698 -7036 228934
rect -7636 193254 -7036 228698
rect -7636 193018 -7454 193254
rect -7218 193018 -7036 193254
rect -7636 192934 -7036 193018
rect -7636 192698 -7454 192934
rect -7218 192698 -7036 192934
rect -7636 157254 -7036 192698
rect -7636 157018 -7454 157254
rect -7218 157018 -7036 157254
rect -7636 156934 -7036 157018
rect -7636 156698 -7454 156934
rect -7218 156698 -7036 156934
rect -7636 121254 -7036 156698
rect -7636 121018 -7454 121254
rect -7218 121018 -7036 121254
rect -7636 120934 -7036 121018
rect -7636 120698 -7454 120934
rect -7218 120698 -7036 120934
rect -7636 85254 -7036 120698
rect -7636 85018 -7454 85254
rect -7218 85018 -7036 85254
rect -7636 84934 -7036 85018
rect -7636 84698 -7454 84934
rect -7218 84698 -7036 84934
rect -7636 49254 -7036 84698
rect -7636 49018 -7454 49254
rect -7218 49018 -7036 49254
rect -7636 48934 -7036 49018
rect -7636 48698 -7454 48934
rect -7218 48698 -7036 48934
rect -7636 13254 -7036 48698
rect -7636 13018 -7454 13254
rect -7218 13018 -7036 13254
rect -7636 12934 -7036 13018
rect -7636 12698 -7454 12934
rect -7218 12698 -7036 12934
rect -7636 -5986 -7036 12698
rect -6696 709538 -6096 709560
rect -6696 709302 -6514 709538
rect -6278 709302 -6096 709538
rect -6696 709218 -6096 709302
rect -6696 708982 -6514 709218
rect -6278 708982 -6096 709218
rect -6696 675654 -6096 708982
rect -6696 675418 -6514 675654
rect -6278 675418 -6096 675654
rect -6696 675334 -6096 675418
rect -6696 675098 -6514 675334
rect -6278 675098 -6096 675334
rect -6696 639654 -6096 675098
rect -6696 639418 -6514 639654
rect -6278 639418 -6096 639654
rect -6696 639334 -6096 639418
rect -6696 639098 -6514 639334
rect -6278 639098 -6096 639334
rect -6696 603654 -6096 639098
rect -6696 603418 -6514 603654
rect -6278 603418 -6096 603654
rect -6696 603334 -6096 603418
rect -6696 603098 -6514 603334
rect -6278 603098 -6096 603334
rect -6696 567654 -6096 603098
rect -6696 567418 -6514 567654
rect -6278 567418 -6096 567654
rect -6696 567334 -6096 567418
rect -6696 567098 -6514 567334
rect -6278 567098 -6096 567334
rect -6696 531654 -6096 567098
rect -6696 531418 -6514 531654
rect -6278 531418 -6096 531654
rect -6696 531334 -6096 531418
rect -6696 531098 -6514 531334
rect -6278 531098 -6096 531334
rect -6696 495654 -6096 531098
rect -6696 495418 -6514 495654
rect -6278 495418 -6096 495654
rect -6696 495334 -6096 495418
rect -6696 495098 -6514 495334
rect -6278 495098 -6096 495334
rect -6696 459654 -6096 495098
rect -6696 459418 -6514 459654
rect -6278 459418 -6096 459654
rect -6696 459334 -6096 459418
rect -6696 459098 -6514 459334
rect -6278 459098 -6096 459334
rect -6696 423654 -6096 459098
rect -6696 423418 -6514 423654
rect -6278 423418 -6096 423654
rect -6696 423334 -6096 423418
rect -6696 423098 -6514 423334
rect -6278 423098 -6096 423334
rect -6696 387654 -6096 423098
rect -6696 387418 -6514 387654
rect -6278 387418 -6096 387654
rect -6696 387334 -6096 387418
rect -6696 387098 -6514 387334
rect -6278 387098 -6096 387334
rect -6696 351654 -6096 387098
rect -6696 351418 -6514 351654
rect -6278 351418 -6096 351654
rect -6696 351334 -6096 351418
rect -6696 351098 -6514 351334
rect -6278 351098 -6096 351334
rect -6696 315654 -6096 351098
rect -6696 315418 -6514 315654
rect -6278 315418 -6096 315654
rect -6696 315334 -6096 315418
rect -6696 315098 -6514 315334
rect -6278 315098 -6096 315334
rect -6696 279654 -6096 315098
rect -6696 279418 -6514 279654
rect -6278 279418 -6096 279654
rect -6696 279334 -6096 279418
rect -6696 279098 -6514 279334
rect -6278 279098 -6096 279334
rect -6696 243654 -6096 279098
rect -6696 243418 -6514 243654
rect -6278 243418 -6096 243654
rect -6696 243334 -6096 243418
rect -6696 243098 -6514 243334
rect -6278 243098 -6096 243334
rect -6696 207654 -6096 243098
rect -6696 207418 -6514 207654
rect -6278 207418 -6096 207654
rect -6696 207334 -6096 207418
rect -6696 207098 -6514 207334
rect -6278 207098 -6096 207334
rect -6696 171654 -6096 207098
rect -6696 171418 -6514 171654
rect -6278 171418 -6096 171654
rect -6696 171334 -6096 171418
rect -6696 171098 -6514 171334
rect -6278 171098 -6096 171334
rect -6696 135654 -6096 171098
rect -6696 135418 -6514 135654
rect -6278 135418 -6096 135654
rect -6696 135334 -6096 135418
rect -6696 135098 -6514 135334
rect -6278 135098 -6096 135334
rect -6696 99654 -6096 135098
rect -6696 99418 -6514 99654
rect -6278 99418 -6096 99654
rect -6696 99334 -6096 99418
rect -6696 99098 -6514 99334
rect -6278 99098 -6096 99334
rect -6696 63654 -6096 99098
rect -6696 63418 -6514 63654
rect -6278 63418 -6096 63654
rect -6696 63334 -6096 63418
rect -6696 63098 -6514 63334
rect -6278 63098 -6096 63334
rect -6696 27654 -6096 63098
rect -6696 27418 -6514 27654
rect -6278 27418 -6096 27654
rect -6696 27334 -6096 27418
rect -6696 27098 -6514 27334
rect -6278 27098 -6096 27334
rect -6696 -5046 -6096 27098
rect -5756 708598 -5156 708620
rect -5756 708362 -5574 708598
rect -5338 708362 -5156 708598
rect -5756 708278 -5156 708362
rect -5756 708042 -5574 708278
rect -5338 708042 -5156 708278
rect -5756 693654 -5156 708042
rect 8004 708598 8604 709560
rect 8004 708362 8186 708598
rect 8422 708362 8604 708598
rect 8004 708278 8604 708362
rect 8004 708042 8186 708278
rect 8422 708042 8604 708278
rect -5756 693418 -5574 693654
rect -5338 693418 -5156 693654
rect -5756 693334 -5156 693418
rect -5756 693098 -5574 693334
rect -5338 693098 -5156 693334
rect -5756 657654 -5156 693098
rect -5756 657418 -5574 657654
rect -5338 657418 -5156 657654
rect -5756 657334 -5156 657418
rect -5756 657098 -5574 657334
rect -5338 657098 -5156 657334
rect -5756 621654 -5156 657098
rect -5756 621418 -5574 621654
rect -5338 621418 -5156 621654
rect -5756 621334 -5156 621418
rect -5756 621098 -5574 621334
rect -5338 621098 -5156 621334
rect -5756 585654 -5156 621098
rect -5756 585418 -5574 585654
rect -5338 585418 -5156 585654
rect -5756 585334 -5156 585418
rect -5756 585098 -5574 585334
rect -5338 585098 -5156 585334
rect -5756 549654 -5156 585098
rect -5756 549418 -5574 549654
rect -5338 549418 -5156 549654
rect -5756 549334 -5156 549418
rect -5756 549098 -5574 549334
rect -5338 549098 -5156 549334
rect -5756 513654 -5156 549098
rect -5756 513418 -5574 513654
rect -5338 513418 -5156 513654
rect -5756 513334 -5156 513418
rect -5756 513098 -5574 513334
rect -5338 513098 -5156 513334
rect -5756 477654 -5156 513098
rect -5756 477418 -5574 477654
rect -5338 477418 -5156 477654
rect -5756 477334 -5156 477418
rect -5756 477098 -5574 477334
rect -5338 477098 -5156 477334
rect -5756 441654 -5156 477098
rect -5756 441418 -5574 441654
rect -5338 441418 -5156 441654
rect -5756 441334 -5156 441418
rect -5756 441098 -5574 441334
rect -5338 441098 -5156 441334
rect -5756 405654 -5156 441098
rect -5756 405418 -5574 405654
rect -5338 405418 -5156 405654
rect -5756 405334 -5156 405418
rect -5756 405098 -5574 405334
rect -5338 405098 -5156 405334
rect -5756 369654 -5156 405098
rect -5756 369418 -5574 369654
rect -5338 369418 -5156 369654
rect -5756 369334 -5156 369418
rect -5756 369098 -5574 369334
rect -5338 369098 -5156 369334
rect -5756 333654 -5156 369098
rect -5756 333418 -5574 333654
rect -5338 333418 -5156 333654
rect -5756 333334 -5156 333418
rect -5756 333098 -5574 333334
rect -5338 333098 -5156 333334
rect -5756 297654 -5156 333098
rect -5756 297418 -5574 297654
rect -5338 297418 -5156 297654
rect -5756 297334 -5156 297418
rect -5756 297098 -5574 297334
rect -5338 297098 -5156 297334
rect -5756 261654 -5156 297098
rect -5756 261418 -5574 261654
rect -5338 261418 -5156 261654
rect -5756 261334 -5156 261418
rect -5756 261098 -5574 261334
rect -5338 261098 -5156 261334
rect -5756 225654 -5156 261098
rect -5756 225418 -5574 225654
rect -5338 225418 -5156 225654
rect -5756 225334 -5156 225418
rect -5756 225098 -5574 225334
rect -5338 225098 -5156 225334
rect -5756 189654 -5156 225098
rect -5756 189418 -5574 189654
rect -5338 189418 -5156 189654
rect -5756 189334 -5156 189418
rect -5756 189098 -5574 189334
rect -5338 189098 -5156 189334
rect -5756 153654 -5156 189098
rect -5756 153418 -5574 153654
rect -5338 153418 -5156 153654
rect -5756 153334 -5156 153418
rect -5756 153098 -5574 153334
rect -5338 153098 -5156 153334
rect -5756 117654 -5156 153098
rect -5756 117418 -5574 117654
rect -5338 117418 -5156 117654
rect -5756 117334 -5156 117418
rect -5756 117098 -5574 117334
rect -5338 117098 -5156 117334
rect -5756 81654 -5156 117098
rect -5756 81418 -5574 81654
rect -5338 81418 -5156 81654
rect -5756 81334 -5156 81418
rect -5756 81098 -5574 81334
rect -5338 81098 -5156 81334
rect -5756 45654 -5156 81098
rect -5756 45418 -5574 45654
rect -5338 45418 -5156 45654
rect -5756 45334 -5156 45418
rect -5756 45098 -5574 45334
rect -5338 45098 -5156 45334
rect -5756 9654 -5156 45098
rect -5756 9418 -5574 9654
rect -5338 9418 -5156 9654
rect -5756 9334 -5156 9418
rect -5756 9098 -5574 9334
rect -5338 9098 -5156 9334
rect -5756 -4106 -5156 9098
rect -4816 707658 -4216 707680
rect -4816 707422 -4634 707658
rect -4398 707422 -4216 707658
rect -4816 707338 -4216 707422
rect -4816 707102 -4634 707338
rect -4398 707102 -4216 707338
rect -4816 672054 -4216 707102
rect -4816 671818 -4634 672054
rect -4398 671818 -4216 672054
rect -4816 671734 -4216 671818
rect -4816 671498 -4634 671734
rect -4398 671498 -4216 671734
rect -4816 636054 -4216 671498
rect -4816 635818 -4634 636054
rect -4398 635818 -4216 636054
rect -4816 635734 -4216 635818
rect -4816 635498 -4634 635734
rect -4398 635498 -4216 635734
rect -4816 600054 -4216 635498
rect -4816 599818 -4634 600054
rect -4398 599818 -4216 600054
rect -4816 599734 -4216 599818
rect -4816 599498 -4634 599734
rect -4398 599498 -4216 599734
rect -4816 564054 -4216 599498
rect -4816 563818 -4634 564054
rect -4398 563818 -4216 564054
rect -4816 563734 -4216 563818
rect -4816 563498 -4634 563734
rect -4398 563498 -4216 563734
rect -4816 528054 -4216 563498
rect -4816 527818 -4634 528054
rect -4398 527818 -4216 528054
rect -4816 527734 -4216 527818
rect -4816 527498 -4634 527734
rect -4398 527498 -4216 527734
rect -4816 492054 -4216 527498
rect -4816 491818 -4634 492054
rect -4398 491818 -4216 492054
rect -4816 491734 -4216 491818
rect -4816 491498 -4634 491734
rect -4398 491498 -4216 491734
rect -4816 456054 -4216 491498
rect -4816 455818 -4634 456054
rect -4398 455818 -4216 456054
rect -4816 455734 -4216 455818
rect -4816 455498 -4634 455734
rect -4398 455498 -4216 455734
rect -4816 420054 -4216 455498
rect -4816 419818 -4634 420054
rect -4398 419818 -4216 420054
rect -4816 419734 -4216 419818
rect -4816 419498 -4634 419734
rect -4398 419498 -4216 419734
rect -4816 384054 -4216 419498
rect -4816 383818 -4634 384054
rect -4398 383818 -4216 384054
rect -4816 383734 -4216 383818
rect -4816 383498 -4634 383734
rect -4398 383498 -4216 383734
rect -4816 348054 -4216 383498
rect -4816 347818 -4634 348054
rect -4398 347818 -4216 348054
rect -4816 347734 -4216 347818
rect -4816 347498 -4634 347734
rect -4398 347498 -4216 347734
rect -4816 312054 -4216 347498
rect -4816 311818 -4634 312054
rect -4398 311818 -4216 312054
rect -4816 311734 -4216 311818
rect -4816 311498 -4634 311734
rect -4398 311498 -4216 311734
rect -4816 276054 -4216 311498
rect -4816 275818 -4634 276054
rect -4398 275818 -4216 276054
rect -4816 275734 -4216 275818
rect -4816 275498 -4634 275734
rect -4398 275498 -4216 275734
rect -4816 240054 -4216 275498
rect -4816 239818 -4634 240054
rect -4398 239818 -4216 240054
rect -4816 239734 -4216 239818
rect -4816 239498 -4634 239734
rect -4398 239498 -4216 239734
rect -4816 204054 -4216 239498
rect -4816 203818 -4634 204054
rect -4398 203818 -4216 204054
rect -4816 203734 -4216 203818
rect -4816 203498 -4634 203734
rect -4398 203498 -4216 203734
rect -4816 168054 -4216 203498
rect -4816 167818 -4634 168054
rect -4398 167818 -4216 168054
rect -4816 167734 -4216 167818
rect -4816 167498 -4634 167734
rect -4398 167498 -4216 167734
rect -4816 132054 -4216 167498
rect -4816 131818 -4634 132054
rect -4398 131818 -4216 132054
rect -4816 131734 -4216 131818
rect -4816 131498 -4634 131734
rect -4398 131498 -4216 131734
rect -4816 96054 -4216 131498
rect -4816 95818 -4634 96054
rect -4398 95818 -4216 96054
rect -4816 95734 -4216 95818
rect -4816 95498 -4634 95734
rect -4398 95498 -4216 95734
rect -4816 60054 -4216 95498
rect -4816 59818 -4634 60054
rect -4398 59818 -4216 60054
rect -4816 59734 -4216 59818
rect -4816 59498 -4634 59734
rect -4398 59498 -4216 59734
rect -4816 24054 -4216 59498
rect -4816 23818 -4634 24054
rect -4398 23818 -4216 24054
rect -4816 23734 -4216 23818
rect -4816 23498 -4634 23734
rect -4398 23498 -4216 23734
rect -4816 -3166 -4216 23498
rect -3876 706718 -3276 706740
rect -3876 706482 -3694 706718
rect -3458 706482 -3276 706718
rect -3876 706398 -3276 706482
rect -3876 706162 -3694 706398
rect -3458 706162 -3276 706398
rect -3876 690054 -3276 706162
rect 4404 706718 5004 707680
rect 4404 706482 4586 706718
rect 4822 706482 5004 706718
rect 4404 706398 5004 706482
rect 4404 706162 4586 706398
rect 4822 706162 5004 706398
rect -3876 689818 -3694 690054
rect -3458 689818 -3276 690054
rect -3876 689734 -3276 689818
rect -3876 689498 -3694 689734
rect -3458 689498 -3276 689734
rect -3876 654054 -3276 689498
rect -3876 653818 -3694 654054
rect -3458 653818 -3276 654054
rect -3876 653734 -3276 653818
rect -3876 653498 -3694 653734
rect -3458 653498 -3276 653734
rect -3876 618054 -3276 653498
rect -3876 617818 -3694 618054
rect -3458 617818 -3276 618054
rect -3876 617734 -3276 617818
rect -3876 617498 -3694 617734
rect -3458 617498 -3276 617734
rect -3876 582054 -3276 617498
rect -3876 581818 -3694 582054
rect -3458 581818 -3276 582054
rect -3876 581734 -3276 581818
rect -3876 581498 -3694 581734
rect -3458 581498 -3276 581734
rect -3876 546054 -3276 581498
rect -3876 545818 -3694 546054
rect -3458 545818 -3276 546054
rect -3876 545734 -3276 545818
rect -3876 545498 -3694 545734
rect -3458 545498 -3276 545734
rect -3876 510054 -3276 545498
rect -3876 509818 -3694 510054
rect -3458 509818 -3276 510054
rect -3876 509734 -3276 509818
rect -3876 509498 -3694 509734
rect -3458 509498 -3276 509734
rect -3876 474054 -3276 509498
rect -3876 473818 -3694 474054
rect -3458 473818 -3276 474054
rect -3876 473734 -3276 473818
rect -3876 473498 -3694 473734
rect -3458 473498 -3276 473734
rect -3876 438054 -3276 473498
rect -3876 437818 -3694 438054
rect -3458 437818 -3276 438054
rect -3876 437734 -3276 437818
rect -3876 437498 -3694 437734
rect -3458 437498 -3276 437734
rect -3876 402054 -3276 437498
rect -3876 401818 -3694 402054
rect -3458 401818 -3276 402054
rect -3876 401734 -3276 401818
rect -3876 401498 -3694 401734
rect -3458 401498 -3276 401734
rect -3876 366054 -3276 401498
rect -3876 365818 -3694 366054
rect -3458 365818 -3276 366054
rect -3876 365734 -3276 365818
rect -3876 365498 -3694 365734
rect -3458 365498 -3276 365734
rect -3876 330054 -3276 365498
rect -3876 329818 -3694 330054
rect -3458 329818 -3276 330054
rect -3876 329734 -3276 329818
rect -3876 329498 -3694 329734
rect -3458 329498 -3276 329734
rect -3876 294054 -3276 329498
rect -3876 293818 -3694 294054
rect -3458 293818 -3276 294054
rect -3876 293734 -3276 293818
rect -3876 293498 -3694 293734
rect -3458 293498 -3276 293734
rect -3876 258054 -3276 293498
rect -3876 257818 -3694 258054
rect -3458 257818 -3276 258054
rect -3876 257734 -3276 257818
rect -3876 257498 -3694 257734
rect -3458 257498 -3276 257734
rect -3876 222054 -3276 257498
rect -3876 221818 -3694 222054
rect -3458 221818 -3276 222054
rect -3876 221734 -3276 221818
rect -3876 221498 -3694 221734
rect -3458 221498 -3276 221734
rect -3876 186054 -3276 221498
rect -3876 185818 -3694 186054
rect -3458 185818 -3276 186054
rect -3876 185734 -3276 185818
rect -3876 185498 -3694 185734
rect -3458 185498 -3276 185734
rect -3876 150054 -3276 185498
rect -3876 149818 -3694 150054
rect -3458 149818 -3276 150054
rect -3876 149734 -3276 149818
rect -3876 149498 -3694 149734
rect -3458 149498 -3276 149734
rect -3876 114054 -3276 149498
rect -3876 113818 -3694 114054
rect -3458 113818 -3276 114054
rect -3876 113734 -3276 113818
rect -3876 113498 -3694 113734
rect -3458 113498 -3276 113734
rect -3876 78054 -3276 113498
rect -3876 77818 -3694 78054
rect -3458 77818 -3276 78054
rect -3876 77734 -3276 77818
rect -3876 77498 -3694 77734
rect -3458 77498 -3276 77734
rect -3876 42054 -3276 77498
rect -3876 41818 -3694 42054
rect -3458 41818 -3276 42054
rect -3876 41734 -3276 41818
rect -3876 41498 -3694 41734
rect -3458 41498 -3276 41734
rect -3876 6054 -3276 41498
rect -3876 5818 -3694 6054
rect -3458 5818 -3276 6054
rect -3876 5734 -3276 5818
rect -3876 5498 -3694 5734
rect -3458 5498 -3276 5734
rect -3876 -2226 -3276 5498
rect -2936 705778 -2336 705800
rect -2936 705542 -2754 705778
rect -2518 705542 -2336 705778
rect -2936 705458 -2336 705542
rect -2936 705222 -2754 705458
rect -2518 705222 -2336 705458
rect -2936 668454 -2336 705222
rect -2936 668218 -2754 668454
rect -2518 668218 -2336 668454
rect -2936 668134 -2336 668218
rect -2936 667898 -2754 668134
rect -2518 667898 -2336 668134
rect -2936 632454 -2336 667898
rect -2936 632218 -2754 632454
rect -2518 632218 -2336 632454
rect -2936 632134 -2336 632218
rect -2936 631898 -2754 632134
rect -2518 631898 -2336 632134
rect -2936 596454 -2336 631898
rect -2936 596218 -2754 596454
rect -2518 596218 -2336 596454
rect -2936 596134 -2336 596218
rect -2936 595898 -2754 596134
rect -2518 595898 -2336 596134
rect -2936 560454 -2336 595898
rect -2936 560218 -2754 560454
rect -2518 560218 -2336 560454
rect -2936 560134 -2336 560218
rect -2936 559898 -2754 560134
rect -2518 559898 -2336 560134
rect -2936 524454 -2336 559898
rect -2936 524218 -2754 524454
rect -2518 524218 -2336 524454
rect -2936 524134 -2336 524218
rect -2936 523898 -2754 524134
rect -2518 523898 -2336 524134
rect -2936 488454 -2336 523898
rect -2936 488218 -2754 488454
rect -2518 488218 -2336 488454
rect -2936 488134 -2336 488218
rect -2936 487898 -2754 488134
rect -2518 487898 -2336 488134
rect -2936 452454 -2336 487898
rect -2936 452218 -2754 452454
rect -2518 452218 -2336 452454
rect -2936 452134 -2336 452218
rect -2936 451898 -2754 452134
rect -2518 451898 -2336 452134
rect -2936 416454 -2336 451898
rect -2936 416218 -2754 416454
rect -2518 416218 -2336 416454
rect -2936 416134 -2336 416218
rect -2936 415898 -2754 416134
rect -2518 415898 -2336 416134
rect -2936 380454 -2336 415898
rect -2936 380218 -2754 380454
rect -2518 380218 -2336 380454
rect -2936 380134 -2336 380218
rect -2936 379898 -2754 380134
rect -2518 379898 -2336 380134
rect -2936 344454 -2336 379898
rect -2936 344218 -2754 344454
rect -2518 344218 -2336 344454
rect -2936 344134 -2336 344218
rect -2936 343898 -2754 344134
rect -2518 343898 -2336 344134
rect -2936 308454 -2336 343898
rect -2936 308218 -2754 308454
rect -2518 308218 -2336 308454
rect -2936 308134 -2336 308218
rect -2936 307898 -2754 308134
rect -2518 307898 -2336 308134
rect -2936 272454 -2336 307898
rect -2936 272218 -2754 272454
rect -2518 272218 -2336 272454
rect -2936 272134 -2336 272218
rect -2936 271898 -2754 272134
rect -2518 271898 -2336 272134
rect -2936 236454 -2336 271898
rect -2936 236218 -2754 236454
rect -2518 236218 -2336 236454
rect -2936 236134 -2336 236218
rect -2936 235898 -2754 236134
rect -2518 235898 -2336 236134
rect -2936 200454 -2336 235898
rect -2936 200218 -2754 200454
rect -2518 200218 -2336 200454
rect -2936 200134 -2336 200218
rect -2936 199898 -2754 200134
rect -2518 199898 -2336 200134
rect -2936 164454 -2336 199898
rect -2936 164218 -2754 164454
rect -2518 164218 -2336 164454
rect -2936 164134 -2336 164218
rect -2936 163898 -2754 164134
rect -2518 163898 -2336 164134
rect -2936 128454 -2336 163898
rect -2936 128218 -2754 128454
rect -2518 128218 -2336 128454
rect -2936 128134 -2336 128218
rect -2936 127898 -2754 128134
rect -2518 127898 -2336 128134
rect -2936 92454 -2336 127898
rect -2936 92218 -2754 92454
rect -2518 92218 -2336 92454
rect -2936 92134 -2336 92218
rect -2936 91898 -2754 92134
rect -2518 91898 -2336 92134
rect -2936 56454 -2336 91898
rect -2936 56218 -2754 56454
rect -2518 56218 -2336 56454
rect -2936 56134 -2336 56218
rect -2936 55898 -2754 56134
rect -2518 55898 -2336 56134
rect -2936 20454 -2336 55898
rect -2936 20218 -2754 20454
rect -2518 20218 -2336 20454
rect -2936 20134 -2336 20218
rect -2936 19898 -2754 20134
rect -2518 19898 -2336 20134
rect -2936 -1286 -2336 19898
rect -1996 704838 -1396 704860
rect -1996 704602 -1814 704838
rect -1578 704602 -1396 704838
rect -1996 704518 -1396 704602
rect -1996 704282 -1814 704518
rect -1578 704282 -1396 704518
rect -1996 686454 -1396 704282
rect -1996 686218 -1814 686454
rect -1578 686218 -1396 686454
rect -1996 686134 -1396 686218
rect -1996 685898 -1814 686134
rect -1578 685898 -1396 686134
rect -1996 650454 -1396 685898
rect -1996 650218 -1814 650454
rect -1578 650218 -1396 650454
rect -1996 650134 -1396 650218
rect -1996 649898 -1814 650134
rect -1578 649898 -1396 650134
rect -1996 614454 -1396 649898
rect -1996 614218 -1814 614454
rect -1578 614218 -1396 614454
rect -1996 614134 -1396 614218
rect -1996 613898 -1814 614134
rect -1578 613898 -1396 614134
rect -1996 578454 -1396 613898
rect -1996 578218 -1814 578454
rect -1578 578218 -1396 578454
rect -1996 578134 -1396 578218
rect -1996 577898 -1814 578134
rect -1578 577898 -1396 578134
rect -1996 542454 -1396 577898
rect -1996 542218 -1814 542454
rect -1578 542218 -1396 542454
rect -1996 542134 -1396 542218
rect -1996 541898 -1814 542134
rect -1578 541898 -1396 542134
rect -1996 506454 -1396 541898
rect -1996 506218 -1814 506454
rect -1578 506218 -1396 506454
rect -1996 506134 -1396 506218
rect -1996 505898 -1814 506134
rect -1578 505898 -1396 506134
rect -1996 470454 -1396 505898
rect -1996 470218 -1814 470454
rect -1578 470218 -1396 470454
rect -1996 470134 -1396 470218
rect -1996 469898 -1814 470134
rect -1578 469898 -1396 470134
rect -1996 434454 -1396 469898
rect -1996 434218 -1814 434454
rect -1578 434218 -1396 434454
rect -1996 434134 -1396 434218
rect -1996 433898 -1814 434134
rect -1578 433898 -1396 434134
rect -1996 398454 -1396 433898
rect -1996 398218 -1814 398454
rect -1578 398218 -1396 398454
rect -1996 398134 -1396 398218
rect -1996 397898 -1814 398134
rect -1578 397898 -1396 398134
rect -1996 362454 -1396 397898
rect -1996 362218 -1814 362454
rect -1578 362218 -1396 362454
rect -1996 362134 -1396 362218
rect -1996 361898 -1814 362134
rect -1578 361898 -1396 362134
rect -1996 326454 -1396 361898
rect -1996 326218 -1814 326454
rect -1578 326218 -1396 326454
rect -1996 326134 -1396 326218
rect -1996 325898 -1814 326134
rect -1578 325898 -1396 326134
rect -1996 290454 -1396 325898
rect -1996 290218 -1814 290454
rect -1578 290218 -1396 290454
rect -1996 290134 -1396 290218
rect -1996 289898 -1814 290134
rect -1578 289898 -1396 290134
rect -1996 254454 -1396 289898
rect -1996 254218 -1814 254454
rect -1578 254218 -1396 254454
rect -1996 254134 -1396 254218
rect -1996 253898 -1814 254134
rect -1578 253898 -1396 254134
rect -1996 218454 -1396 253898
rect -1996 218218 -1814 218454
rect -1578 218218 -1396 218454
rect -1996 218134 -1396 218218
rect -1996 217898 -1814 218134
rect -1578 217898 -1396 218134
rect -1996 182454 -1396 217898
rect -1996 182218 -1814 182454
rect -1578 182218 -1396 182454
rect -1996 182134 -1396 182218
rect -1996 181898 -1814 182134
rect -1578 181898 -1396 182134
rect -1996 146454 -1396 181898
rect -1996 146218 -1814 146454
rect -1578 146218 -1396 146454
rect -1996 146134 -1396 146218
rect -1996 145898 -1814 146134
rect -1578 145898 -1396 146134
rect -1996 110454 -1396 145898
rect -1996 110218 -1814 110454
rect -1578 110218 -1396 110454
rect -1996 110134 -1396 110218
rect -1996 109898 -1814 110134
rect -1578 109898 -1396 110134
rect -1996 74454 -1396 109898
rect -1996 74218 -1814 74454
rect -1578 74218 -1396 74454
rect -1996 74134 -1396 74218
rect -1996 73898 -1814 74134
rect -1578 73898 -1396 74134
rect -1996 38454 -1396 73898
rect -1996 38218 -1814 38454
rect -1578 38218 -1396 38454
rect -1996 38134 -1396 38218
rect -1996 37898 -1814 38134
rect -1578 37898 -1396 38134
rect -1996 2454 -1396 37898
rect -1996 2218 -1814 2454
rect -1578 2218 -1396 2454
rect -1996 2134 -1396 2218
rect -1996 1898 -1814 2134
rect -1578 1898 -1396 2134
rect -1996 -346 -1396 1898
rect -1996 -582 -1814 -346
rect -1578 -582 -1396 -346
rect -1996 -666 -1396 -582
rect -1996 -902 -1814 -666
rect -1578 -902 -1396 -666
rect -1996 -924 -1396 -902
rect 804 704838 1404 705800
rect 804 704602 986 704838
rect 1222 704602 1404 704838
rect 804 704518 1404 704602
rect 804 704282 986 704518
rect 1222 704282 1404 704518
rect 804 686454 1404 704282
rect 804 686218 986 686454
rect 1222 686218 1404 686454
rect 804 686134 1404 686218
rect 804 685898 986 686134
rect 1222 685898 1404 686134
rect 804 650454 1404 685898
rect 804 650218 986 650454
rect 1222 650218 1404 650454
rect 804 650134 1404 650218
rect 804 649898 986 650134
rect 1222 649898 1404 650134
rect 804 614454 1404 649898
rect 804 614218 986 614454
rect 1222 614218 1404 614454
rect 804 614134 1404 614218
rect 804 613898 986 614134
rect 1222 613898 1404 614134
rect 804 578454 1404 613898
rect 804 578218 986 578454
rect 1222 578218 1404 578454
rect 804 578134 1404 578218
rect 804 577898 986 578134
rect 1222 577898 1404 578134
rect 804 542454 1404 577898
rect 804 542218 986 542454
rect 1222 542218 1404 542454
rect 804 542134 1404 542218
rect 804 541898 986 542134
rect 1222 541898 1404 542134
rect 804 506454 1404 541898
rect 804 506218 986 506454
rect 1222 506218 1404 506454
rect 804 506134 1404 506218
rect 804 505898 986 506134
rect 1222 505898 1404 506134
rect 804 470454 1404 505898
rect 804 470218 986 470454
rect 1222 470218 1404 470454
rect 804 470134 1404 470218
rect 804 469898 986 470134
rect 1222 469898 1404 470134
rect 804 434454 1404 469898
rect 804 434218 986 434454
rect 1222 434218 1404 434454
rect 804 434134 1404 434218
rect 804 433898 986 434134
rect 1222 433898 1404 434134
rect 804 398454 1404 433898
rect 804 398218 986 398454
rect 1222 398218 1404 398454
rect 804 398134 1404 398218
rect 804 397898 986 398134
rect 1222 397898 1404 398134
rect 804 362454 1404 397898
rect 804 362218 986 362454
rect 1222 362218 1404 362454
rect 804 362134 1404 362218
rect 804 361898 986 362134
rect 1222 361898 1404 362134
rect 804 326454 1404 361898
rect 804 326218 986 326454
rect 1222 326218 1404 326454
rect 804 326134 1404 326218
rect 804 325898 986 326134
rect 1222 325898 1404 326134
rect 804 290454 1404 325898
rect 804 290218 986 290454
rect 1222 290218 1404 290454
rect 804 290134 1404 290218
rect 804 289898 986 290134
rect 1222 289898 1404 290134
rect 804 254454 1404 289898
rect 804 254218 986 254454
rect 1222 254218 1404 254454
rect 804 254134 1404 254218
rect 804 253898 986 254134
rect 1222 253898 1404 254134
rect 804 218454 1404 253898
rect 804 218218 986 218454
rect 1222 218218 1404 218454
rect 804 218134 1404 218218
rect 804 217898 986 218134
rect 1222 217898 1404 218134
rect 804 182454 1404 217898
rect 804 182218 986 182454
rect 1222 182218 1404 182454
rect 804 182134 1404 182218
rect 804 181898 986 182134
rect 1222 181898 1404 182134
rect 804 146454 1404 181898
rect 804 146218 986 146454
rect 1222 146218 1404 146454
rect 804 146134 1404 146218
rect 804 145898 986 146134
rect 1222 145898 1404 146134
rect 804 110454 1404 145898
rect 804 110218 986 110454
rect 1222 110218 1404 110454
rect 804 110134 1404 110218
rect 804 109898 986 110134
rect 1222 109898 1404 110134
rect 804 74454 1404 109898
rect 804 74218 986 74454
rect 1222 74218 1404 74454
rect 804 74134 1404 74218
rect 804 73898 986 74134
rect 1222 73898 1404 74134
rect 804 38454 1404 73898
rect 804 38218 986 38454
rect 1222 38218 1404 38454
rect 804 38134 1404 38218
rect 804 37898 986 38134
rect 1222 37898 1404 38134
rect 804 2454 1404 37898
rect 804 2218 986 2454
rect 1222 2218 1404 2454
rect 804 2134 1404 2218
rect 804 1898 986 2134
rect 1222 1898 1404 2134
rect 804 -346 1404 1898
rect 804 -582 986 -346
rect 1222 -582 1404 -346
rect 804 -666 1404 -582
rect 804 -902 986 -666
rect 1222 -902 1404 -666
rect -2936 -1522 -2754 -1286
rect -2518 -1522 -2336 -1286
rect -2936 -1606 -2336 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 -2336 -1606
rect -2936 -1864 -2336 -1842
rect 804 -1864 1404 -902
rect 4404 690054 5004 706162
rect 4404 689818 4586 690054
rect 4822 689818 5004 690054
rect 4404 689734 5004 689818
rect 4404 689498 4586 689734
rect 4822 689498 5004 689734
rect 4404 654054 5004 689498
rect 4404 653818 4586 654054
rect 4822 653818 5004 654054
rect 4404 653734 5004 653818
rect 4404 653498 4586 653734
rect 4822 653498 5004 653734
rect 4404 618054 5004 653498
rect 4404 617818 4586 618054
rect 4822 617818 5004 618054
rect 4404 617734 5004 617818
rect 4404 617498 4586 617734
rect 4822 617498 5004 617734
rect 4404 582054 5004 617498
rect 4404 581818 4586 582054
rect 4822 581818 5004 582054
rect 4404 581734 5004 581818
rect 4404 581498 4586 581734
rect 4822 581498 5004 581734
rect 4404 546054 5004 581498
rect 4404 545818 4586 546054
rect 4822 545818 5004 546054
rect 4404 545734 5004 545818
rect 4404 545498 4586 545734
rect 4822 545498 5004 545734
rect 4404 510054 5004 545498
rect 4404 509818 4586 510054
rect 4822 509818 5004 510054
rect 4404 509734 5004 509818
rect 4404 509498 4586 509734
rect 4822 509498 5004 509734
rect 4404 474054 5004 509498
rect 4404 473818 4586 474054
rect 4822 473818 5004 474054
rect 4404 473734 5004 473818
rect 4404 473498 4586 473734
rect 4822 473498 5004 473734
rect 4404 438054 5004 473498
rect 4404 437818 4586 438054
rect 4822 437818 5004 438054
rect 4404 437734 5004 437818
rect 4404 437498 4586 437734
rect 4822 437498 5004 437734
rect 4404 402054 5004 437498
rect 4404 401818 4586 402054
rect 4822 401818 5004 402054
rect 4404 401734 5004 401818
rect 4404 401498 4586 401734
rect 4822 401498 5004 401734
rect 4404 366054 5004 401498
rect 4404 365818 4586 366054
rect 4822 365818 5004 366054
rect 4404 365734 5004 365818
rect 4404 365498 4586 365734
rect 4822 365498 5004 365734
rect 4404 330054 5004 365498
rect 4404 329818 4586 330054
rect 4822 329818 5004 330054
rect 4404 329734 5004 329818
rect 4404 329498 4586 329734
rect 4822 329498 5004 329734
rect 4404 294054 5004 329498
rect 4404 293818 4586 294054
rect 4822 293818 5004 294054
rect 4404 293734 5004 293818
rect 4404 293498 4586 293734
rect 4822 293498 5004 293734
rect 4404 258054 5004 293498
rect 4404 257818 4586 258054
rect 4822 257818 5004 258054
rect 4404 257734 5004 257818
rect 4404 257498 4586 257734
rect 4822 257498 5004 257734
rect 4404 222054 5004 257498
rect 4404 221818 4586 222054
rect 4822 221818 5004 222054
rect 4404 221734 5004 221818
rect 4404 221498 4586 221734
rect 4822 221498 5004 221734
rect 4404 186054 5004 221498
rect 4404 185818 4586 186054
rect 4822 185818 5004 186054
rect 4404 185734 5004 185818
rect 4404 185498 4586 185734
rect 4822 185498 5004 185734
rect 4404 150054 5004 185498
rect 4404 149818 4586 150054
rect 4822 149818 5004 150054
rect 4404 149734 5004 149818
rect 4404 149498 4586 149734
rect 4822 149498 5004 149734
rect 4404 114054 5004 149498
rect 4404 113818 4586 114054
rect 4822 113818 5004 114054
rect 4404 113734 5004 113818
rect 4404 113498 4586 113734
rect 4822 113498 5004 113734
rect 4404 78054 5004 113498
rect 4404 77818 4586 78054
rect 4822 77818 5004 78054
rect 4404 77734 5004 77818
rect 4404 77498 4586 77734
rect 4822 77498 5004 77734
rect 4404 42054 5004 77498
rect 4404 41818 4586 42054
rect 4822 41818 5004 42054
rect 4404 41734 5004 41818
rect 4404 41498 4586 41734
rect 4822 41498 5004 41734
rect 4404 6054 5004 41498
rect 4404 5818 4586 6054
rect 4822 5818 5004 6054
rect 4404 5734 5004 5818
rect 4404 5498 4586 5734
rect 4822 5498 5004 5734
rect -3876 -2462 -3694 -2226
rect -3458 -2462 -3276 -2226
rect -3876 -2546 -3276 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 -3276 -2546
rect -3876 -2804 -3276 -2782
rect 4404 -2226 5004 5498
rect 4404 -2462 4586 -2226
rect 4822 -2462 5004 -2226
rect 4404 -2546 5004 -2462
rect 4404 -2782 4586 -2546
rect 4822 -2782 5004 -2546
rect -4816 -3402 -4634 -3166
rect -4398 -3402 -4216 -3166
rect -4816 -3486 -4216 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 -4216 -3486
rect -4816 -3744 -4216 -3722
rect 4404 -3744 5004 -2782
rect 8004 693654 8604 708042
rect 8004 693418 8186 693654
rect 8422 693418 8604 693654
rect 8004 693334 8604 693418
rect 8004 693098 8186 693334
rect 8422 693098 8604 693334
rect 8004 657654 8604 693098
rect 8004 657418 8186 657654
rect 8422 657418 8604 657654
rect 8004 657334 8604 657418
rect 8004 657098 8186 657334
rect 8422 657098 8604 657334
rect 8004 621654 8604 657098
rect 8004 621418 8186 621654
rect 8422 621418 8604 621654
rect 8004 621334 8604 621418
rect 8004 621098 8186 621334
rect 8422 621098 8604 621334
rect 8004 585654 8604 621098
rect 8004 585418 8186 585654
rect 8422 585418 8604 585654
rect 8004 585334 8604 585418
rect 8004 585098 8186 585334
rect 8422 585098 8604 585334
rect 8004 549654 8604 585098
rect 8004 549418 8186 549654
rect 8422 549418 8604 549654
rect 8004 549334 8604 549418
rect 8004 549098 8186 549334
rect 8422 549098 8604 549334
rect 8004 513654 8604 549098
rect 8004 513418 8186 513654
rect 8422 513418 8604 513654
rect 8004 513334 8604 513418
rect 8004 513098 8186 513334
rect 8422 513098 8604 513334
rect 8004 477654 8604 513098
rect 8004 477418 8186 477654
rect 8422 477418 8604 477654
rect 8004 477334 8604 477418
rect 8004 477098 8186 477334
rect 8422 477098 8604 477334
rect 8004 441654 8604 477098
rect 8004 441418 8186 441654
rect 8422 441418 8604 441654
rect 8004 441334 8604 441418
rect 8004 441098 8186 441334
rect 8422 441098 8604 441334
rect 8004 405654 8604 441098
rect 8004 405418 8186 405654
rect 8422 405418 8604 405654
rect 8004 405334 8604 405418
rect 8004 405098 8186 405334
rect 8422 405098 8604 405334
rect 8004 369654 8604 405098
rect 8004 369418 8186 369654
rect 8422 369418 8604 369654
rect 8004 369334 8604 369418
rect 8004 369098 8186 369334
rect 8422 369098 8604 369334
rect 8004 333654 8604 369098
rect 8004 333418 8186 333654
rect 8422 333418 8604 333654
rect 8004 333334 8604 333418
rect 8004 333098 8186 333334
rect 8422 333098 8604 333334
rect 8004 297654 8604 333098
rect 8004 297418 8186 297654
rect 8422 297418 8604 297654
rect 8004 297334 8604 297418
rect 8004 297098 8186 297334
rect 8422 297098 8604 297334
rect 8004 261654 8604 297098
rect 8004 261418 8186 261654
rect 8422 261418 8604 261654
rect 8004 261334 8604 261418
rect 8004 261098 8186 261334
rect 8422 261098 8604 261334
rect 8004 225654 8604 261098
rect 8004 225418 8186 225654
rect 8422 225418 8604 225654
rect 8004 225334 8604 225418
rect 8004 225098 8186 225334
rect 8422 225098 8604 225334
rect 8004 189654 8604 225098
rect 8004 189418 8186 189654
rect 8422 189418 8604 189654
rect 8004 189334 8604 189418
rect 8004 189098 8186 189334
rect 8422 189098 8604 189334
rect 8004 153654 8604 189098
rect 8004 153418 8186 153654
rect 8422 153418 8604 153654
rect 8004 153334 8604 153418
rect 8004 153098 8186 153334
rect 8422 153098 8604 153334
rect 8004 117654 8604 153098
rect 8004 117418 8186 117654
rect 8422 117418 8604 117654
rect 8004 117334 8604 117418
rect 8004 117098 8186 117334
rect 8422 117098 8604 117334
rect 8004 81654 8604 117098
rect 8004 81418 8186 81654
rect 8422 81418 8604 81654
rect 8004 81334 8604 81418
rect 8004 81098 8186 81334
rect 8422 81098 8604 81334
rect 8004 45654 8604 81098
rect 8004 45418 8186 45654
rect 8422 45418 8604 45654
rect 8004 45334 8604 45418
rect 8004 45098 8186 45334
rect 8422 45098 8604 45334
rect 8004 9654 8604 45098
rect 8004 9418 8186 9654
rect 8422 9418 8604 9654
rect 8004 9334 8604 9418
rect 8004 9098 8186 9334
rect 8422 9098 8604 9334
rect -5756 -4342 -5574 -4106
rect -5338 -4342 -5156 -4106
rect -5756 -4426 -5156 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 -5156 -4426
rect -5756 -4684 -5156 -4662
rect 8004 -4106 8604 9098
rect 8004 -4342 8186 -4106
rect 8422 -4342 8604 -4106
rect 8004 -4426 8604 -4342
rect 8004 -4662 8186 -4426
rect 8422 -4662 8604 -4426
rect -6696 -5282 -6514 -5046
rect -6278 -5282 -6096 -5046
rect -6696 -5366 -6096 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 -6096 -5366
rect -6696 -5624 -6096 -5602
rect 8004 -5624 8604 -4662
rect 11604 697254 12204 709922
rect 29604 711418 30204 711440
rect 29604 711182 29786 711418
rect 30022 711182 30204 711418
rect 29604 711098 30204 711182
rect 29604 710862 29786 711098
rect 30022 710862 30204 711098
rect 26004 709538 26604 709560
rect 26004 709302 26186 709538
rect 26422 709302 26604 709538
rect 26004 709218 26604 709302
rect 26004 708982 26186 709218
rect 26422 708982 26604 709218
rect 22404 707658 23004 707680
rect 22404 707422 22586 707658
rect 22822 707422 23004 707658
rect 22404 707338 23004 707422
rect 22404 707102 22586 707338
rect 22822 707102 23004 707338
rect 11604 697018 11786 697254
rect 12022 697018 12204 697254
rect 11604 696934 12204 697018
rect 11604 696698 11786 696934
rect 12022 696698 12204 696934
rect 11604 661254 12204 696698
rect 11604 661018 11786 661254
rect 12022 661018 12204 661254
rect 11604 660934 12204 661018
rect 11604 660698 11786 660934
rect 12022 660698 12204 660934
rect 11604 625254 12204 660698
rect 11604 625018 11786 625254
rect 12022 625018 12204 625254
rect 11604 624934 12204 625018
rect 11604 624698 11786 624934
rect 12022 624698 12204 624934
rect 11604 589254 12204 624698
rect 11604 589018 11786 589254
rect 12022 589018 12204 589254
rect 11604 588934 12204 589018
rect 11604 588698 11786 588934
rect 12022 588698 12204 588934
rect 11604 553254 12204 588698
rect 11604 553018 11786 553254
rect 12022 553018 12204 553254
rect 11604 552934 12204 553018
rect 11604 552698 11786 552934
rect 12022 552698 12204 552934
rect 11604 517254 12204 552698
rect 11604 517018 11786 517254
rect 12022 517018 12204 517254
rect 11604 516934 12204 517018
rect 11604 516698 11786 516934
rect 12022 516698 12204 516934
rect 11604 481254 12204 516698
rect 11604 481018 11786 481254
rect 12022 481018 12204 481254
rect 11604 480934 12204 481018
rect 11604 480698 11786 480934
rect 12022 480698 12204 480934
rect 11604 445254 12204 480698
rect 11604 445018 11786 445254
rect 12022 445018 12204 445254
rect 11604 444934 12204 445018
rect 11604 444698 11786 444934
rect 12022 444698 12204 444934
rect 11604 409254 12204 444698
rect 11604 409018 11786 409254
rect 12022 409018 12204 409254
rect 11604 408934 12204 409018
rect 11604 408698 11786 408934
rect 12022 408698 12204 408934
rect 11604 373254 12204 408698
rect 11604 373018 11786 373254
rect 12022 373018 12204 373254
rect 11604 372934 12204 373018
rect 11604 372698 11786 372934
rect 12022 372698 12204 372934
rect 11604 337254 12204 372698
rect 11604 337018 11786 337254
rect 12022 337018 12204 337254
rect 11604 336934 12204 337018
rect 11604 336698 11786 336934
rect 12022 336698 12204 336934
rect 11604 301254 12204 336698
rect 11604 301018 11786 301254
rect 12022 301018 12204 301254
rect 11604 300934 12204 301018
rect 11604 300698 11786 300934
rect 12022 300698 12204 300934
rect 11604 265254 12204 300698
rect 11604 265018 11786 265254
rect 12022 265018 12204 265254
rect 11604 264934 12204 265018
rect 11604 264698 11786 264934
rect 12022 264698 12204 264934
rect 11604 229254 12204 264698
rect 11604 229018 11786 229254
rect 12022 229018 12204 229254
rect 11604 228934 12204 229018
rect 11604 228698 11786 228934
rect 12022 228698 12204 228934
rect 11604 193254 12204 228698
rect 11604 193018 11786 193254
rect 12022 193018 12204 193254
rect 11604 192934 12204 193018
rect 11604 192698 11786 192934
rect 12022 192698 12204 192934
rect 11604 157254 12204 192698
rect 11604 157018 11786 157254
rect 12022 157018 12204 157254
rect 11604 156934 12204 157018
rect 11604 156698 11786 156934
rect 12022 156698 12204 156934
rect 11604 121254 12204 156698
rect 11604 121018 11786 121254
rect 12022 121018 12204 121254
rect 11604 120934 12204 121018
rect 11604 120698 11786 120934
rect 12022 120698 12204 120934
rect 11604 85254 12204 120698
rect 11604 85018 11786 85254
rect 12022 85018 12204 85254
rect 11604 84934 12204 85018
rect 11604 84698 11786 84934
rect 12022 84698 12204 84934
rect 11604 49254 12204 84698
rect 11604 49018 11786 49254
rect 12022 49018 12204 49254
rect 11604 48934 12204 49018
rect 11604 48698 11786 48934
rect 12022 48698 12204 48934
rect 11604 13254 12204 48698
rect 11604 13018 11786 13254
rect 12022 13018 12204 13254
rect 11604 12934 12204 13018
rect 11604 12698 11786 12934
rect 12022 12698 12204 12934
rect -7636 -6222 -7454 -5986
rect -7218 -6222 -7036 -5986
rect -7636 -6306 -7036 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 -7036 -6306
rect -7636 -6564 -7036 -6542
rect 11604 -5986 12204 12698
rect 18804 705778 19404 705800
rect 18804 705542 18986 705778
rect 19222 705542 19404 705778
rect 18804 705458 19404 705542
rect 18804 705222 18986 705458
rect 19222 705222 19404 705458
rect 18804 668454 19404 705222
rect 18804 668218 18986 668454
rect 19222 668218 19404 668454
rect 18804 668134 19404 668218
rect 18804 667898 18986 668134
rect 19222 667898 19404 668134
rect 18804 632454 19404 667898
rect 18804 632218 18986 632454
rect 19222 632218 19404 632454
rect 18804 632134 19404 632218
rect 18804 631898 18986 632134
rect 19222 631898 19404 632134
rect 18804 596454 19404 631898
rect 18804 596218 18986 596454
rect 19222 596218 19404 596454
rect 18804 596134 19404 596218
rect 18804 595898 18986 596134
rect 19222 595898 19404 596134
rect 18804 560454 19404 595898
rect 18804 560218 18986 560454
rect 19222 560218 19404 560454
rect 18804 560134 19404 560218
rect 18804 559898 18986 560134
rect 19222 559898 19404 560134
rect 18804 524454 19404 559898
rect 18804 524218 18986 524454
rect 19222 524218 19404 524454
rect 18804 524134 19404 524218
rect 18804 523898 18986 524134
rect 19222 523898 19404 524134
rect 18804 488454 19404 523898
rect 18804 488218 18986 488454
rect 19222 488218 19404 488454
rect 18804 488134 19404 488218
rect 18804 487898 18986 488134
rect 19222 487898 19404 488134
rect 18804 452454 19404 487898
rect 18804 452218 18986 452454
rect 19222 452218 19404 452454
rect 18804 452134 19404 452218
rect 18804 451898 18986 452134
rect 19222 451898 19404 452134
rect 18804 416454 19404 451898
rect 18804 416218 18986 416454
rect 19222 416218 19404 416454
rect 18804 416134 19404 416218
rect 18804 415898 18986 416134
rect 19222 415898 19404 416134
rect 18804 380454 19404 415898
rect 18804 380218 18986 380454
rect 19222 380218 19404 380454
rect 18804 380134 19404 380218
rect 18804 379898 18986 380134
rect 19222 379898 19404 380134
rect 18804 344454 19404 379898
rect 18804 344218 18986 344454
rect 19222 344218 19404 344454
rect 18804 344134 19404 344218
rect 18804 343898 18986 344134
rect 19222 343898 19404 344134
rect 18804 308454 19404 343898
rect 18804 308218 18986 308454
rect 19222 308218 19404 308454
rect 18804 308134 19404 308218
rect 18804 307898 18986 308134
rect 19222 307898 19404 308134
rect 18804 272454 19404 307898
rect 18804 272218 18986 272454
rect 19222 272218 19404 272454
rect 18804 272134 19404 272218
rect 18804 271898 18986 272134
rect 19222 271898 19404 272134
rect 18804 236454 19404 271898
rect 18804 236218 18986 236454
rect 19222 236218 19404 236454
rect 18804 236134 19404 236218
rect 18804 235898 18986 236134
rect 19222 235898 19404 236134
rect 18804 200454 19404 235898
rect 18804 200218 18986 200454
rect 19222 200218 19404 200454
rect 18804 200134 19404 200218
rect 18804 199898 18986 200134
rect 19222 199898 19404 200134
rect 18804 164454 19404 199898
rect 18804 164218 18986 164454
rect 19222 164218 19404 164454
rect 18804 164134 19404 164218
rect 18804 163898 18986 164134
rect 19222 163898 19404 164134
rect 18804 128454 19404 163898
rect 18804 128218 18986 128454
rect 19222 128218 19404 128454
rect 18804 128134 19404 128218
rect 18804 127898 18986 128134
rect 19222 127898 19404 128134
rect 18804 92454 19404 127898
rect 18804 92218 18986 92454
rect 19222 92218 19404 92454
rect 18804 92134 19404 92218
rect 18804 91898 18986 92134
rect 19222 91898 19404 92134
rect 18804 56454 19404 91898
rect 18804 56218 18986 56454
rect 19222 56218 19404 56454
rect 18804 56134 19404 56218
rect 18804 55898 18986 56134
rect 19222 55898 19404 56134
rect 18804 20454 19404 55898
rect 18804 20218 18986 20454
rect 19222 20218 19404 20454
rect 18804 20134 19404 20218
rect 18804 19898 18986 20134
rect 19222 19898 19404 20134
rect 18804 -1286 19404 19898
rect 18804 -1522 18986 -1286
rect 19222 -1522 19404 -1286
rect 18804 -1606 19404 -1522
rect 18804 -1842 18986 -1606
rect 19222 -1842 19404 -1606
rect 18804 -1864 19404 -1842
rect 22404 672054 23004 707102
rect 22404 671818 22586 672054
rect 22822 671818 23004 672054
rect 22404 671734 23004 671818
rect 22404 671498 22586 671734
rect 22822 671498 23004 671734
rect 22404 636054 23004 671498
rect 22404 635818 22586 636054
rect 22822 635818 23004 636054
rect 22404 635734 23004 635818
rect 22404 635498 22586 635734
rect 22822 635498 23004 635734
rect 22404 600054 23004 635498
rect 22404 599818 22586 600054
rect 22822 599818 23004 600054
rect 22404 599734 23004 599818
rect 22404 599498 22586 599734
rect 22822 599498 23004 599734
rect 22404 564054 23004 599498
rect 22404 563818 22586 564054
rect 22822 563818 23004 564054
rect 22404 563734 23004 563818
rect 22404 563498 22586 563734
rect 22822 563498 23004 563734
rect 22404 528054 23004 563498
rect 22404 527818 22586 528054
rect 22822 527818 23004 528054
rect 22404 527734 23004 527818
rect 22404 527498 22586 527734
rect 22822 527498 23004 527734
rect 22404 492054 23004 527498
rect 22404 491818 22586 492054
rect 22822 491818 23004 492054
rect 22404 491734 23004 491818
rect 22404 491498 22586 491734
rect 22822 491498 23004 491734
rect 22404 456054 23004 491498
rect 22404 455818 22586 456054
rect 22822 455818 23004 456054
rect 22404 455734 23004 455818
rect 22404 455498 22586 455734
rect 22822 455498 23004 455734
rect 22404 420054 23004 455498
rect 22404 419818 22586 420054
rect 22822 419818 23004 420054
rect 22404 419734 23004 419818
rect 22404 419498 22586 419734
rect 22822 419498 23004 419734
rect 22404 384054 23004 419498
rect 22404 383818 22586 384054
rect 22822 383818 23004 384054
rect 22404 383734 23004 383818
rect 22404 383498 22586 383734
rect 22822 383498 23004 383734
rect 22404 348054 23004 383498
rect 22404 347818 22586 348054
rect 22822 347818 23004 348054
rect 22404 347734 23004 347818
rect 22404 347498 22586 347734
rect 22822 347498 23004 347734
rect 22404 312054 23004 347498
rect 22404 311818 22586 312054
rect 22822 311818 23004 312054
rect 22404 311734 23004 311818
rect 22404 311498 22586 311734
rect 22822 311498 23004 311734
rect 22404 276054 23004 311498
rect 22404 275818 22586 276054
rect 22822 275818 23004 276054
rect 22404 275734 23004 275818
rect 22404 275498 22586 275734
rect 22822 275498 23004 275734
rect 22404 240054 23004 275498
rect 22404 239818 22586 240054
rect 22822 239818 23004 240054
rect 22404 239734 23004 239818
rect 22404 239498 22586 239734
rect 22822 239498 23004 239734
rect 22404 204054 23004 239498
rect 22404 203818 22586 204054
rect 22822 203818 23004 204054
rect 22404 203734 23004 203818
rect 22404 203498 22586 203734
rect 22822 203498 23004 203734
rect 22404 168054 23004 203498
rect 22404 167818 22586 168054
rect 22822 167818 23004 168054
rect 22404 167734 23004 167818
rect 22404 167498 22586 167734
rect 22822 167498 23004 167734
rect 22404 132054 23004 167498
rect 22404 131818 22586 132054
rect 22822 131818 23004 132054
rect 22404 131734 23004 131818
rect 22404 131498 22586 131734
rect 22822 131498 23004 131734
rect 22404 96054 23004 131498
rect 22404 95818 22586 96054
rect 22822 95818 23004 96054
rect 22404 95734 23004 95818
rect 22404 95498 22586 95734
rect 22822 95498 23004 95734
rect 22404 60054 23004 95498
rect 22404 59818 22586 60054
rect 22822 59818 23004 60054
rect 22404 59734 23004 59818
rect 22404 59498 22586 59734
rect 22822 59498 23004 59734
rect 22404 24054 23004 59498
rect 22404 23818 22586 24054
rect 22822 23818 23004 24054
rect 22404 23734 23004 23818
rect 22404 23498 22586 23734
rect 22822 23498 23004 23734
rect 22404 -3166 23004 23498
rect 22404 -3402 22586 -3166
rect 22822 -3402 23004 -3166
rect 22404 -3486 23004 -3402
rect 22404 -3722 22586 -3486
rect 22822 -3722 23004 -3486
rect 22404 -3744 23004 -3722
rect 26004 675654 26604 708982
rect 26004 675418 26186 675654
rect 26422 675418 26604 675654
rect 26004 675334 26604 675418
rect 26004 675098 26186 675334
rect 26422 675098 26604 675334
rect 26004 639654 26604 675098
rect 26004 639418 26186 639654
rect 26422 639418 26604 639654
rect 26004 639334 26604 639418
rect 26004 639098 26186 639334
rect 26422 639098 26604 639334
rect 26004 603654 26604 639098
rect 26004 603418 26186 603654
rect 26422 603418 26604 603654
rect 26004 603334 26604 603418
rect 26004 603098 26186 603334
rect 26422 603098 26604 603334
rect 26004 567654 26604 603098
rect 26004 567418 26186 567654
rect 26422 567418 26604 567654
rect 26004 567334 26604 567418
rect 26004 567098 26186 567334
rect 26422 567098 26604 567334
rect 26004 531654 26604 567098
rect 26004 531418 26186 531654
rect 26422 531418 26604 531654
rect 26004 531334 26604 531418
rect 26004 531098 26186 531334
rect 26422 531098 26604 531334
rect 26004 495654 26604 531098
rect 26004 495418 26186 495654
rect 26422 495418 26604 495654
rect 26004 495334 26604 495418
rect 26004 495098 26186 495334
rect 26422 495098 26604 495334
rect 26004 459654 26604 495098
rect 26004 459418 26186 459654
rect 26422 459418 26604 459654
rect 26004 459334 26604 459418
rect 26004 459098 26186 459334
rect 26422 459098 26604 459334
rect 26004 423654 26604 459098
rect 26004 423418 26186 423654
rect 26422 423418 26604 423654
rect 26004 423334 26604 423418
rect 26004 423098 26186 423334
rect 26422 423098 26604 423334
rect 26004 387654 26604 423098
rect 26004 387418 26186 387654
rect 26422 387418 26604 387654
rect 26004 387334 26604 387418
rect 26004 387098 26186 387334
rect 26422 387098 26604 387334
rect 26004 351654 26604 387098
rect 26004 351418 26186 351654
rect 26422 351418 26604 351654
rect 26004 351334 26604 351418
rect 26004 351098 26186 351334
rect 26422 351098 26604 351334
rect 26004 315654 26604 351098
rect 26004 315418 26186 315654
rect 26422 315418 26604 315654
rect 26004 315334 26604 315418
rect 26004 315098 26186 315334
rect 26422 315098 26604 315334
rect 26004 279654 26604 315098
rect 26004 279418 26186 279654
rect 26422 279418 26604 279654
rect 26004 279334 26604 279418
rect 26004 279098 26186 279334
rect 26422 279098 26604 279334
rect 26004 243654 26604 279098
rect 26004 243418 26186 243654
rect 26422 243418 26604 243654
rect 26004 243334 26604 243418
rect 26004 243098 26186 243334
rect 26422 243098 26604 243334
rect 26004 207654 26604 243098
rect 26004 207418 26186 207654
rect 26422 207418 26604 207654
rect 26004 207334 26604 207418
rect 26004 207098 26186 207334
rect 26422 207098 26604 207334
rect 26004 171654 26604 207098
rect 26004 171418 26186 171654
rect 26422 171418 26604 171654
rect 26004 171334 26604 171418
rect 26004 171098 26186 171334
rect 26422 171098 26604 171334
rect 26004 135654 26604 171098
rect 26004 135418 26186 135654
rect 26422 135418 26604 135654
rect 26004 135334 26604 135418
rect 26004 135098 26186 135334
rect 26422 135098 26604 135334
rect 26004 99654 26604 135098
rect 26004 99418 26186 99654
rect 26422 99418 26604 99654
rect 26004 99334 26604 99418
rect 26004 99098 26186 99334
rect 26422 99098 26604 99334
rect 26004 63654 26604 99098
rect 26004 63418 26186 63654
rect 26422 63418 26604 63654
rect 26004 63334 26604 63418
rect 26004 63098 26186 63334
rect 26422 63098 26604 63334
rect 26004 27654 26604 63098
rect 26004 27418 26186 27654
rect 26422 27418 26604 27654
rect 26004 27334 26604 27418
rect 26004 27098 26186 27334
rect 26422 27098 26604 27334
rect 26004 -5046 26604 27098
rect 26004 -5282 26186 -5046
rect 26422 -5282 26604 -5046
rect 26004 -5366 26604 -5282
rect 26004 -5602 26186 -5366
rect 26422 -5602 26604 -5366
rect 26004 -5624 26604 -5602
rect 29604 679254 30204 710862
rect 47604 710478 48204 711440
rect 47604 710242 47786 710478
rect 48022 710242 48204 710478
rect 47604 710158 48204 710242
rect 47604 709922 47786 710158
rect 48022 709922 48204 710158
rect 44004 708598 44604 709560
rect 44004 708362 44186 708598
rect 44422 708362 44604 708598
rect 44004 708278 44604 708362
rect 44004 708042 44186 708278
rect 44422 708042 44604 708278
rect 40404 706718 41004 707680
rect 40404 706482 40586 706718
rect 40822 706482 41004 706718
rect 40404 706398 41004 706482
rect 40404 706162 40586 706398
rect 40822 706162 41004 706398
rect 29604 679018 29786 679254
rect 30022 679018 30204 679254
rect 29604 678934 30204 679018
rect 29604 678698 29786 678934
rect 30022 678698 30204 678934
rect 29604 643254 30204 678698
rect 29604 643018 29786 643254
rect 30022 643018 30204 643254
rect 29604 642934 30204 643018
rect 29604 642698 29786 642934
rect 30022 642698 30204 642934
rect 29604 607254 30204 642698
rect 29604 607018 29786 607254
rect 30022 607018 30204 607254
rect 29604 606934 30204 607018
rect 29604 606698 29786 606934
rect 30022 606698 30204 606934
rect 29604 571254 30204 606698
rect 29604 571018 29786 571254
rect 30022 571018 30204 571254
rect 29604 570934 30204 571018
rect 29604 570698 29786 570934
rect 30022 570698 30204 570934
rect 29604 535254 30204 570698
rect 29604 535018 29786 535254
rect 30022 535018 30204 535254
rect 29604 534934 30204 535018
rect 29604 534698 29786 534934
rect 30022 534698 30204 534934
rect 29604 499254 30204 534698
rect 29604 499018 29786 499254
rect 30022 499018 30204 499254
rect 29604 498934 30204 499018
rect 29604 498698 29786 498934
rect 30022 498698 30204 498934
rect 29604 463254 30204 498698
rect 29604 463018 29786 463254
rect 30022 463018 30204 463254
rect 29604 462934 30204 463018
rect 29604 462698 29786 462934
rect 30022 462698 30204 462934
rect 29604 427254 30204 462698
rect 29604 427018 29786 427254
rect 30022 427018 30204 427254
rect 29604 426934 30204 427018
rect 29604 426698 29786 426934
rect 30022 426698 30204 426934
rect 29604 391254 30204 426698
rect 29604 391018 29786 391254
rect 30022 391018 30204 391254
rect 29604 390934 30204 391018
rect 29604 390698 29786 390934
rect 30022 390698 30204 390934
rect 29604 355254 30204 390698
rect 29604 355018 29786 355254
rect 30022 355018 30204 355254
rect 29604 354934 30204 355018
rect 29604 354698 29786 354934
rect 30022 354698 30204 354934
rect 29604 319254 30204 354698
rect 29604 319018 29786 319254
rect 30022 319018 30204 319254
rect 29604 318934 30204 319018
rect 29604 318698 29786 318934
rect 30022 318698 30204 318934
rect 29604 283254 30204 318698
rect 29604 283018 29786 283254
rect 30022 283018 30204 283254
rect 29604 282934 30204 283018
rect 29604 282698 29786 282934
rect 30022 282698 30204 282934
rect 29604 247254 30204 282698
rect 29604 247018 29786 247254
rect 30022 247018 30204 247254
rect 29604 246934 30204 247018
rect 29604 246698 29786 246934
rect 30022 246698 30204 246934
rect 29604 211254 30204 246698
rect 29604 211018 29786 211254
rect 30022 211018 30204 211254
rect 29604 210934 30204 211018
rect 29604 210698 29786 210934
rect 30022 210698 30204 210934
rect 29604 175254 30204 210698
rect 29604 175018 29786 175254
rect 30022 175018 30204 175254
rect 29604 174934 30204 175018
rect 29604 174698 29786 174934
rect 30022 174698 30204 174934
rect 29604 139254 30204 174698
rect 29604 139018 29786 139254
rect 30022 139018 30204 139254
rect 29604 138934 30204 139018
rect 29604 138698 29786 138934
rect 30022 138698 30204 138934
rect 29604 103254 30204 138698
rect 29604 103018 29786 103254
rect 30022 103018 30204 103254
rect 29604 102934 30204 103018
rect 29604 102698 29786 102934
rect 30022 102698 30204 102934
rect 29604 67254 30204 102698
rect 29604 67018 29786 67254
rect 30022 67018 30204 67254
rect 29604 66934 30204 67018
rect 29604 66698 29786 66934
rect 30022 66698 30204 66934
rect 29604 31254 30204 66698
rect 29604 31018 29786 31254
rect 30022 31018 30204 31254
rect 29604 30934 30204 31018
rect 29604 30698 29786 30934
rect 30022 30698 30204 30934
rect 11604 -6222 11786 -5986
rect 12022 -6222 12204 -5986
rect 11604 -6306 12204 -6222
rect 11604 -6542 11786 -6306
rect 12022 -6542 12204 -6306
rect -8576 -7162 -8394 -6926
rect -8158 -7162 -7976 -6926
rect -8576 -7246 -7976 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 -7976 -7246
rect -8576 -7504 -7976 -7482
rect 11604 -7504 12204 -6542
rect 29604 -6926 30204 30698
rect 36804 704838 37404 705800
rect 36804 704602 36986 704838
rect 37222 704602 37404 704838
rect 36804 704518 37404 704602
rect 36804 704282 36986 704518
rect 37222 704282 37404 704518
rect 36804 686454 37404 704282
rect 36804 686218 36986 686454
rect 37222 686218 37404 686454
rect 36804 686134 37404 686218
rect 36804 685898 36986 686134
rect 37222 685898 37404 686134
rect 36804 650454 37404 685898
rect 36804 650218 36986 650454
rect 37222 650218 37404 650454
rect 36804 650134 37404 650218
rect 36804 649898 36986 650134
rect 37222 649898 37404 650134
rect 36804 614454 37404 649898
rect 36804 614218 36986 614454
rect 37222 614218 37404 614454
rect 36804 614134 37404 614218
rect 36804 613898 36986 614134
rect 37222 613898 37404 614134
rect 36804 578454 37404 613898
rect 36804 578218 36986 578454
rect 37222 578218 37404 578454
rect 36804 578134 37404 578218
rect 36804 577898 36986 578134
rect 37222 577898 37404 578134
rect 36804 542454 37404 577898
rect 36804 542218 36986 542454
rect 37222 542218 37404 542454
rect 36804 542134 37404 542218
rect 36804 541898 36986 542134
rect 37222 541898 37404 542134
rect 36804 506454 37404 541898
rect 36804 506218 36986 506454
rect 37222 506218 37404 506454
rect 36804 506134 37404 506218
rect 36804 505898 36986 506134
rect 37222 505898 37404 506134
rect 36804 470454 37404 505898
rect 36804 470218 36986 470454
rect 37222 470218 37404 470454
rect 36804 470134 37404 470218
rect 36804 469898 36986 470134
rect 37222 469898 37404 470134
rect 36804 434454 37404 469898
rect 36804 434218 36986 434454
rect 37222 434218 37404 434454
rect 36804 434134 37404 434218
rect 36804 433898 36986 434134
rect 37222 433898 37404 434134
rect 36804 398454 37404 433898
rect 36804 398218 36986 398454
rect 37222 398218 37404 398454
rect 36804 398134 37404 398218
rect 36804 397898 36986 398134
rect 37222 397898 37404 398134
rect 36804 362454 37404 397898
rect 36804 362218 36986 362454
rect 37222 362218 37404 362454
rect 36804 362134 37404 362218
rect 36804 361898 36986 362134
rect 37222 361898 37404 362134
rect 36804 326454 37404 361898
rect 36804 326218 36986 326454
rect 37222 326218 37404 326454
rect 36804 326134 37404 326218
rect 36804 325898 36986 326134
rect 37222 325898 37404 326134
rect 36804 290454 37404 325898
rect 36804 290218 36986 290454
rect 37222 290218 37404 290454
rect 36804 290134 37404 290218
rect 36804 289898 36986 290134
rect 37222 289898 37404 290134
rect 36804 254454 37404 289898
rect 36804 254218 36986 254454
rect 37222 254218 37404 254454
rect 36804 254134 37404 254218
rect 36804 253898 36986 254134
rect 37222 253898 37404 254134
rect 36804 218454 37404 253898
rect 36804 218218 36986 218454
rect 37222 218218 37404 218454
rect 36804 218134 37404 218218
rect 36804 217898 36986 218134
rect 37222 217898 37404 218134
rect 36804 182454 37404 217898
rect 36804 182218 36986 182454
rect 37222 182218 37404 182454
rect 36804 182134 37404 182218
rect 36804 181898 36986 182134
rect 37222 181898 37404 182134
rect 36804 146454 37404 181898
rect 36804 146218 36986 146454
rect 37222 146218 37404 146454
rect 36804 146134 37404 146218
rect 36804 145898 36986 146134
rect 37222 145898 37404 146134
rect 36804 110454 37404 145898
rect 36804 110218 36986 110454
rect 37222 110218 37404 110454
rect 36804 110134 37404 110218
rect 36804 109898 36986 110134
rect 37222 109898 37404 110134
rect 36804 74454 37404 109898
rect 36804 74218 36986 74454
rect 37222 74218 37404 74454
rect 36804 74134 37404 74218
rect 36804 73898 36986 74134
rect 37222 73898 37404 74134
rect 36804 38454 37404 73898
rect 36804 38218 36986 38454
rect 37222 38218 37404 38454
rect 36804 38134 37404 38218
rect 36804 37898 36986 38134
rect 37222 37898 37404 38134
rect 36804 2454 37404 37898
rect 36804 2218 36986 2454
rect 37222 2218 37404 2454
rect 36804 2134 37404 2218
rect 36804 1898 36986 2134
rect 37222 1898 37404 2134
rect 36804 -346 37404 1898
rect 36804 -582 36986 -346
rect 37222 -582 37404 -346
rect 36804 -666 37404 -582
rect 36804 -902 36986 -666
rect 37222 -902 37404 -666
rect 36804 -1864 37404 -902
rect 40404 690054 41004 706162
rect 40404 689818 40586 690054
rect 40822 689818 41004 690054
rect 40404 689734 41004 689818
rect 40404 689498 40586 689734
rect 40822 689498 41004 689734
rect 40404 654054 41004 689498
rect 40404 653818 40586 654054
rect 40822 653818 41004 654054
rect 40404 653734 41004 653818
rect 40404 653498 40586 653734
rect 40822 653498 41004 653734
rect 40404 618054 41004 653498
rect 40404 617818 40586 618054
rect 40822 617818 41004 618054
rect 40404 617734 41004 617818
rect 40404 617498 40586 617734
rect 40822 617498 41004 617734
rect 40404 582054 41004 617498
rect 40404 581818 40586 582054
rect 40822 581818 41004 582054
rect 40404 581734 41004 581818
rect 40404 581498 40586 581734
rect 40822 581498 41004 581734
rect 40404 546054 41004 581498
rect 40404 545818 40586 546054
rect 40822 545818 41004 546054
rect 40404 545734 41004 545818
rect 40404 545498 40586 545734
rect 40822 545498 41004 545734
rect 40404 510054 41004 545498
rect 40404 509818 40586 510054
rect 40822 509818 41004 510054
rect 40404 509734 41004 509818
rect 40404 509498 40586 509734
rect 40822 509498 41004 509734
rect 40404 474054 41004 509498
rect 40404 473818 40586 474054
rect 40822 473818 41004 474054
rect 40404 473734 41004 473818
rect 40404 473498 40586 473734
rect 40822 473498 41004 473734
rect 40404 438054 41004 473498
rect 40404 437818 40586 438054
rect 40822 437818 41004 438054
rect 40404 437734 41004 437818
rect 40404 437498 40586 437734
rect 40822 437498 41004 437734
rect 40404 402054 41004 437498
rect 40404 401818 40586 402054
rect 40822 401818 41004 402054
rect 40404 401734 41004 401818
rect 40404 401498 40586 401734
rect 40822 401498 41004 401734
rect 40404 366054 41004 401498
rect 40404 365818 40586 366054
rect 40822 365818 41004 366054
rect 40404 365734 41004 365818
rect 40404 365498 40586 365734
rect 40822 365498 41004 365734
rect 40404 330054 41004 365498
rect 40404 329818 40586 330054
rect 40822 329818 41004 330054
rect 40404 329734 41004 329818
rect 40404 329498 40586 329734
rect 40822 329498 41004 329734
rect 40404 294054 41004 329498
rect 40404 293818 40586 294054
rect 40822 293818 41004 294054
rect 40404 293734 41004 293818
rect 40404 293498 40586 293734
rect 40822 293498 41004 293734
rect 40404 258054 41004 293498
rect 40404 257818 40586 258054
rect 40822 257818 41004 258054
rect 40404 257734 41004 257818
rect 40404 257498 40586 257734
rect 40822 257498 41004 257734
rect 40404 222054 41004 257498
rect 40404 221818 40586 222054
rect 40822 221818 41004 222054
rect 40404 221734 41004 221818
rect 40404 221498 40586 221734
rect 40822 221498 41004 221734
rect 40404 186054 41004 221498
rect 40404 185818 40586 186054
rect 40822 185818 41004 186054
rect 40404 185734 41004 185818
rect 40404 185498 40586 185734
rect 40822 185498 41004 185734
rect 40404 150054 41004 185498
rect 40404 149818 40586 150054
rect 40822 149818 41004 150054
rect 40404 149734 41004 149818
rect 40404 149498 40586 149734
rect 40822 149498 41004 149734
rect 40404 114054 41004 149498
rect 40404 113818 40586 114054
rect 40822 113818 41004 114054
rect 40404 113734 41004 113818
rect 40404 113498 40586 113734
rect 40822 113498 41004 113734
rect 40404 78054 41004 113498
rect 40404 77818 40586 78054
rect 40822 77818 41004 78054
rect 40404 77734 41004 77818
rect 40404 77498 40586 77734
rect 40822 77498 41004 77734
rect 40404 42054 41004 77498
rect 40404 41818 40586 42054
rect 40822 41818 41004 42054
rect 40404 41734 41004 41818
rect 40404 41498 40586 41734
rect 40822 41498 41004 41734
rect 40404 6054 41004 41498
rect 40404 5818 40586 6054
rect 40822 5818 41004 6054
rect 40404 5734 41004 5818
rect 40404 5498 40586 5734
rect 40822 5498 41004 5734
rect 40404 -2226 41004 5498
rect 40404 -2462 40586 -2226
rect 40822 -2462 41004 -2226
rect 40404 -2546 41004 -2462
rect 40404 -2782 40586 -2546
rect 40822 -2782 41004 -2546
rect 40404 -3744 41004 -2782
rect 44004 693654 44604 708042
rect 44004 693418 44186 693654
rect 44422 693418 44604 693654
rect 44004 693334 44604 693418
rect 44004 693098 44186 693334
rect 44422 693098 44604 693334
rect 44004 657654 44604 693098
rect 44004 657418 44186 657654
rect 44422 657418 44604 657654
rect 44004 657334 44604 657418
rect 44004 657098 44186 657334
rect 44422 657098 44604 657334
rect 44004 621654 44604 657098
rect 44004 621418 44186 621654
rect 44422 621418 44604 621654
rect 44004 621334 44604 621418
rect 44004 621098 44186 621334
rect 44422 621098 44604 621334
rect 44004 585654 44604 621098
rect 44004 585418 44186 585654
rect 44422 585418 44604 585654
rect 44004 585334 44604 585418
rect 44004 585098 44186 585334
rect 44422 585098 44604 585334
rect 44004 549654 44604 585098
rect 44004 549418 44186 549654
rect 44422 549418 44604 549654
rect 44004 549334 44604 549418
rect 44004 549098 44186 549334
rect 44422 549098 44604 549334
rect 44004 513654 44604 549098
rect 44004 513418 44186 513654
rect 44422 513418 44604 513654
rect 44004 513334 44604 513418
rect 44004 513098 44186 513334
rect 44422 513098 44604 513334
rect 44004 477654 44604 513098
rect 44004 477418 44186 477654
rect 44422 477418 44604 477654
rect 44004 477334 44604 477418
rect 44004 477098 44186 477334
rect 44422 477098 44604 477334
rect 44004 441654 44604 477098
rect 44004 441418 44186 441654
rect 44422 441418 44604 441654
rect 44004 441334 44604 441418
rect 44004 441098 44186 441334
rect 44422 441098 44604 441334
rect 44004 405654 44604 441098
rect 44004 405418 44186 405654
rect 44422 405418 44604 405654
rect 44004 405334 44604 405418
rect 44004 405098 44186 405334
rect 44422 405098 44604 405334
rect 44004 369654 44604 405098
rect 44004 369418 44186 369654
rect 44422 369418 44604 369654
rect 44004 369334 44604 369418
rect 44004 369098 44186 369334
rect 44422 369098 44604 369334
rect 44004 333654 44604 369098
rect 44004 333418 44186 333654
rect 44422 333418 44604 333654
rect 44004 333334 44604 333418
rect 44004 333098 44186 333334
rect 44422 333098 44604 333334
rect 44004 297654 44604 333098
rect 44004 297418 44186 297654
rect 44422 297418 44604 297654
rect 44004 297334 44604 297418
rect 44004 297098 44186 297334
rect 44422 297098 44604 297334
rect 44004 261654 44604 297098
rect 44004 261418 44186 261654
rect 44422 261418 44604 261654
rect 44004 261334 44604 261418
rect 44004 261098 44186 261334
rect 44422 261098 44604 261334
rect 44004 225654 44604 261098
rect 44004 225418 44186 225654
rect 44422 225418 44604 225654
rect 44004 225334 44604 225418
rect 44004 225098 44186 225334
rect 44422 225098 44604 225334
rect 44004 189654 44604 225098
rect 44004 189418 44186 189654
rect 44422 189418 44604 189654
rect 44004 189334 44604 189418
rect 44004 189098 44186 189334
rect 44422 189098 44604 189334
rect 44004 153654 44604 189098
rect 44004 153418 44186 153654
rect 44422 153418 44604 153654
rect 44004 153334 44604 153418
rect 44004 153098 44186 153334
rect 44422 153098 44604 153334
rect 44004 117654 44604 153098
rect 44004 117418 44186 117654
rect 44422 117418 44604 117654
rect 44004 117334 44604 117418
rect 44004 117098 44186 117334
rect 44422 117098 44604 117334
rect 44004 81654 44604 117098
rect 44004 81418 44186 81654
rect 44422 81418 44604 81654
rect 44004 81334 44604 81418
rect 44004 81098 44186 81334
rect 44422 81098 44604 81334
rect 44004 45654 44604 81098
rect 44004 45418 44186 45654
rect 44422 45418 44604 45654
rect 44004 45334 44604 45418
rect 44004 45098 44186 45334
rect 44422 45098 44604 45334
rect 44004 9654 44604 45098
rect 44004 9418 44186 9654
rect 44422 9418 44604 9654
rect 44004 9334 44604 9418
rect 44004 9098 44186 9334
rect 44422 9098 44604 9334
rect 44004 -4106 44604 9098
rect 44004 -4342 44186 -4106
rect 44422 -4342 44604 -4106
rect 44004 -4426 44604 -4342
rect 44004 -4662 44186 -4426
rect 44422 -4662 44604 -4426
rect 44004 -5624 44604 -4662
rect 47604 697254 48204 709922
rect 65604 711418 66204 711440
rect 65604 711182 65786 711418
rect 66022 711182 66204 711418
rect 65604 711098 66204 711182
rect 65604 710862 65786 711098
rect 66022 710862 66204 711098
rect 62004 709538 62604 709560
rect 62004 709302 62186 709538
rect 62422 709302 62604 709538
rect 62004 709218 62604 709302
rect 62004 708982 62186 709218
rect 62422 708982 62604 709218
rect 58404 707658 59004 707680
rect 58404 707422 58586 707658
rect 58822 707422 59004 707658
rect 58404 707338 59004 707422
rect 58404 707102 58586 707338
rect 58822 707102 59004 707338
rect 47604 697018 47786 697254
rect 48022 697018 48204 697254
rect 47604 696934 48204 697018
rect 47604 696698 47786 696934
rect 48022 696698 48204 696934
rect 47604 661254 48204 696698
rect 47604 661018 47786 661254
rect 48022 661018 48204 661254
rect 47604 660934 48204 661018
rect 47604 660698 47786 660934
rect 48022 660698 48204 660934
rect 47604 625254 48204 660698
rect 47604 625018 47786 625254
rect 48022 625018 48204 625254
rect 47604 624934 48204 625018
rect 47604 624698 47786 624934
rect 48022 624698 48204 624934
rect 47604 589254 48204 624698
rect 47604 589018 47786 589254
rect 48022 589018 48204 589254
rect 47604 588934 48204 589018
rect 47604 588698 47786 588934
rect 48022 588698 48204 588934
rect 47604 553254 48204 588698
rect 47604 553018 47786 553254
rect 48022 553018 48204 553254
rect 47604 552934 48204 553018
rect 47604 552698 47786 552934
rect 48022 552698 48204 552934
rect 47604 517254 48204 552698
rect 47604 517018 47786 517254
rect 48022 517018 48204 517254
rect 47604 516934 48204 517018
rect 47604 516698 47786 516934
rect 48022 516698 48204 516934
rect 47604 481254 48204 516698
rect 47604 481018 47786 481254
rect 48022 481018 48204 481254
rect 47604 480934 48204 481018
rect 47604 480698 47786 480934
rect 48022 480698 48204 480934
rect 47604 445254 48204 480698
rect 47604 445018 47786 445254
rect 48022 445018 48204 445254
rect 47604 444934 48204 445018
rect 47604 444698 47786 444934
rect 48022 444698 48204 444934
rect 47604 409254 48204 444698
rect 47604 409018 47786 409254
rect 48022 409018 48204 409254
rect 47604 408934 48204 409018
rect 47604 408698 47786 408934
rect 48022 408698 48204 408934
rect 47604 373254 48204 408698
rect 47604 373018 47786 373254
rect 48022 373018 48204 373254
rect 47604 372934 48204 373018
rect 47604 372698 47786 372934
rect 48022 372698 48204 372934
rect 47604 337254 48204 372698
rect 47604 337018 47786 337254
rect 48022 337018 48204 337254
rect 47604 336934 48204 337018
rect 47604 336698 47786 336934
rect 48022 336698 48204 336934
rect 47604 301254 48204 336698
rect 47604 301018 47786 301254
rect 48022 301018 48204 301254
rect 47604 300934 48204 301018
rect 47604 300698 47786 300934
rect 48022 300698 48204 300934
rect 47604 265254 48204 300698
rect 47604 265018 47786 265254
rect 48022 265018 48204 265254
rect 47604 264934 48204 265018
rect 47604 264698 47786 264934
rect 48022 264698 48204 264934
rect 47604 229254 48204 264698
rect 47604 229018 47786 229254
rect 48022 229018 48204 229254
rect 47604 228934 48204 229018
rect 47604 228698 47786 228934
rect 48022 228698 48204 228934
rect 47604 193254 48204 228698
rect 47604 193018 47786 193254
rect 48022 193018 48204 193254
rect 47604 192934 48204 193018
rect 47604 192698 47786 192934
rect 48022 192698 48204 192934
rect 47604 157254 48204 192698
rect 47604 157018 47786 157254
rect 48022 157018 48204 157254
rect 47604 156934 48204 157018
rect 47604 156698 47786 156934
rect 48022 156698 48204 156934
rect 47604 121254 48204 156698
rect 47604 121018 47786 121254
rect 48022 121018 48204 121254
rect 47604 120934 48204 121018
rect 47604 120698 47786 120934
rect 48022 120698 48204 120934
rect 47604 85254 48204 120698
rect 47604 85018 47786 85254
rect 48022 85018 48204 85254
rect 47604 84934 48204 85018
rect 47604 84698 47786 84934
rect 48022 84698 48204 84934
rect 47604 49254 48204 84698
rect 47604 49018 47786 49254
rect 48022 49018 48204 49254
rect 47604 48934 48204 49018
rect 47604 48698 47786 48934
rect 48022 48698 48204 48934
rect 47604 13254 48204 48698
rect 47604 13018 47786 13254
rect 48022 13018 48204 13254
rect 47604 12934 48204 13018
rect 47604 12698 47786 12934
rect 48022 12698 48204 12934
rect 29604 -7162 29786 -6926
rect 30022 -7162 30204 -6926
rect 29604 -7246 30204 -7162
rect 29604 -7482 29786 -7246
rect 30022 -7482 30204 -7246
rect 29604 -7504 30204 -7482
rect 47604 -5986 48204 12698
rect 54804 705778 55404 705800
rect 54804 705542 54986 705778
rect 55222 705542 55404 705778
rect 54804 705458 55404 705542
rect 54804 705222 54986 705458
rect 55222 705222 55404 705458
rect 54804 668454 55404 705222
rect 54804 668218 54986 668454
rect 55222 668218 55404 668454
rect 54804 668134 55404 668218
rect 54804 667898 54986 668134
rect 55222 667898 55404 668134
rect 54804 632454 55404 667898
rect 54804 632218 54986 632454
rect 55222 632218 55404 632454
rect 54804 632134 55404 632218
rect 54804 631898 54986 632134
rect 55222 631898 55404 632134
rect 54804 596454 55404 631898
rect 54804 596218 54986 596454
rect 55222 596218 55404 596454
rect 54804 596134 55404 596218
rect 54804 595898 54986 596134
rect 55222 595898 55404 596134
rect 54804 560454 55404 595898
rect 54804 560218 54986 560454
rect 55222 560218 55404 560454
rect 54804 560134 55404 560218
rect 54804 559898 54986 560134
rect 55222 559898 55404 560134
rect 54804 524454 55404 559898
rect 54804 524218 54986 524454
rect 55222 524218 55404 524454
rect 54804 524134 55404 524218
rect 54804 523898 54986 524134
rect 55222 523898 55404 524134
rect 54804 488454 55404 523898
rect 54804 488218 54986 488454
rect 55222 488218 55404 488454
rect 54804 488134 55404 488218
rect 54804 487898 54986 488134
rect 55222 487898 55404 488134
rect 54804 452454 55404 487898
rect 54804 452218 54986 452454
rect 55222 452218 55404 452454
rect 54804 452134 55404 452218
rect 54804 451898 54986 452134
rect 55222 451898 55404 452134
rect 54804 416454 55404 451898
rect 54804 416218 54986 416454
rect 55222 416218 55404 416454
rect 54804 416134 55404 416218
rect 54804 415898 54986 416134
rect 55222 415898 55404 416134
rect 54804 380454 55404 415898
rect 54804 380218 54986 380454
rect 55222 380218 55404 380454
rect 54804 380134 55404 380218
rect 54804 379898 54986 380134
rect 55222 379898 55404 380134
rect 54804 344454 55404 379898
rect 54804 344218 54986 344454
rect 55222 344218 55404 344454
rect 54804 344134 55404 344218
rect 54804 343898 54986 344134
rect 55222 343898 55404 344134
rect 54804 308454 55404 343898
rect 54804 308218 54986 308454
rect 55222 308218 55404 308454
rect 54804 308134 55404 308218
rect 54804 307898 54986 308134
rect 55222 307898 55404 308134
rect 54804 272454 55404 307898
rect 54804 272218 54986 272454
rect 55222 272218 55404 272454
rect 54804 272134 55404 272218
rect 54804 271898 54986 272134
rect 55222 271898 55404 272134
rect 54804 236454 55404 271898
rect 54804 236218 54986 236454
rect 55222 236218 55404 236454
rect 54804 236134 55404 236218
rect 54804 235898 54986 236134
rect 55222 235898 55404 236134
rect 54804 200454 55404 235898
rect 54804 200218 54986 200454
rect 55222 200218 55404 200454
rect 54804 200134 55404 200218
rect 54804 199898 54986 200134
rect 55222 199898 55404 200134
rect 54804 164454 55404 199898
rect 54804 164218 54986 164454
rect 55222 164218 55404 164454
rect 54804 164134 55404 164218
rect 54804 163898 54986 164134
rect 55222 163898 55404 164134
rect 54804 128454 55404 163898
rect 54804 128218 54986 128454
rect 55222 128218 55404 128454
rect 54804 128134 55404 128218
rect 54804 127898 54986 128134
rect 55222 127898 55404 128134
rect 54804 92454 55404 127898
rect 54804 92218 54986 92454
rect 55222 92218 55404 92454
rect 54804 92134 55404 92218
rect 54804 91898 54986 92134
rect 55222 91898 55404 92134
rect 54804 56454 55404 91898
rect 54804 56218 54986 56454
rect 55222 56218 55404 56454
rect 54804 56134 55404 56218
rect 54804 55898 54986 56134
rect 55222 55898 55404 56134
rect 54804 20454 55404 55898
rect 54804 20218 54986 20454
rect 55222 20218 55404 20454
rect 54804 20134 55404 20218
rect 54804 19898 54986 20134
rect 55222 19898 55404 20134
rect 54804 -1286 55404 19898
rect 54804 -1522 54986 -1286
rect 55222 -1522 55404 -1286
rect 54804 -1606 55404 -1522
rect 54804 -1842 54986 -1606
rect 55222 -1842 55404 -1606
rect 54804 -1864 55404 -1842
rect 58404 672054 59004 707102
rect 58404 671818 58586 672054
rect 58822 671818 59004 672054
rect 58404 671734 59004 671818
rect 58404 671498 58586 671734
rect 58822 671498 59004 671734
rect 58404 636054 59004 671498
rect 58404 635818 58586 636054
rect 58822 635818 59004 636054
rect 58404 635734 59004 635818
rect 58404 635498 58586 635734
rect 58822 635498 59004 635734
rect 58404 600054 59004 635498
rect 58404 599818 58586 600054
rect 58822 599818 59004 600054
rect 58404 599734 59004 599818
rect 58404 599498 58586 599734
rect 58822 599498 59004 599734
rect 58404 564054 59004 599498
rect 58404 563818 58586 564054
rect 58822 563818 59004 564054
rect 58404 563734 59004 563818
rect 58404 563498 58586 563734
rect 58822 563498 59004 563734
rect 58404 528054 59004 563498
rect 58404 527818 58586 528054
rect 58822 527818 59004 528054
rect 58404 527734 59004 527818
rect 58404 527498 58586 527734
rect 58822 527498 59004 527734
rect 58404 492054 59004 527498
rect 58404 491818 58586 492054
rect 58822 491818 59004 492054
rect 58404 491734 59004 491818
rect 58404 491498 58586 491734
rect 58822 491498 59004 491734
rect 58404 456054 59004 491498
rect 58404 455818 58586 456054
rect 58822 455818 59004 456054
rect 58404 455734 59004 455818
rect 58404 455498 58586 455734
rect 58822 455498 59004 455734
rect 58404 420054 59004 455498
rect 58404 419818 58586 420054
rect 58822 419818 59004 420054
rect 58404 419734 59004 419818
rect 58404 419498 58586 419734
rect 58822 419498 59004 419734
rect 58404 384054 59004 419498
rect 58404 383818 58586 384054
rect 58822 383818 59004 384054
rect 58404 383734 59004 383818
rect 58404 383498 58586 383734
rect 58822 383498 59004 383734
rect 58404 348054 59004 383498
rect 58404 347818 58586 348054
rect 58822 347818 59004 348054
rect 58404 347734 59004 347818
rect 58404 347498 58586 347734
rect 58822 347498 59004 347734
rect 58404 312054 59004 347498
rect 58404 311818 58586 312054
rect 58822 311818 59004 312054
rect 58404 311734 59004 311818
rect 58404 311498 58586 311734
rect 58822 311498 59004 311734
rect 58404 276054 59004 311498
rect 58404 275818 58586 276054
rect 58822 275818 59004 276054
rect 58404 275734 59004 275818
rect 58404 275498 58586 275734
rect 58822 275498 59004 275734
rect 58404 240054 59004 275498
rect 58404 239818 58586 240054
rect 58822 239818 59004 240054
rect 58404 239734 59004 239818
rect 58404 239498 58586 239734
rect 58822 239498 59004 239734
rect 58404 204054 59004 239498
rect 58404 203818 58586 204054
rect 58822 203818 59004 204054
rect 58404 203734 59004 203818
rect 58404 203498 58586 203734
rect 58822 203498 59004 203734
rect 58404 168054 59004 203498
rect 58404 167818 58586 168054
rect 58822 167818 59004 168054
rect 58404 167734 59004 167818
rect 58404 167498 58586 167734
rect 58822 167498 59004 167734
rect 58404 132054 59004 167498
rect 58404 131818 58586 132054
rect 58822 131818 59004 132054
rect 58404 131734 59004 131818
rect 58404 131498 58586 131734
rect 58822 131498 59004 131734
rect 58404 96054 59004 131498
rect 58404 95818 58586 96054
rect 58822 95818 59004 96054
rect 58404 95734 59004 95818
rect 58404 95498 58586 95734
rect 58822 95498 59004 95734
rect 58404 60054 59004 95498
rect 58404 59818 58586 60054
rect 58822 59818 59004 60054
rect 58404 59734 59004 59818
rect 58404 59498 58586 59734
rect 58822 59498 59004 59734
rect 58404 24054 59004 59498
rect 58404 23818 58586 24054
rect 58822 23818 59004 24054
rect 58404 23734 59004 23818
rect 58404 23498 58586 23734
rect 58822 23498 59004 23734
rect 58404 -3166 59004 23498
rect 58404 -3402 58586 -3166
rect 58822 -3402 59004 -3166
rect 58404 -3486 59004 -3402
rect 58404 -3722 58586 -3486
rect 58822 -3722 59004 -3486
rect 58404 -3744 59004 -3722
rect 62004 675654 62604 708982
rect 62004 675418 62186 675654
rect 62422 675418 62604 675654
rect 62004 675334 62604 675418
rect 62004 675098 62186 675334
rect 62422 675098 62604 675334
rect 62004 639654 62604 675098
rect 62004 639418 62186 639654
rect 62422 639418 62604 639654
rect 62004 639334 62604 639418
rect 62004 639098 62186 639334
rect 62422 639098 62604 639334
rect 62004 603654 62604 639098
rect 62004 603418 62186 603654
rect 62422 603418 62604 603654
rect 62004 603334 62604 603418
rect 62004 603098 62186 603334
rect 62422 603098 62604 603334
rect 62004 567654 62604 603098
rect 62004 567418 62186 567654
rect 62422 567418 62604 567654
rect 62004 567334 62604 567418
rect 62004 567098 62186 567334
rect 62422 567098 62604 567334
rect 62004 531654 62604 567098
rect 62004 531418 62186 531654
rect 62422 531418 62604 531654
rect 62004 531334 62604 531418
rect 62004 531098 62186 531334
rect 62422 531098 62604 531334
rect 62004 495654 62604 531098
rect 62004 495418 62186 495654
rect 62422 495418 62604 495654
rect 62004 495334 62604 495418
rect 62004 495098 62186 495334
rect 62422 495098 62604 495334
rect 62004 459654 62604 495098
rect 62004 459418 62186 459654
rect 62422 459418 62604 459654
rect 62004 459334 62604 459418
rect 62004 459098 62186 459334
rect 62422 459098 62604 459334
rect 62004 423654 62604 459098
rect 62004 423418 62186 423654
rect 62422 423418 62604 423654
rect 62004 423334 62604 423418
rect 62004 423098 62186 423334
rect 62422 423098 62604 423334
rect 62004 387654 62604 423098
rect 62004 387418 62186 387654
rect 62422 387418 62604 387654
rect 62004 387334 62604 387418
rect 62004 387098 62186 387334
rect 62422 387098 62604 387334
rect 62004 351654 62604 387098
rect 62004 351418 62186 351654
rect 62422 351418 62604 351654
rect 62004 351334 62604 351418
rect 62004 351098 62186 351334
rect 62422 351098 62604 351334
rect 62004 315654 62604 351098
rect 62004 315418 62186 315654
rect 62422 315418 62604 315654
rect 62004 315334 62604 315418
rect 62004 315098 62186 315334
rect 62422 315098 62604 315334
rect 62004 279654 62604 315098
rect 62004 279418 62186 279654
rect 62422 279418 62604 279654
rect 62004 279334 62604 279418
rect 62004 279098 62186 279334
rect 62422 279098 62604 279334
rect 62004 243654 62604 279098
rect 62004 243418 62186 243654
rect 62422 243418 62604 243654
rect 62004 243334 62604 243418
rect 62004 243098 62186 243334
rect 62422 243098 62604 243334
rect 62004 207654 62604 243098
rect 62004 207418 62186 207654
rect 62422 207418 62604 207654
rect 62004 207334 62604 207418
rect 62004 207098 62186 207334
rect 62422 207098 62604 207334
rect 62004 171654 62604 207098
rect 62004 171418 62186 171654
rect 62422 171418 62604 171654
rect 62004 171334 62604 171418
rect 62004 171098 62186 171334
rect 62422 171098 62604 171334
rect 62004 135654 62604 171098
rect 62004 135418 62186 135654
rect 62422 135418 62604 135654
rect 62004 135334 62604 135418
rect 62004 135098 62186 135334
rect 62422 135098 62604 135334
rect 62004 99654 62604 135098
rect 62004 99418 62186 99654
rect 62422 99418 62604 99654
rect 62004 99334 62604 99418
rect 62004 99098 62186 99334
rect 62422 99098 62604 99334
rect 62004 63654 62604 99098
rect 62004 63418 62186 63654
rect 62422 63418 62604 63654
rect 62004 63334 62604 63418
rect 62004 63098 62186 63334
rect 62422 63098 62604 63334
rect 62004 27654 62604 63098
rect 62004 27418 62186 27654
rect 62422 27418 62604 27654
rect 62004 27334 62604 27418
rect 62004 27098 62186 27334
rect 62422 27098 62604 27334
rect 62004 -5046 62604 27098
rect 62004 -5282 62186 -5046
rect 62422 -5282 62604 -5046
rect 62004 -5366 62604 -5282
rect 62004 -5602 62186 -5366
rect 62422 -5602 62604 -5366
rect 62004 -5624 62604 -5602
rect 65604 679254 66204 710862
rect 83604 710478 84204 711440
rect 83604 710242 83786 710478
rect 84022 710242 84204 710478
rect 83604 710158 84204 710242
rect 83604 709922 83786 710158
rect 84022 709922 84204 710158
rect 80004 708598 80604 709560
rect 80004 708362 80186 708598
rect 80422 708362 80604 708598
rect 80004 708278 80604 708362
rect 80004 708042 80186 708278
rect 80422 708042 80604 708278
rect 76404 706718 77004 707680
rect 76404 706482 76586 706718
rect 76822 706482 77004 706718
rect 76404 706398 77004 706482
rect 76404 706162 76586 706398
rect 76822 706162 77004 706398
rect 65604 679018 65786 679254
rect 66022 679018 66204 679254
rect 65604 678934 66204 679018
rect 65604 678698 65786 678934
rect 66022 678698 66204 678934
rect 65604 643254 66204 678698
rect 65604 643018 65786 643254
rect 66022 643018 66204 643254
rect 65604 642934 66204 643018
rect 65604 642698 65786 642934
rect 66022 642698 66204 642934
rect 65604 607254 66204 642698
rect 65604 607018 65786 607254
rect 66022 607018 66204 607254
rect 65604 606934 66204 607018
rect 65604 606698 65786 606934
rect 66022 606698 66204 606934
rect 65604 571254 66204 606698
rect 65604 571018 65786 571254
rect 66022 571018 66204 571254
rect 65604 570934 66204 571018
rect 65604 570698 65786 570934
rect 66022 570698 66204 570934
rect 65604 535254 66204 570698
rect 65604 535018 65786 535254
rect 66022 535018 66204 535254
rect 65604 534934 66204 535018
rect 65604 534698 65786 534934
rect 66022 534698 66204 534934
rect 65604 499254 66204 534698
rect 65604 499018 65786 499254
rect 66022 499018 66204 499254
rect 65604 498934 66204 499018
rect 65604 498698 65786 498934
rect 66022 498698 66204 498934
rect 65604 463254 66204 498698
rect 65604 463018 65786 463254
rect 66022 463018 66204 463254
rect 65604 462934 66204 463018
rect 65604 462698 65786 462934
rect 66022 462698 66204 462934
rect 65604 427254 66204 462698
rect 65604 427018 65786 427254
rect 66022 427018 66204 427254
rect 65604 426934 66204 427018
rect 65604 426698 65786 426934
rect 66022 426698 66204 426934
rect 65604 391254 66204 426698
rect 65604 391018 65786 391254
rect 66022 391018 66204 391254
rect 65604 390934 66204 391018
rect 65604 390698 65786 390934
rect 66022 390698 66204 390934
rect 65604 355254 66204 390698
rect 65604 355018 65786 355254
rect 66022 355018 66204 355254
rect 65604 354934 66204 355018
rect 65604 354698 65786 354934
rect 66022 354698 66204 354934
rect 65604 319254 66204 354698
rect 65604 319018 65786 319254
rect 66022 319018 66204 319254
rect 65604 318934 66204 319018
rect 65604 318698 65786 318934
rect 66022 318698 66204 318934
rect 65604 283254 66204 318698
rect 65604 283018 65786 283254
rect 66022 283018 66204 283254
rect 65604 282934 66204 283018
rect 65604 282698 65786 282934
rect 66022 282698 66204 282934
rect 65604 247254 66204 282698
rect 65604 247018 65786 247254
rect 66022 247018 66204 247254
rect 65604 246934 66204 247018
rect 65604 246698 65786 246934
rect 66022 246698 66204 246934
rect 65604 211254 66204 246698
rect 65604 211018 65786 211254
rect 66022 211018 66204 211254
rect 65604 210934 66204 211018
rect 65604 210698 65786 210934
rect 66022 210698 66204 210934
rect 65604 175254 66204 210698
rect 65604 175018 65786 175254
rect 66022 175018 66204 175254
rect 65604 174934 66204 175018
rect 65604 174698 65786 174934
rect 66022 174698 66204 174934
rect 65604 139254 66204 174698
rect 65604 139018 65786 139254
rect 66022 139018 66204 139254
rect 65604 138934 66204 139018
rect 65604 138698 65786 138934
rect 66022 138698 66204 138934
rect 65604 103254 66204 138698
rect 65604 103018 65786 103254
rect 66022 103018 66204 103254
rect 65604 102934 66204 103018
rect 65604 102698 65786 102934
rect 66022 102698 66204 102934
rect 65604 67254 66204 102698
rect 65604 67018 65786 67254
rect 66022 67018 66204 67254
rect 65604 66934 66204 67018
rect 65604 66698 65786 66934
rect 66022 66698 66204 66934
rect 65604 31254 66204 66698
rect 65604 31018 65786 31254
rect 66022 31018 66204 31254
rect 65604 30934 66204 31018
rect 65604 30698 65786 30934
rect 66022 30698 66204 30934
rect 47604 -6222 47786 -5986
rect 48022 -6222 48204 -5986
rect 47604 -6306 48204 -6222
rect 47604 -6542 47786 -6306
rect 48022 -6542 48204 -6306
rect 47604 -7504 48204 -6542
rect 65604 -6926 66204 30698
rect 72804 704838 73404 705800
rect 72804 704602 72986 704838
rect 73222 704602 73404 704838
rect 72804 704518 73404 704602
rect 72804 704282 72986 704518
rect 73222 704282 73404 704518
rect 72804 686454 73404 704282
rect 72804 686218 72986 686454
rect 73222 686218 73404 686454
rect 72804 686134 73404 686218
rect 72804 685898 72986 686134
rect 73222 685898 73404 686134
rect 72804 650454 73404 685898
rect 72804 650218 72986 650454
rect 73222 650218 73404 650454
rect 72804 650134 73404 650218
rect 72804 649898 72986 650134
rect 73222 649898 73404 650134
rect 72804 614454 73404 649898
rect 72804 614218 72986 614454
rect 73222 614218 73404 614454
rect 72804 614134 73404 614218
rect 72804 613898 72986 614134
rect 73222 613898 73404 614134
rect 72804 578454 73404 613898
rect 72804 578218 72986 578454
rect 73222 578218 73404 578454
rect 72804 578134 73404 578218
rect 72804 577898 72986 578134
rect 73222 577898 73404 578134
rect 72804 542454 73404 577898
rect 72804 542218 72986 542454
rect 73222 542218 73404 542454
rect 72804 542134 73404 542218
rect 72804 541898 72986 542134
rect 73222 541898 73404 542134
rect 72804 506454 73404 541898
rect 72804 506218 72986 506454
rect 73222 506218 73404 506454
rect 72804 506134 73404 506218
rect 72804 505898 72986 506134
rect 73222 505898 73404 506134
rect 72804 470454 73404 505898
rect 72804 470218 72986 470454
rect 73222 470218 73404 470454
rect 72804 470134 73404 470218
rect 72804 469898 72986 470134
rect 73222 469898 73404 470134
rect 72804 434454 73404 469898
rect 72804 434218 72986 434454
rect 73222 434218 73404 434454
rect 72804 434134 73404 434218
rect 72804 433898 72986 434134
rect 73222 433898 73404 434134
rect 72804 398454 73404 433898
rect 72804 398218 72986 398454
rect 73222 398218 73404 398454
rect 72804 398134 73404 398218
rect 72804 397898 72986 398134
rect 73222 397898 73404 398134
rect 72804 362454 73404 397898
rect 72804 362218 72986 362454
rect 73222 362218 73404 362454
rect 72804 362134 73404 362218
rect 72804 361898 72986 362134
rect 73222 361898 73404 362134
rect 72804 326454 73404 361898
rect 72804 326218 72986 326454
rect 73222 326218 73404 326454
rect 72804 326134 73404 326218
rect 72804 325898 72986 326134
rect 73222 325898 73404 326134
rect 72804 290454 73404 325898
rect 72804 290218 72986 290454
rect 73222 290218 73404 290454
rect 72804 290134 73404 290218
rect 72804 289898 72986 290134
rect 73222 289898 73404 290134
rect 72804 254454 73404 289898
rect 72804 254218 72986 254454
rect 73222 254218 73404 254454
rect 72804 254134 73404 254218
rect 72804 253898 72986 254134
rect 73222 253898 73404 254134
rect 72804 218454 73404 253898
rect 72804 218218 72986 218454
rect 73222 218218 73404 218454
rect 72804 218134 73404 218218
rect 72804 217898 72986 218134
rect 73222 217898 73404 218134
rect 72804 182454 73404 217898
rect 72804 182218 72986 182454
rect 73222 182218 73404 182454
rect 72804 182134 73404 182218
rect 72804 181898 72986 182134
rect 73222 181898 73404 182134
rect 72804 146454 73404 181898
rect 72804 146218 72986 146454
rect 73222 146218 73404 146454
rect 72804 146134 73404 146218
rect 72804 145898 72986 146134
rect 73222 145898 73404 146134
rect 72804 110454 73404 145898
rect 72804 110218 72986 110454
rect 73222 110218 73404 110454
rect 72804 110134 73404 110218
rect 72804 109898 72986 110134
rect 73222 109898 73404 110134
rect 72804 74454 73404 109898
rect 72804 74218 72986 74454
rect 73222 74218 73404 74454
rect 72804 74134 73404 74218
rect 72804 73898 72986 74134
rect 73222 73898 73404 74134
rect 72804 38454 73404 73898
rect 72804 38218 72986 38454
rect 73222 38218 73404 38454
rect 72804 38134 73404 38218
rect 72804 37898 72986 38134
rect 73222 37898 73404 38134
rect 72804 2454 73404 37898
rect 72804 2218 72986 2454
rect 73222 2218 73404 2454
rect 72804 2134 73404 2218
rect 72804 1898 72986 2134
rect 73222 1898 73404 2134
rect 72804 -346 73404 1898
rect 72804 -582 72986 -346
rect 73222 -582 73404 -346
rect 72804 -666 73404 -582
rect 72804 -902 72986 -666
rect 73222 -902 73404 -666
rect 72804 -1864 73404 -902
rect 76404 690054 77004 706162
rect 76404 689818 76586 690054
rect 76822 689818 77004 690054
rect 76404 689734 77004 689818
rect 76404 689498 76586 689734
rect 76822 689498 77004 689734
rect 76404 654054 77004 689498
rect 76404 653818 76586 654054
rect 76822 653818 77004 654054
rect 76404 653734 77004 653818
rect 76404 653498 76586 653734
rect 76822 653498 77004 653734
rect 76404 618054 77004 653498
rect 76404 617818 76586 618054
rect 76822 617818 77004 618054
rect 76404 617734 77004 617818
rect 76404 617498 76586 617734
rect 76822 617498 77004 617734
rect 76404 582054 77004 617498
rect 76404 581818 76586 582054
rect 76822 581818 77004 582054
rect 76404 581734 77004 581818
rect 76404 581498 76586 581734
rect 76822 581498 77004 581734
rect 76404 546054 77004 581498
rect 76404 545818 76586 546054
rect 76822 545818 77004 546054
rect 76404 545734 77004 545818
rect 76404 545498 76586 545734
rect 76822 545498 77004 545734
rect 76404 510054 77004 545498
rect 76404 509818 76586 510054
rect 76822 509818 77004 510054
rect 76404 509734 77004 509818
rect 76404 509498 76586 509734
rect 76822 509498 77004 509734
rect 76404 474054 77004 509498
rect 76404 473818 76586 474054
rect 76822 473818 77004 474054
rect 76404 473734 77004 473818
rect 76404 473498 76586 473734
rect 76822 473498 77004 473734
rect 76404 438054 77004 473498
rect 76404 437818 76586 438054
rect 76822 437818 77004 438054
rect 76404 437734 77004 437818
rect 76404 437498 76586 437734
rect 76822 437498 77004 437734
rect 76404 402054 77004 437498
rect 76404 401818 76586 402054
rect 76822 401818 77004 402054
rect 76404 401734 77004 401818
rect 76404 401498 76586 401734
rect 76822 401498 77004 401734
rect 76404 366054 77004 401498
rect 76404 365818 76586 366054
rect 76822 365818 77004 366054
rect 76404 365734 77004 365818
rect 76404 365498 76586 365734
rect 76822 365498 77004 365734
rect 76404 330054 77004 365498
rect 76404 329818 76586 330054
rect 76822 329818 77004 330054
rect 76404 329734 77004 329818
rect 76404 329498 76586 329734
rect 76822 329498 77004 329734
rect 76404 294054 77004 329498
rect 76404 293818 76586 294054
rect 76822 293818 77004 294054
rect 76404 293734 77004 293818
rect 76404 293498 76586 293734
rect 76822 293498 77004 293734
rect 76404 258054 77004 293498
rect 76404 257818 76586 258054
rect 76822 257818 77004 258054
rect 76404 257734 77004 257818
rect 76404 257498 76586 257734
rect 76822 257498 77004 257734
rect 76404 222054 77004 257498
rect 76404 221818 76586 222054
rect 76822 221818 77004 222054
rect 76404 221734 77004 221818
rect 76404 221498 76586 221734
rect 76822 221498 77004 221734
rect 76404 186054 77004 221498
rect 76404 185818 76586 186054
rect 76822 185818 77004 186054
rect 76404 185734 77004 185818
rect 76404 185498 76586 185734
rect 76822 185498 77004 185734
rect 76404 150054 77004 185498
rect 76404 149818 76586 150054
rect 76822 149818 77004 150054
rect 76404 149734 77004 149818
rect 76404 149498 76586 149734
rect 76822 149498 77004 149734
rect 76404 114054 77004 149498
rect 76404 113818 76586 114054
rect 76822 113818 77004 114054
rect 76404 113734 77004 113818
rect 76404 113498 76586 113734
rect 76822 113498 77004 113734
rect 76404 78054 77004 113498
rect 76404 77818 76586 78054
rect 76822 77818 77004 78054
rect 76404 77734 77004 77818
rect 76404 77498 76586 77734
rect 76822 77498 77004 77734
rect 76404 42054 77004 77498
rect 76404 41818 76586 42054
rect 76822 41818 77004 42054
rect 76404 41734 77004 41818
rect 76404 41498 76586 41734
rect 76822 41498 77004 41734
rect 76404 6054 77004 41498
rect 76404 5818 76586 6054
rect 76822 5818 77004 6054
rect 76404 5734 77004 5818
rect 76404 5498 76586 5734
rect 76822 5498 77004 5734
rect 76404 -2226 77004 5498
rect 76404 -2462 76586 -2226
rect 76822 -2462 77004 -2226
rect 76404 -2546 77004 -2462
rect 76404 -2782 76586 -2546
rect 76822 -2782 77004 -2546
rect 76404 -3744 77004 -2782
rect 80004 693654 80604 708042
rect 80004 693418 80186 693654
rect 80422 693418 80604 693654
rect 80004 693334 80604 693418
rect 80004 693098 80186 693334
rect 80422 693098 80604 693334
rect 80004 657654 80604 693098
rect 80004 657418 80186 657654
rect 80422 657418 80604 657654
rect 80004 657334 80604 657418
rect 80004 657098 80186 657334
rect 80422 657098 80604 657334
rect 80004 621654 80604 657098
rect 80004 621418 80186 621654
rect 80422 621418 80604 621654
rect 80004 621334 80604 621418
rect 80004 621098 80186 621334
rect 80422 621098 80604 621334
rect 80004 585654 80604 621098
rect 80004 585418 80186 585654
rect 80422 585418 80604 585654
rect 80004 585334 80604 585418
rect 80004 585098 80186 585334
rect 80422 585098 80604 585334
rect 80004 549654 80604 585098
rect 80004 549418 80186 549654
rect 80422 549418 80604 549654
rect 80004 549334 80604 549418
rect 80004 549098 80186 549334
rect 80422 549098 80604 549334
rect 80004 513654 80604 549098
rect 80004 513418 80186 513654
rect 80422 513418 80604 513654
rect 80004 513334 80604 513418
rect 80004 513098 80186 513334
rect 80422 513098 80604 513334
rect 80004 477654 80604 513098
rect 80004 477418 80186 477654
rect 80422 477418 80604 477654
rect 80004 477334 80604 477418
rect 80004 477098 80186 477334
rect 80422 477098 80604 477334
rect 80004 441654 80604 477098
rect 80004 441418 80186 441654
rect 80422 441418 80604 441654
rect 80004 441334 80604 441418
rect 80004 441098 80186 441334
rect 80422 441098 80604 441334
rect 80004 405654 80604 441098
rect 80004 405418 80186 405654
rect 80422 405418 80604 405654
rect 80004 405334 80604 405418
rect 80004 405098 80186 405334
rect 80422 405098 80604 405334
rect 80004 369654 80604 405098
rect 80004 369418 80186 369654
rect 80422 369418 80604 369654
rect 80004 369334 80604 369418
rect 80004 369098 80186 369334
rect 80422 369098 80604 369334
rect 80004 333654 80604 369098
rect 80004 333418 80186 333654
rect 80422 333418 80604 333654
rect 80004 333334 80604 333418
rect 80004 333098 80186 333334
rect 80422 333098 80604 333334
rect 80004 297654 80604 333098
rect 80004 297418 80186 297654
rect 80422 297418 80604 297654
rect 80004 297334 80604 297418
rect 80004 297098 80186 297334
rect 80422 297098 80604 297334
rect 80004 261654 80604 297098
rect 80004 261418 80186 261654
rect 80422 261418 80604 261654
rect 80004 261334 80604 261418
rect 80004 261098 80186 261334
rect 80422 261098 80604 261334
rect 80004 225654 80604 261098
rect 80004 225418 80186 225654
rect 80422 225418 80604 225654
rect 80004 225334 80604 225418
rect 80004 225098 80186 225334
rect 80422 225098 80604 225334
rect 80004 189654 80604 225098
rect 80004 189418 80186 189654
rect 80422 189418 80604 189654
rect 80004 189334 80604 189418
rect 80004 189098 80186 189334
rect 80422 189098 80604 189334
rect 80004 153654 80604 189098
rect 80004 153418 80186 153654
rect 80422 153418 80604 153654
rect 80004 153334 80604 153418
rect 80004 153098 80186 153334
rect 80422 153098 80604 153334
rect 80004 117654 80604 153098
rect 80004 117418 80186 117654
rect 80422 117418 80604 117654
rect 80004 117334 80604 117418
rect 80004 117098 80186 117334
rect 80422 117098 80604 117334
rect 80004 81654 80604 117098
rect 80004 81418 80186 81654
rect 80422 81418 80604 81654
rect 80004 81334 80604 81418
rect 80004 81098 80186 81334
rect 80422 81098 80604 81334
rect 80004 45654 80604 81098
rect 80004 45418 80186 45654
rect 80422 45418 80604 45654
rect 80004 45334 80604 45418
rect 80004 45098 80186 45334
rect 80422 45098 80604 45334
rect 80004 9654 80604 45098
rect 80004 9418 80186 9654
rect 80422 9418 80604 9654
rect 80004 9334 80604 9418
rect 80004 9098 80186 9334
rect 80422 9098 80604 9334
rect 80004 -4106 80604 9098
rect 80004 -4342 80186 -4106
rect 80422 -4342 80604 -4106
rect 80004 -4426 80604 -4342
rect 80004 -4662 80186 -4426
rect 80422 -4662 80604 -4426
rect 80004 -5624 80604 -4662
rect 83604 697254 84204 709922
rect 101604 711418 102204 711440
rect 101604 711182 101786 711418
rect 102022 711182 102204 711418
rect 101604 711098 102204 711182
rect 101604 710862 101786 711098
rect 102022 710862 102204 711098
rect 98004 709538 98604 709560
rect 98004 709302 98186 709538
rect 98422 709302 98604 709538
rect 98004 709218 98604 709302
rect 98004 708982 98186 709218
rect 98422 708982 98604 709218
rect 94404 707658 95004 707680
rect 94404 707422 94586 707658
rect 94822 707422 95004 707658
rect 94404 707338 95004 707422
rect 94404 707102 94586 707338
rect 94822 707102 95004 707338
rect 83604 697018 83786 697254
rect 84022 697018 84204 697254
rect 83604 696934 84204 697018
rect 83604 696698 83786 696934
rect 84022 696698 84204 696934
rect 83604 661254 84204 696698
rect 83604 661018 83786 661254
rect 84022 661018 84204 661254
rect 83604 660934 84204 661018
rect 83604 660698 83786 660934
rect 84022 660698 84204 660934
rect 83604 625254 84204 660698
rect 83604 625018 83786 625254
rect 84022 625018 84204 625254
rect 83604 624934 84204 625018
rect 83604 624698 83786 624934
rect 84022 624698 84204 624934
rect 83604 589254 84204 624698
rect 83604 589018 83786 589254
rect 84022 589018 84204 589254
rect 83604 588934 84204 589018
rect 83604 588698 83786 588934
rect 84022 588698 84204 588934
rect 83604 553254 84204 588698
rect 83604 553018 83786 553254
rect 84022 553018 84204 553254
rect 83604 552934 84204 553018
rect 83604 552698 83786 552934
rect 84022 552698 84204 552934
rect 83604 517254 84204 552698
rect 83604 517018 83786 517254
rect 84022 517018 84204 517254
rect 83604 516934 84204 517018
rect 83604 516698 83786 516934
rect 84022 516698 84204 516934
rect 83604 481254 84204 516698
rect 83604 481018 83786 481254
rect 84022 481018 84204 481254
rect 83604 480934 84204 481018
rect 83604 480698 83786 480934
rect 84022 480698 84204 480934
rect 83604 445254 84204 480698
rect 83604 445018 83786 445254
rect 84022 445018 84204 445254
rect 83604 444934 84204 445018
rect 83604 444698 83786 444934
rect 84022 444698 84204 444934
rect 83604 409254 84204 444698
rect 83604 409018 83786 409254
rect 84022 409018 84204 409254
rect 83604 408934 84204 409018
rect 83604 408698 83786 408934
rect 84022 408698 84204 408934
rect 83604 373254 84204 408698
rect 83604 373018 83786 373254
rect 84022 373018 84204 373254
rect 83604 372934 84204 373018
rect 83604 372698 83786 372934
rect 84022 372698 84204 372934
rect 83604 337254 84204 372698
rect 83604 337018 83786 337254
rect 84022 337018 84204 337254
rect 83604 336934 84204 337018
rect 83604 336698 83786 336934
rect 84022 336698 84204 336934
rect 83604 301254 84204 336698
rect 83604 301018 83786 301254
rect 84022 301018 84204 301254
rect 83604 300934 84204 301018
rect 83604 300698 83786 300934
rect 84022 300698 84204 300934
rect 83604 265254 84204 300698
rect 83604 265018 83786 265254
rect 84022 265018 84204 265254
rect 83604 264934 84204 265018
rect 83604 264698 83786 264934
rect 84022 264698 84204 264934
rect 83604 229254 84204 264698
rect 83604 229018 83786 229254
rect 84022 229018 84204 229254
rect 83604 228934 84204 229018
rect 83604 228698 83786 228934
rect 84022 228698 84204 228934
rect 83604 193254 84204 228698
rect 83604 193018 83786 193254
rect 84022 193018 84204 193254
rect 83604 192934 84204 193018
rect 83604 192698 83786 192934
rect 84022 192698 84204 192934
rect 83604 157254 84204 192698
rect 83604 157018 83786 157254
rect 84022 157018 84204 157254
rect 83604 156934 84204 157018
rect 83604 156698 83786 156934
rect 84022 156698 84204 156934
rect 83604 121254 84204 156698
rect 83604 121018 83786 121254
rect 84022 121018 84204 121254
rect 83604 120934 84204 121018
rect 83604 120698 83786 120934
rect 84022 120698 84204 120934
rect 83604 85254 84204 120698
rect 83604 85018 83786 85254
rect 84022 85018 84204 85254
rect 83604 84934 84204 85018
rect 83604 84698 83786 84934
rect 84022 84698 84204 84934
rect 83604 49254 84204 84698
rect 83604 49018 83786 49254
rect 84022 49018 84204 49254
rect 83604 48934 84204 49018
rect 83604 48698 83786 48934
rect 84022 48698 84204 48934
rect 83604 13254 84204 48698
rect 83604 13018 83786 13254
rect 84022 13018 84204 13254
rect 83604 12934 84204 13018
rect 83604 12698 83786 12934
rect 84022 12698 84204 12934
rect 65604 -7162 65786 -6926
rect 66022 -7162 66204 -6926
rect 65604 -7246 66204 -7162
rect 65604 -7482 65786 -7246
rect 66022 -7482 66204 -7246
rect 65604 -7504 66204 -7482
rect 83604 -5986 84204 12698
rect 90804 705778 91404 705800
rect 90804 705542 90986 705778
rect 91222 705542 91404 705778
rect 90804 705458 91404 705542
rect 90804 705222 90986 705458
rect 91222 705222 91404 705458
rect 90804 668454 91404 705222
rect 90804 668218 90986 668454
rect 91222 668218 91404 668454
rect 90804 668134 91404 668218
rect 90804 667898 90986 668134
rect 91222 667898 91404 668134
rect 90804 632454 91404 667898
rect 90804 632218 90986 632454
rect 91222 632218 91404 632454
rect 90804 632134 91404 632218
rect 90804 631898 90986 632134
rect 91222 631898 91404 632134
rect 90804 596454 91404 631898
rect 90804 596218 90986 596454
rect 91222 596218 91404 596454
rect 90804 596134 91404 596218
rect 90804 595898 90986 596134
rect 91222 595898 91404 596134
rect 90804 560454 91404 595898
rect 90804 560218 90986 560454
rect 91222 560218 91404 560454
rect 90804 560134 91404 560218
rect 90804 559898 90986 560134
rect 91222 559898 91404 560134
rect 90804 524454 91404 559898
rect 90804 524218 90986 524454
rect 91222 524218 91404 524454
rect 90804 524134 91404 524218
rect 90804 523898 90986 524134
rect 91222 523898 91404 524134
rect 90804 488454 91404 523898
rect 90804 488218 90986 488454
rect 91222 488218 91404 488454
rect 90804 488134 91404 488218
rect 90804 487898 90986 488134
rect 91222 487898 91404 488134
rect 90804 452454 91404 487898
rect 90804 452218 90986 452454
rect 91222 452218 91404 452454
rect 90804 452134 91404 452218
rect 90804 451898 90986 452134
rect 91222 451898 91404 452134
rect 90804 416454 91404 451898
rect 90804 416218 90986 416454
rect 91222 416218 91404 416454
rect 90804 416134 91404 416218
rect 90804 415898 90986 416134
rect 91222 415898 91404 416134
rect 90804 380454 91404 415898
rect 90804 380218 90986 380454
rect 91222 380218 91404 380454
rect 90804 380134 91404 380218
rect 90804 379898 90986 380134
rect 91222 379898 91404 380134
rect 90804 344454 91404 379898
rect 90804 344218 90986 344454
rect 91222 344218 91404 344454
rect 90804 344134 91404 344218
rect 90804 343898 90986 344134
rect 91222 343898 91404 344134
rect 90804 308454 91404 343898
rect 90804 308218 90986 308454
rect 91222 308218 91404 308454
rect 90804 308134 91404 308218
rect 90804 307898 90986 308134
rect 91222 307898 91404 308134
rect 90804 272454 91404 307898
rect 90804 272218 90986 272454
rect 91222 272218 91404 272454
rect 90804 272134 91404 272218
rect 90804 271898 90986 272134
rect 91222 271898 91404 272134
rect 90804 236454 91404 271898
rect 90804 236218 90986 236454
rect 91222 236218 91404 236454
rect 90804 236134 91404 236218
rect 90804 235898 90986 236134
rect 91222 235898 91404 236134
rect 90804 200454 91404 235898
rect 90804 200218 90986 200454
rect 91222 200218 91404 200454
rect 90804 200134 91404 200218
rect 90804 199898 90986 200134
rect 91222 199898 91404 200134
rect 90804 164454 91404 199898
rect 90804 164218 90986 164454
rect 91222 164218 91404 164454
rect 90804 164134 91404 164218
rect 90804 163898 90986 164134
rect 91222 163898 91404 164134
rect 90804 128454 91404 163898
rect 90804 128218 90986 128454
rect 91222 128218 91404 128454
rect 90804 128134 91404 128218
rect 90804 127898 90986 128134
rect 91222 127898 91404 128134
rect 90804 92454 91404 127898
rect 90804 92218 90986 92454
rect 91222 92218 91404 92454
rect 90804 92134 91404 92218
rect 90804 91898 90986 92134
rect 91222 91898 91404 92134
rect 90804 56454 91404 91898
rect 90804 56218 90986 56454
rect 91222 56218 91404 56454
rect 90804 56134 91404 56218
rect 90804 55898 90986 56134
rect 91222 55898 91404 56134
rect 90804 20454 91404 55898
rect 90804 20218 90986 20454
rect 91222 20218 91404 20454
rect 90804 20134 91404 20218
rect 90804 19898 90986 20134
rect 91222 19898 91404 20134
rect 90804 -1286 91404 19898
rect 90804 -1522 90986 -1286
rect 91222 -1522 91404 -1286
rect 90804 -1606 91404 -1522
rect 90804 -1842 90986 -1606
rect 91222 -1842 91404 -1606
rect 90804 -1864 91404 -1842
rect 94404 672054 95004 707102
rect 94404 671818 94586 672054
rect 94822 671818 95004 672054
rect 94404 671734 95004 671818
rect 94404 671498 94586 671734
rect 94822 671498 95004 671734
rect 94404 636054 95004 671498
rect 94404 635818 94586 636054
rect 94822 635818 95004 636054
rect 94404 635734 95004 635818
rect 94404 635498 94586 635734
rect 94822 635498 95004 635734
rect 94404 600054 95004 635498
rect 94404 599818 94586 600054
rect 94822 599818 95004 600054
rect 94404 599734 95004 599818
rect 94404 599498 94586 599734
rect 94822 599498 95004 599734
rect 94404 564054 95004 599498
rect 94404 563818 94586 564054
rect 94822 563818 95004 564054
rect 94404 563734 95004 563818
rect 94404 563498 94586 563734
rect 94822 563498 95004 563734
rect 94404 528054 95004 563498
rect 94404 527818 94586 528054
rect 94822 527818 95004 528054
rect 94404 527734 95004 527818
rect 94404 527498 94586 527734
rect 94822 527498 95004 527734
rect 94404 492054 95004 527498
rect 94404 491818 94586 492054
rect 94822 491818 95004 492054
rect 94404 491734 95004 491818
rect 94404 491498 94586 491734
rect 94822 491498 95004 491734
rect 94404 456054 95004 491498
rect 94404 455818 94586 456054
rect 94822 455818 95004 456054
rect 94404 455734 95004 455818
rect 94404 455498 94586 455734
rect 94822 455498 95004 455734
rect 94404 420054 95004 455498
rect 94404 419818 94586 420054
rect 94822 419818 95004 420054
rect 94404 419734 95004 419818
rect 94404 419498 94586 419734
rect 94822 419498 95004 419734
rect 94404 384054 95004 419498
rect 94404 383818 94586 384054
rect 94822 383818 95004 384054
rect 94404 383734 95004 383818
rect 94404 383498 94586 383734
rect 94822 383498 95004 383734
rect 94404 348054 95004 383498
rect 94404 347818 94586 348054
rect 94822 347818 95004 348054
rect 94404 347734 95004 347818
rect 94404 347498 94586 347734
rect 94822 347498 95004 347734
rect 94404 312054 95004 347498
rect 94404 311818 94586 312054
rect 94822 311818 95004 312054
rect 94404 311734 95004 311818
rect 94404 311498 94586 311734
rect 94822 311498 95004 311734
rect 94404 276054 95004 311498
rect 94404 275818 94586 276054
rect 94822 275818 95004 276054
rect 94404 275734 95004 275818
rect 94404 275498 94586 275734
rect 94822 275498 95004 275734
rect 94404 240054 95004 275498
rect 94404 239818 94586 240054
rect 94822 239818 95004 240054
rect 94404 239734 95004 239818
rect 94404 239498 94586 239734
rect 94822 239498 95004 239734
rect 94404 204054 95004 239498
rect 94404 203818 94586 204054
rect 94822 203818 95004 204054
rect 94404 203734 95004 203818
rect 94404 203498 94586 203734
rect 94822 203498 95004 203734
rect 94404 168054 95004 203498
rect 94404 167818 94586 168054
rect 94822 167818 95004 168054
rect 94404 167734 95004 167818
rect 94404 167498 94586 167734
rect 94822 167498 95004 167734
rect 94404 132054 95004 167498
rect 94404 131818 94586 132054
rect 94822 131818 95004 132054
rect 94404 131734 95004 131818
rect 94404 131498 94586 131734
rect 94822 131498 95004 131734
rect 94404 96054 95004 131498
rect 94404 95818 94586 96054
rect 94822 95818 95004 96054
rect 94404 95734 95004 95818
rect 94404 95498 94586 95734
rect 94822 95498 95004 95734
rect 94404 60054 95004 95498
rect 94404 59818 94586 60054
rect 94822 59818 95004 60054
rect 94404 59734 95004 59818
rect 94404 59498 94586 59734
rect 94822 59498 95004 59734
rect 94404 24054 95004 59498
rect 94404 23818 94586 24054
rect 94822 23818 95004 24054
rect 94404 23734 95004 23818
rect 94404 23498 94586 23734
rect 94822 23498 95004 23734
rect 94404 -3166 95004 23498
rect 94404 -3402 94586 -3166
rect 94822 -3402 95004 -3166
rect 94404 -3486 95004 -3402
rect 94404 -3722 94586 -3486
rect 94822 -3722 95004 -3486
rect 94404 -3744 95004 -3722
rect 98004 675654 98604 708982
rect 98004 675418 98186 675654
rect 98422 675418 98604 675654
rect 98004 675334 98604 675418
rect 98004 675098 98186 675334
rect 98422 675098 98604 675334
rect 98004 639654 98604 675098
rect 98004 639418 98186 639654
rect 98422 639418 98604 639654
rect 98004 639334 98604 639418
rect 98004 639098 98186 639334
rect 98422 639098 98604 639334
rect 98004 603654 98604 639098
rect 98004 603418 98186 603654
rect 98422 603418 98604 603654
rect 98004 603334 98604 603418
rect 98004 603098 98186 603334
rect 98422 603098 98604 603334
rect 98004 567654 98604 603098
rect 98004 567418 98186 567654
rect 98422 567418 98604 567654
rect 98004 567334 98604 567418
rect 98004 567098 98186 567334
rect 98422 567098 98604 567334
rect 98004 531654 98604 567098
rect 98004 531418 98186 531654
rect 98422 531418 98604 531654
rect 98004 531334 98604 531418
rect 98004 531098 98186 531334
rect 98422 531098 98604 531334
rect 98004 495654 98604 531098
rect 98004 495418 98186 495654
rect 98422 495418 98604 495654
rect 98004 495334 98604 495418
rect 98004 495098 98186 495334
rect 98422 495098 98604 495334
rect 98004 459654 98604 495098
rect 98004 459418 98186 459654
rect 98422 459418 98604 459654
rect 98004 459334 98604 459418
rect 98004 459098 98186 459334
rect 98422 459098 98604 459334
rect 98004 423654 98604 459098
rect 98004 423418 98186 423654
rect 98422 423418 98604 423654
rect 98004 423334 98604 423418
rect 98004 423098 98186 423334
rect 98422 423098 98604 423334
rect 98004 387654 98604 423098
rect 98004 387418 98186 387654
rect 98422 387418 98604 387654
rect 98004 387334 98604 387418
rect 98004 387098 98186 387334
rect 98422 387098 98604 387334
rect 98004 351654 98604 387098
rect 98004 351418 98186 351654
rect 98422 351418 98604 351654
rect 98004 351334 98604 351418
rect 98004 351098 98186 351334
rect 98422 351098 98604 351334
rect 98004 315654 98604 351098
rect 98004 315418 98186 315654
rect 98422 315418 98604 315654
rect 98004 315334 98604 315418
rect 98004 315098 98186 315334
rect 98422 315098 98604 315334
rect 98004 279654 98604 315098
rect 98004 279418 98186 279654
rect 98422 279418 98604 279654
rect 98004 279334 98604 279418
rect 98004 279098 98186 279334
rect 98422 279098 98604 279334
rect 98004 243654 98604 279098
rect 98004 243418 98186 243654
rect 98422 243418 98604 243654
rect 98004 243334 98604 243418
rect 98004 243098 98186 243334
rect 98422 243098 98604 243334
rect 98004 207654 98604 243098
rect 98004 207418 98186 207654
rect 98422 207418 98604 207654
rect 98004 207334 98604 207418
rect 98004 207098 98186 207334
rect 98422 207098 98604 207334
rect 98004 171654 98604 207098
rect 98004 171418 98186 171654
rect 98422 171418 98604 171654
rect 98004 171334 98604 171418
rect 98004 171098 98186 171334
rect 98422 171098 98604 171334
rect 98004 135654 98604 171098
rect 98004 135418 98186 135654
rect 98422 135418 98604 135654
rect 98004 135334 98604 135418
rect 98004 135098 98186 135334
rect 98422 135098 98604 135334
rect 98004 99654 98604 135098
rect 98004 99418 98186 99654
rect 98422 99418 98604 99654
rect 98004 99334 98604 99418
rect 98004 99098 98186 99334
rect 98422 99098 98604 99334
rect 98004 63654 98604 99098
rect 98004 63418 98186 63654
rect 98422 63418 98604 63654
rect 98004 63334 98604 63418
rect 98004 63098 98186 63334
rect 98422 63098 98604 63334
rect 98004 27654 98604 63098
rect 98004 27418 98186 27654
rect 98422 27418 98604 27654
rect 98004 27334 98604 27418
rect 98004 27098 98186 27334
rect 98422 27098 98604 27334
rect 98004 -5046 98604 27098
rect 98004 -5282 98186 -5046
rect 98422 -5282 98604 -5046
rect 98004 -5366 98604 -5282
rect 98004 -5602 98186 -5366
rect 98422 -5602 98604 -5366
rect 98004 -5624 98604 -5602
rect 101604 679254 102204 710862
rect 119604 710478 120204 711440
rect 119604 710242 119786 710478
rect 120022 710242 120204 710478
rect 119604 710158 120204 710242
rect 119604 709922 119786 710158
rect 120022 709922 120204 710158
rect 116004 708598 116604 709560
rect 116004 708362 116186 708598
rect 116422 708362 116604 708598
rect 116004 708278 116604 708362
rect 116004 708042 116186 708278
rect 116422 708042 116604 708278
rect 112404 706718 113004 707680
rect 112404 706482 112586 706718
rect 112822 706482 113004 706718
rect 112404 706398 113004 706482
rect 112404 706162 112586 706398
rect 112822 706162 113004 706398
rect 101604 679018 101786 679254
rect 102022 679018 102204 679254
rect 101604 678934 102204 679018
rect 101604 678698 101786 678934
rect 102022 678698 102204 678934
rect 101604 643254 102204 678698
rect 101604 643018 101786 643254
rect 102022 643018 102204 643254
rect 101604 642934 102204 643018
rect 101604 642698 101786 642934
rect 102022 642698 102204 642934
rect 101604 607254 102204 642698
rect 101604 607018 101786 607254
rect 102022 607018 102204 607254
rect 101604 606934 102204 607018
rect 101604 606698 101786 606934
rect 102022 606698 102204 606934
rect 101604 571254 102204 606698
rect 101604 571018 101786 571254
rect 102022 571018 102204 571254
rect 101604 570934 102204 571018
rect 101604 570698 101786 570934
rect 102022 570698 102204 570934
rect 101604 535254 102204 570698
rect 101604 535018 101786 535254
rect 102022 535018 102204 535254
rect 101604 534934 102204 535018
rect 101604 534698 101786 534934
rect 102022 534698 102204 534934
rect 101604 499254 102204 534698
rect 101604 499018 101786 499254
rect 102022 499018 102204 499254
rect 101604 498934 102204 499018
rect 101604 498698 101786 498934
rect 102022 498698 102204 498934
rect 101604 463254 102204 498698
rect 101604 463018 101786 463254
rect 102022 463018 102204 463254
rect 101604 462934 102204 463018
rect 101604 462698 101786 462934
rect 102022 462698 102204 462934
rect 101604 427254 102204 462698
rect 101604 427018 101786 427254
rect 102022 427018 102204 427254
rect 101604 426934 102204 427018
rect 101604 426698 101786 426934
rect 102022 426698 102204 426934
rect 101604 391254 102204 426698
rect 101604 391018 101786 391254
rect 102022 391018 102204 391254
rect 101604 390934 102204 391018
rect 101604 390698 101786 390934
rect 102022 390698 102204 390934
rect 101604 355254 102204 390698
rect 101604 355018 101786 355254
rect 102022 355018 102204 355254
rect 101604 354934 102204 355018
rect 101604 354698 101786 354934
rect 102022 354698 102204 354934
rect 101604 319254 102204 354698
rect 101604 319018 101786 319254
rect 102022 319018 102204 319254
rect 101604 318934 102204 319018
rect 101604 318698 101786 318934
rect 102022 318698 102204 318934
rect 101604 283254 102204 318698
rect 101604 283018 101786 283254
rect 102022 283018 102204 283254
rect 101604 282934 102204 283018
rect 101604 282698 101786 282934
rect 102022 282698 102204 282934
rect 101604 247254 102204 282698
rect 101604 247018 101786 247254
rect 102022 247018 102204 247254
rect 101604 246934 102204 247018
rect 101604 246698 101786 246934
rect 102022 246698 102204 246934
rect 101604 211254 102204 246698
rect 101604 211018 101786 211254
rect 102022 211018 102204 211254
rect 101604 210934 102204 211018
rect 101604 210698 101786 210934
rect 102022 210698 102204 210934
rect 101604 175254 102204 210698
rect 101604 175018 101786 175254
rect 102022 175018 102204 175254
rect 101604 174934 102204 175018
rect 101604 174698 101786 174934
rect 102022 174698 102204 174934
rect 101604 139254 102204 174698
rect 101604 139018 101786 139254
rect 102022 139018 102204 139254
rect 101604 138934 102204 139018
rect 101604 138698 101786 138934
rect 102022 138698 102204 138934
rect 101604 103254 102204 138698
rect 101604 103018 101786 103254
rect 102022 103018 102204 103254
rect 101604 102934 102204 103018
rect 101604 102698 101786 102934
rect 102022 102698 102204 102934
rect 101604 67254 102204 102698
rect 101604 67018 101786 67254
rect 102022 67018 102204 67254
rect 101604 66934 102204 67018
rect 101604 66698 101786 66934
rect 102022 66698 102204 66934
rect 101604 31254 102204 66698
rect 101604 31018 101786 31254
rect 102022 31018 102204 31254
rect 101604 30934 102204 31018
rect 101604 30698 101786 30934
rect 102022 30698 102204 30934
rect 83604 -6222 83786 -5986
rect 84022 -6222 84204 -5986
rect 83604 -6306 84204 -6222
rect 83604 -6542 83786 -6306
rect 84022 -6542 84204 -6306
rect 83604 -7504 84204 -6542
rect 101604 -6926 102204 30698
rect 108804 704838 109404 705800
rect 108804 704602 108986 704838
rect 109222 704602 109404 704838
rect 108804 704518 109404 704602
rect 108804 704282 108986 704518
rect 109222 704282 109404 704518
rect 108804 686454 109404 704282
rect 108804 686218 108986 686454
rect 109222 686218 109404 686454
rect 108804 686134 109404 686218
rect 108804 685898 108986 686134
rect 109222 685898 109404 686134
rect 108804 650454 109404 685898
rect 108804 650218 108986 650454
rect 109222 650218 109404 650454
rect 108804 650134 109404 650218
rect 108804 649898 108986 650134
rect 109222 649898 109404 650134
rect 108804 614454 109404 649898
rect 108804 614218 108986 614454
rect 109222 614218 109404 614454
rect 108804 614134 109404 614218
rect 108804 613898 108986 614134
rect 109222 613898 109404 614134
rect 108804 578454 109404 613898
rect 108804 578218 108986 578454
rect 109222 578218 109404 578454
rect 108804 578134 109404 578218
rect 108804 577898 108986 578134
rect 109222 577898 109404 578134
rect 108804 542454 109404 577898
rect 108804 542218 108986 542454
rect 109222 542218 109404 542454
rect 108804 542134 109404 542218
rect 108804 541898 108986 542134
rect 109222 541898 109404 542134
rect 108804 506454 109404 541898
rect 108804 506218 108986 506454
rect 109222 506218 109404 506454
rect 108804 506134 109404 506218
rect 108804 505898 108986 506134
rect 109222 505898 109404 506134
rect 108804 470454 109404 505898
rect 108804 470218 108986 470454
rect 109222 470218 109404 470454
rect 108804 470134 109404 470218
rect 108804 469898 108986 470134
rect 109222 469898 109404 470134
rect 108804 434454 109404 469898
rect 108804 434218 108986 434454
rect 109222 434218 109404 434454
rect 108804 434134 109404 434218
rect 108804 433898 108986 434134
rect 109222 433898 109404 434134
rect 108804 398454 109404 433898
rect 108804 398218 108986 398454
rect 109222 398218 109404 398454
rect 108804 398134 109404 398218
rect 108804 397898 108986 398134
rect 109222 397898 109404 398134
rect 108804 362454 109404 397898
rect 108804 362218 108986 362454
rect 109222 362218 109404 362454
rect 108804 362134 109404 362218
rect 108804 361898 108986 362134
rect 109222 361898 109404 362134
rect 108804 326454 109404 361898
rect 108804 326218 108986 326454
rect 109222 326218 109404 326454
rect 108804 326134 109404 326218
rect 108804 325898 108986 326134
rect 109222 325898 109404 326134
rect 108804 290454 109404 325898
rect 108804 290218 108986 290454
rect 109222 290218 109404 290454
rect 108804 290134 109404 290218
rect 108804 289898 108986 290134
rect 109222 289898 109404 290134
rect 108804 254454 109404 289898
rect 108804 254218 108986 254454
rect 109222 254218 109404 254454
rect 108804 254134 109404 254218
rect 108804 253898 108986 254134
rect 109222 253898 109404 254134
rect 108804 218454 109404 253898
rect 108804 218218 108986 218454
rect 109222 218218 109404 218454
rect 108804 218134 109404 218218
rect 108804 217898 108986 218134
rect 109222 217898 109404 218134
rect 108804 182454 109404 217898
rect 108804 182218 108986 182454
rect 109222 182218 109404 182454
rect 108804 182134 109404 182218
rect 108804 181898 108986 182134
rect 109222 181898 109404 182134
rect 108804 146454 109404 181898
rect 108804 146218 108986 146454
rect 109222 146218 109404 146454
rect 108804 146134 109404 146218
rect 108804 145898 108986 146134
rect 109222 145898 109404 146134
rect 108804 110454 109404 145898
rect 108804 110218 108986 110454
rect 109222 110218 109404 110454
rect 108804 110134 109404 110218
rect 108804 109898 108986 110134
rect 109222 109898 109404 110134
rect 108804 74454 109404 109898
rect 108804 74218 108986 74454
rect 109222 74218 109404 74454
rect 108804 74134 109404 74218
rect 108804 73898 108986 74134
rect 109222 73898 109404 74134
rect 108804 38454 109404 73898
rect 108804 38218 108986 38454
rect 109222 38218 109404 38454
rect 108804 38134 109404 38218
rect 108804 37898 108986 38134
rect 109222 37898 109404 38134
rect 108804 2454 109404 37898
rect 108804 2218 108986 2454
rect 109222 2218 109404 2454
rect 108804 2134 109404 2218
rect 108804 1898 108986 2134
rect 109222 1898 109404 2134
rect 108804 -346 109404 1898
rect 108804 -582 108986 -346
rect 109222 -582 109404 -346
rect 108804 -666 109404 -582
rect 108804 -902 108986 -666
rect 109222 -902 109404 -666
rect 108804 -1864 109404 -902
rect 112404 690054 113004 706162
rect 112404 689818 112586 690054
rect 112822 689818 113004 690054
rect 112404 689734 113004 689818
rect 112404 689498 112586 689734
rect 112822 689498 113004 689734
rect 112404 654054 113004 689498
rect 112404 653818 112586 654054
rect 112822 653818 113004 654054
rect 112404 653734 113004 653818
rect 112404 653498 112586 653734
rect 112822 653498 113004 653734
rect 112404 618054 113004 653498
rect 112404 617818 112586 618054
rect 112822 617818 113004 618054
rect 112404 617734 113004 617818
rect 112404 617498 112586 617734
rect 112822 617498 113004 617734
rect 112404 582054 113004 617498
rect 112404 581818 112586 582054
rect 112822 581818 113004 582054
rect 112404 581734 113004 581818
rect 112404 581498 112586 581734
rect 112822 581498 113004 581734
rect 112404 546054 113004 581498
rect 112404 545818 112586 546054
rect 112822 545818 113004 546054
rect 112404 545734 113004 545818
rect 112404 545498 112586 545734
rect 112822 545498 113004 545734
rect 112404 510054 113004 545498
rect 112404 509818 112586 510054
rect 112822 509818 113004 510054
rect 112404 509734 113004 509818
rect 112404 509498 112586 509734
rect 112822 509498 113004 509734
rect 112404 474054 113004 509498
rect 112404 473818 112586 474054
rect 112822 473818 113004 474054
rect 112404 473734 113004 473818
rect 112404 473498 112586 473734
rect 112822 473498 113004 473734
rect 112404 438054 113004 473498
rect 112404 437818 112586 438054
rect 112822 437818 113004 438054
rect 112404 437734 113004 437818
rect 112404 437498 112586 437734
rect 112822 437498 113004 437734
rect 112404 402054 113004 437498
rect 112404 401818 112586 402054
rect 112822 401818 113004 402054
rect 112404 401734 113004 401818
rect 112404 401498 112586 401734
rect 112822 401498 113004 401734
rect 112404 366054 113004 401498
rect 112404 365818 112586 366054
rect 112822 365818 113004 366054
rect 112404 365734 113004 365818
rect 112404 365498 112586 365734
rect 112822 365498 113004 365734
rect 112404 330054 113004 365498
rect 112404 329818 112586 330054
rect 112822 329818 113004 330054
rect 112404 329734 113004 329818
rect 112404 329498 112586 329734
rect 112822 329498 113004 329734
rect 112404 294054 113004 329498
rect 112404 293818 112586 294054
rect 112822 293818 113004 294054
rect 112404 293734 113004 293818
rect 112404 293498 112586 293734
rect 112822 293498 113004 293734
rect 112404 258054 113004 293498
rect 112404 257818 112586 258054
rect 112822 257818 113004 258054
rect 112404 257734 113004 257818
rect 112404 257498 112586 257734
rect 112822 257498 113004 257734
rect 112404 222054 113004 257498
rect 112404 221818 112586 222054
rect 112822 221818 113004 222054
rect 112404 221734 113004 221818
rect 112404 221498 112586 221734
rect 112822 221498 113004 221734
rect 112404 186054 113004 221498
rect 112404 185818 112586 186054
rect 112822 185818 113004 186054
rect 112404 185734 113004 185818
rect 112404 185498 112586 185734
rect 112822 185498 113004 185734
rect 112404 150054 113004 185498
rect 112404 149818 112586 150054
rect 112822 149818 113004 150054
rect 112404 149734 113004 149818
rect 112404 149498 112586 149734
rect 112822 149498 113004 149734
rect 112404 114054 113004 149498
rect 112404 113818 112586 114054
rect 112822 113818 113004 114054
rect 112404 113734 113004 113818
rect 112404 113498 112586 113734
rect 112822 113498 113004 113734
rect 112404 78054 113004 113498
rect 112404 77818 112586 78054
rect 112822 77818 113004 78054
rect 112404 77734 113004 77818
rect 112404 77498 112586 77734
rect 112822 77498 113004 77734
rect 112404 42054 113004 77498
rect 112404 41818 112586 42054
rect 112822 41818 113004 42054
rect 112404 41734 113004 41818
rect 112404 41498 112586 41734
rect 112822 41498 113004 41734
rect 112404 6054 113004 41498
rect 112404 5818 112586 6054
rect 112822 5818 113004 6054
rect 112404 5734 113004 5818
rect 112404 5498 112586 5734
rect 112822 5498 113004 5734
rect 112404 -2226 113004 5498
rect 112404 -2462 112586 -2226
rect 112822 -2462 113004 -2226
rect 112404 -2546 113004 -2462
rect 112404 -2782 112586 -2546
rect 112822 -2782 113004 -2546
rect 112404 -3744 113004 -2782
rect 116004 693654 116604 708042
rect 116004 693418 116186 693654
rect 116422 693418 116604 693654
rect 116004 693334 116604 693418
rect 116004 693098 116186 693334
rect 116422 693098 116604 693334
rect 116004 657654 116604 693098
rect 116004 657418 116186 657654
rect 116422 657418 116604 657654
rect 116004 657334 116604 657418
rect 116004 657098 116186 657334
rect 116422 657098 116604 657334
rect 116004 621654 116604 657098
rect 116004 621418 116186 621654
rect 116422 621418 116604 621654
rect 116004 621334 116604 621418
rect 116004 621098 116186 621334
rect 116422 621098 116604 621334
rect 116004 585654 116604 621098
rect 116004 585418 116186 585654
rect 116422 585418 116604 585654
rect 116004 585334 116604 585418
rect 116004 585098 116186 585334
rect 116422 585098 116604 585334
rect 116004 549654 116604 585098
rect 116004 549418 116186 549654
rect 116422 549418 116604 549654
rect 116004 549334 116604 549418
rect 116004 549098 116186 549334
rect 116422 549098 116604 549334
rect 116004 513654 116604 549098
rect 116004 513418 116186 513654
rect 116422 513418 116604 513654
rect 116004 513334 116604 513418
rect 116004 513098 116186 513334
rect 116422 513098 116604 513334
rect 116004 477654 116604 513098
rect 116004 477418 116186 477654
rect 116422 477418 116604 477654
rect 116004 477334 116604 477418
rect 116004 477098 116186 477334
rect 116422 477098 116604 477334
rect 116004 441654 116604 477098
rect 116004 441418 116186 441654
rect 116422 441418 116604 441654
rect 116004 441334 116604 441418
rect 116004 441098 116186 441334
rect 116422 441098 116604 441334
rect 116004 405654 116604 441098
rect 116004 405418 116186 405654
rect 116422 405418 116604 405654
rect 116004 405334 116604 405418
rect 116004 405098 116186 405334
rect 116422 405098 116604 405334
rect 116004 369654 116604 405098
rect 116004 369418 116186 369654
rect 116422 369418 116604 369654
rect 116004 369334 116604 369418
rect 116004 369098 116186 369334
rect 116422 369098 116604 369334
rect 116004 333654 116604 369098
rect 116004 333418 116186 333654
rect 116422 333418 116604 333654
rect 116004 333334 116604 333418
rect 116004 333098 116186 333334
rect 116422 333098 116604 333334
rect 116004 297654 116604 333098
rect 116004 297418 116186 297654
rect 116422 297418 116604 297654
rect 116004 297334 116604 297418
rect 116004 297098 116186 297334
rect 116422 297098 116604 297334
rect 116004 261654 116604 297098
rect 116004 261418 116186 261654
rect 116422 261418 116604 261654
rect 116004 261334 116604 261418
rect 116004 261098 116186 261334
rect 116422 261098 116604 261334
rect 116004 225654 116604 261098
rect 116004 225418 116186 225654
rect 116422 225418 116604 225654
rect 116004 225334 116604 225418
rect 116004 225098 116186 225334
rect 116422 225098 116604 225334
rect 116004 189654 116604 225098
rect 116004 189418 116186 189654
rect 116422 189418 116604 189654
rect 116004 189334 116604 189418
rect 116004 189098 116186 189334
rect 116422 189098 116604 189334
rect 116004 153654 116604 189098
rect 116004 153418 116186 153654
rect 116422 153418 116604 153654
rect 116004 153334 116604 153418
rect 116004 153098 116186 153334
rect 116422 153098 116604 153334
rect 116004 117654 116604 153098
rect 116004 117418 116186 117654
rect 116422 117418 116604 117654
rect 116004 117334 116604 117418
rect 116004 117098 116186 117334
rect 116422 117098 116604 117334
rect 116004 81654 116604 117098
rect 116004 81418 116186 81654
rect 116422 81418 116604 81654
rect 116004 81334 116604 81418
rect 116004 81098 116186 81334
rect 116422 81098 116604 81334
rect 116004 45654 116604 81098
rect 116004 45418 116186 45654
rect 116422 45418 116604 45654
rect 116004 45334 116604 45418
rect 116004 45098 116186 45334
rect 116422 45098 116604 45334
rect 116004 9654 116604 45098
rect 116004 9418 116186 9654
rect 116422 9418 116604 9654
rect 116004 9334 116604 9418
rect 116004 9098 116186 9334
rect 116422 9098 116604 9334
rect 116004 -4106 116604 9098
rect 116004 -4342 116186 -4106
rect 116422 -4342 116604 -4106
rect 116004 -4426 116604 -4342
rect 116004 -4662 116186 -4426
rect 116422 -4662 116604 -4426
rect 116004 -5624 116604 -4662
rect 119604 697254 120204 709922
rect 137604 711418 138204 711440
rect 137604 711182 137786 711418
rect 138022 711182 138204 711418
rect 137604 711098 138204 711182
rect 137604 710862 137786 711098
rect 138022 710862 138204 711098
rect 134004 709538 134604 709560
rect 134004 709302 134186 709538
rect 134422 709302 134604 709538
rect 134004 709218 134604 709302
rect 134004 708982 134186 709218
rect 134422 708982 134604 709218
rect 130404 707658 131004 707680
rect 130404 707422 130586 707658
rect 130822 707422 131004 707658
rect 130404 707338 131004 707422
rect 130404 707102 130586 707338
rect 130822 707102 131004 707338
rect 119604 697018 119786 697254
rect 120022 697018 120204 697254
rect 119604 696934 120204 697018
rect 119604 696698 119786 696934
rect 120022 696698 120204 696934
rect 119604 661254 120204 696698
rect 119604 661018 119786 661254
rect 120022 661018 120204 661254
rect 119604 660934 120204 661018
rect 119604 660698 119786 660934
rect 120022 660698 120204 660934
rect 119604 625254 120204 660698
rect 119604 625018 119786 625254
rect 120022 625018 120204 625254
rect 119604 624934 120204 625018
rect 119604 624698 119786 624934
rect 120022 624698 120204 624934
rect 119604 589254 120204 624698
rect 119604 589018 119786 589254
rect 120022 589018 120204 589254
rect 119604 588934 120204 589018
rect 119604 588698 119786 588934
rect 120022 588698 120204 588934
rect 119604 553254 120204 588698
rect 119604 553018 119786 553254
rect 120022 553018 120204 553254
rect 119604 552934 120204 553018
rect 119604 552698 119786 552934
rect 120022 552698 120204 552934
rect 119604 517254 120204 552698
rect 119604 517018 119786 517254
rect 120022 517018 120204 517254
rect 119604 516934 120204 517018
rect 119604 516698 119786 516934
rect 120022 516698 120204 516934
rect 119604 481254 120204 516698
rect 126804 705778 127404 705800
rect 126804 705542 126986 705778
rect 127222 705542 127404 705778
rect 126804 705458 127404 705542
rect 126804 705222 126986 705458
rect 127222 705222 127404 705458
rect 126804 668454 127404 705222
rect 126804 668218 126986 668454
rect 127222 668218 127404 668454
rect 126804 668134 127404 668218
rect 126804 667898 126986 668134
rect 127222 667898 127404 668134
rect 126804 632454 127404 667898
rect 126804 632218 126986 632454
rect 127222 632218 127404 632454
rect 126804 632134 127404 632218
rect 126804 631898 126986 632134
rect 127222 631898 127404 632134
rect 126804 596454 127404 631898
rect 126804 596218 126986 596454
rect 127222 596218 127404 596454
rect 126804 596134 127404 596218
rect 126804 595898 126986 596134
rect 127222 595898 127404 596134
rect 126804 560454 127404 595898
rect 126804 560218 126986 560454
rect 127222 560218 127404 560454
rect 126804 560134 127404 560218
rect 126804 559898 126986 560134
rect 127222 559898 127404 560134
rect 126804 524454 127404 559898
rect 126804 524218 126986 524454
rect 127222 524218 127404 524454
rect 126804 524134 127404 524218
rect 126804 523898 126986 524134
rect 127222 523898 127404 524134
rect 125915 495548 125981 495549
rect 125915 495484 125916 495548
rect 125980 495484 125981 495548
rect 125915 495483 125981 495484
rect 125918 492693 125978 495483
rect 125915 492692 125981 492693
rect 125915 492628 125916 492692
rect 125980 492628 125981 492692
rect 125915 492627 125981 492628
rect 119604 481018 119786 481254
rect 120022 481018 120204 481254
rect 119604 480934 120204 481018
rect 119604 480698 119786 480934
rect 120022 480698 120204 480934
rect 119604 445254 120204 480698
rect 119604 445018 119786 445254
rect 120022 445018 120204 445254
rect 119604 444934 120204 445018
rect 119604 444698 119786 444934
rect 120022 444698 120204 444934
rect 119604 409254 120204 444698
rect 119604 409018 119786 409254
rect 120022 409018 120204 409254
rect 119604 408934 120204 409018
rect 119604 408698 119786 408934
rect 120022 408698 120204 408934
rect 119604 373254 120204 408698
rect 119604 373018 119786 373254
rect 120022 373018 120204 373254
rect 119604 372934 120204 373018
rect 119604 372698 119786 372934
rect 120022 372698 120204 372934
rect 119604 337254 120204 372698
rect 119604 337018 119786 337254
rect 120022 337018 120204 337254
rect 119604 336934 120204 337018
rect 119604 336698 119786 336934
rect 120022 336698 120204 336934
rect 119604 301254 120204 336698
rect 119604 301018 119786 301254
rect 120022 301018 120204 301254
rect 119604 300934 120204 301018
rect 119604 300698 119786 300934
rect 120022 300698 120204 300934
rect 119604 265254 120204 300698
rect 119604 265018 119786 265254
rect 120022 265018 120204 265254
rect 119604 264934 120204 265018
rect 119604 264698 119786 264934
rect 120022 264698 120204 264934
rect 119604 229254 120204 264698
rect 119604 229018 119786 229254
rect 120022 229018 120204 229254
rect 119604 228934 120204 229018
rect 119604 228698 119786 228934
rect 120022 228698 120204 228934
rect 119604 193254 120204 228698
rect 119604 193018 119786 193254
rect 120022 193018 120204 193254
rect 119604 192934 120204 193018
rect 119604 192698 119786 192934
rect 120022 192698 120204 192934
rect 119604 157254 120204 192698
rect 119604 157018 119786 157254
rect 120022 157018 120204 157254
rect 119604 156934 120204 157018
rect 119604 156698 119786 156934
rect 120022 156698 120204 156934
rect 119604 121254 120204 156698
rect 119604 121018 119786 121254
rect 120022 121018 120204 121254
rect 119604 120934 120204 121018
rect 119604 120698 119786 120934
rect 120022 120698 120204 120934
rect 119604 85254 120204 120698
rect 119604 85018 119786 85254
rect 120022 85018 120204 85254
rect 119604 84934 120204 85018
rect 119604 84698 119786 84934
rect 120022 84698 120204 84934
rect 119604 49254 120204 84698
rect 119604 49018 119786 49254
rect 120022 49018 120204 49254
rect 119604 48934 120204 49018
rect 119604 48698 119786 48934
rect 120022 48698 120204 48934
rect 119604 13254 120204 48698
rect 119604 13018 119786 13254
rect 120022 13018 120204 13254
rect 119604 12934 120204 13018
rect 119604 12698 119786 12934
rect 120022 12698 120204 12934
rect 101604 -7162 101786 -6926
rect 102022 -7162 102204 -6926
rect 101604 -7246 102204 -7162
rect 101604 -7482 101786 -7246
rect 102022 -7482 102204 -7246
rect 101604 -7504 102204 -7482
rect 119604 -5986 120204 12698
rect 126804 488454 127404 523898
rect 126804 488218 126986 488454
rect 127222 488218 127404 488454
rect 126804 488134 127404 488218
rect 126804 487898 126986 488134
rect 127222 487898 127404 488134
rect 126804 452454 127404 487898
rect 126804 452218 126986 452454
rect 127222 452218 127404 452454
rect 126804 452134 127404 452218
rect 126804 451898 126986 452134
rect 127222 451898 127404 452134
rect 126804 416454 127404 451898
rect 126804 416218 126986 416454
rect 127222 416218 127404 416454
rect 126804 416134 127404 416218
rect 126804 415898 126986 416134
rect 127222 415898 127404 416134
rect 126804 380454 127404 415898
rect 126804 380218 126986 380454
rect 127222 380218 127404 380454
rect 126804 380134 127404 380218
rect 126804 379898 126986 380134
rect 127222 379898 127404 380134
rect 126804 344454 127404 379898
rect 126804 344218 126986 344454
rect 127222 344218 127404 344454
rect 126804 344134 127404 344218
rect 126804 343898 126986 344134
rect 127222 343898 127404 344134
rect 126804 308454 127404 343898
rect 126804 308218 126986 308454
rect 127222 308218 127404 308454
rect 126804 308134 127404 308218
rect 126804 307898 126986 308134
rect 127222 307898 127404 308134
rect 126804 272454 127404 307898
rect 126804 272218 126986 272454
rect 127222 272218 127404 272454
rect 126804 272134 127404 272218
rect 126804 271898 126986 272134
rect 127222 271898 127404 272134
rect 126804 236454 127404 271898
rect 126804 236218 126986 236454
rect 127222 236218 127404 236454
rect 126804 236134 127404 236218
rect 126804 235898 126986 236134
rect 127222 235898 127404 236134
rect 126804 200454 127404 235898
rect 126804 200218 126986 200454
rect 127222 200218 127404 200454
rect 126804 200134 127404 200218
rect 126804 199898 126986 200134
rect 127222 199898 127404 200134
rect 126804 164454 127404 199898
rect 126804 164218 126986 164454
rect 127222 164218 127404 164454
rect 126804 164134 127404 164218
rect 126804 163898 126986 164134
rect 127222 163898 127404 164134
rect 126804 128454 127404 163898
rect 126804 128218 126986 128454
rect 127222 128218 127404 128454
rect 126804 128134 127404 128218
rect 126804 127898 126986 128134
rect 127222 127898 127404 128134
rect 126804 92454 127404 127898
rect 126804 92218 126986 92454
rect 127222 92218 127404 92454
rect 126804 92134 127404 92218
rect 126804 91898 126986 92134
rect 127222 91898 127404 92134
rect 126804 56454 127404 91898
rect 126804 56218 126986 56454
rect 127222 56218 127404 56454
rect 126804 56134 127404 56218
rect 126804 55898 126986 56134
rect 127222 55898 127404 56134
rect 126804 20454 127404 55898
rect 126804 20218 126986 20454
rect 127222 20218 127404 20454
rect 126804 20134 127404 20218
rect 126804 19898 126986 20134
rect 127222 19898 127404 20134
rect 126804 -1286 127404 19898
rect 126804 -1522 126986 -1286
rect 127222 -1522 127404 -1286
rect 126804 -1606 127404 -1522
rect 126804 -1842 126986 -1606
rect 127222 -1842 127404 -1606
rect 126804 -1864 127404 -1842
rect 130404 672054 131004 707102
rect 132171 700500 132237 700501
rect 132171 700436 132172 700500
rect 132236 700436 132237 700500
rect 132171 700435 132237 700436
rect 131987 685948 132053 685949
rect 131987 685884 131988 685948
rect 132052 685884 132053 685948
rect 131987 685883 132053 685884
rect 130404 671818 130586 672054
rect 130822 671818 131004 672054
rect 130404 671734 131004 671818
rect 130404 671498 130586 671734
rect 130822 671498 131004 671734
rect 130404 636054 131004 671498
rect 131803 639028 131869 639029
rect 131803 638964 131804 639028
rect 131868 638964 131869 639028
rect 131803 638963 131869 638964
rect 130404 635818 130586 636054
rect 130822 635818 131004 636054
rect 130404 635734 131004 635818
rect 130404 635498 130586 635734
rect 130822 635498 131004 635734
rect 130404 600054 131004 635498
rect 130404 599818 130586 600054
rect 130822 599818 131004 600054
rect 130404 599734 131004 599818
rect 130404 599498 130586 599734
rect 130822 599498 131004 599734
rect 130404 564054 131004 599498
rect 130404 563818 130586 564054
rect 130822 563818 131004 564054
rect 130404 563734 131004 563818
rect 130404 563498 130586 563734
rect 130822 563498 131004 563734
rect 130404 528054 131004 563498
rect 130404 527818 130586 528054
rect 130822 527818 131004 528054
rect 130404 527734 131004 527818
rect 130404 527498 130586 527734
rect 130822 527498 131004 527734
rect 130404 492054 131004 527498
rect 130404 491818 130586 492054
rect 130822 491818 131004 492054
rect 130404 491734 131004 491818
rect 130404 491498 130586 491734
rect 130822 491498 131004 491734
rect 130404 456054 131004 491498
rect 130404 455818 130586 456054
rect 130822 455818 131004 456054
rect 130404 455734 131004 455818
rect 130404 455498 130586 455734
rect 130822 455498 131004 455734
rect 130404 420054 131004 455498
rect 130404 419818 130586 420054
rect 130822 419818 131004 420054
rect 130404 419734 131004 419818
rect 130404 419498 130586 419734
rect 130822 419498 131004 419734
rect 130404 384054 131004 419498
rect 130404 383818 130586 384054
rect 130822 383818 131004 384054
rect 130404 383734 131004 383818
rect 130404 383498 130586 383734
rect 130822 383498 131004 383734
rect 130404 348054 131004 383498
rect 130404 347818 130586 348054
rect 130822 347818 131004 348054
rect 130404 347734 131004 347818
rect 130404 347498 130586 347734
rect 130822 347498 131004 347734
rect 130404 312054 131004 347498
rect 130404 311818 130586 312054
rect 130822 311818 131004 312054
rect 130404 311734 131004 311818
rect 130404 311498 130586 311734
rect 130822 311498 131004 311734
rect 130404 276054 131004 311498
rect 130404 275818 130586 276054
rect 130822 275818 131004 276054
rect 130404 275734 131004 275818
rect 130404 275498 130586 275734
rect 130822 275498 131004 275734
rect 130404 240054 131004 275498
rect 130404 239818 130586 240054
rect 130822 239818 131004 240054
rect 130404 239734 131004 239818
rect 130404 239498 130586 239734
rect 130822 239498 131004 239734
rect 130404 204054 131004 239498
rect 130404 203818 130586 204054
rect 130822 203818 131004 204054
rect 130404 203734 131004 203818
rect 130404 203498 130586 203734
rect 130822 203498 131004 203734
rect 130404 168054 131004 203498
rect 130404 167818 130586 168054
rect 130822 167818 131004 168054
rect 130404 167734 131004 167818
rect 130404 167498 130586 167734
rect 130822 167498 131004 167734
rect 130404 132054 131004 167498
rect 131806 134061 131866 638963
rect 131990 135149 132050 685883
rect 132174 137189 132234 700435
rect 132355 700364 132421 700365
rect 132355 700300 132356 700364
rect 132420 700300 132421 700364
rect 132355 700299 132421 700300
rect 132171 137188 132237 137189
rect 132171 137124 132172 137188
rect 132236 137124 132237 137188
rect 132171 137123 132237 137124
rect 132358 136237 132418 700299
rect 133643 697236 133709 697237
rect 133643 697172 133644 697236
rect 133708 697172 133709 697236
rect 133643 697171 133709 697172
rect 133459 650316 133525 650317
rect 133459 650252 133460 650316
rect 133524 650252 133525 650316
rect 133459 650251 133525 650252
rect 133091 603396 133157 603397
rect 133091 603332 133092 603396
rect 133156 603332 133157 603396
rect 133091 603331 133157 603332
rect 132907 200700 132973 200701
rect 132907 200636 132908 200700
rect 132972 200636 132973 200700
rect 132907 200635 132973 200636
rect 132910 176221 132970 200635
rect 132907 176220 132973 176221
rect 132907 176156 132908 176220
rect 132972 176156 132973 176220
rect 132907 176155 132973 176156
rect 133094 172957 133154 603331
rect 133275 592380 133341 592381
rect 133275 592316 133276 592380
rect 133340 592316 133341 592380
rect 133275 592315 133341 592316
rect 133091 172956 133157 172957
rect 133091 172892 133092 172956
rect 133156 172892 133157 172956
rect 133091 172891 133157 172892
rect 132355 136236 132421 136237
rect 132355 136172 132356 136236
rect 132420 136172 132421 136236
rect 132355 136171 132421 136172
rect 131987 135148 132053 135149
rect 131987 135084 131988 135148
rect 132052 135084 132053 135148
rect 131987 135083 132053 135084
rect 131803 134060 131869 134061
rect 131803 133996 131804 134060
rect 131868 133996 131869 134060
rect 131803 133995 131869 133996
rect 133278 132973 133338 592315
rect 133462 174045 133522 650251
rect 133646 175133 133706 697171
rect 134004 675654 134604 708982
rect 134004 675418 134186 675654
rect 134422 675418 134604 675654
rect 134004 675334 134604 675418
rect 134004 675098 134186 675334
rect 134422 675098 134604 675334
rect 134004 639654 134604 675098
rect 134004 639418 134186 639654
rect 134422 639418 134604 639654
rect 134004 639334 134604 639418
rect 134004 639098 134186 639334
rect 134422 639098 134604 639334
rect 134004 603654 134604 639098
rect 134004 603418 134186 603654
rect 134422 603418 134604 603654
rect 134004 603334 134604 603418
rect 134004 603098 134186 603334
rect 134422 603098 134604 603334
rect 134004 567654 134604 603098
rect 134004 567418 134186 567654
rect 134422 567418 134604 567654
rect 134004 567334 134604 567418
rect 134004 567098 134186 567334
rect 134422 567098 134604 567334
rect 134004 531654 134604 567098
rect 134004 531418 134186 531654
rect 134422 531418 134604 531654
rect 134004 531334 134604 531418
rect 134004 531098 134186 531334
rect 134422 531098 134604 531334
rect 134004 495654 134604 531098
rect 134004 495418 134186 495654
rect 134422 495418 134604 495654
rect 134004 495334 134604 495418
rect 134004 495098 134186 495334
rect 134422 495098 134604 495334
rect 134004 459654 134604 495098
rect 134004 459418 134186 459654
rect 134422 459418 134604 459654
rect 134004 459334 134604 459418
rect 134004 459098 134186 459334
rect 134422 459098 134604 459334
rect 134004 423654 134604 459098
rect 134004 423418 134186 423654
rect 134422 423418 134604 423654
rect 134004 423334 134604 423418
rect 134004 423098 134186 423334
rect 134422 423098 134604 423334
rect 134004 387654 134604 423098
rect 134004 387418 134186 387654
rect 134422 387418 134604 387654
rect 134004 387334 134604 387418
rect 134004 387098 134186 387334
rect 134422 387098 134604 387334
rect 134004 351654 134604 387098
rect 134004 351418 134186 351654
rect 134422 351418 134604 351654
rect 134004 351334 134604 351418
rect 134004 351098 134186 351334
rect 134422 351098 134604 351334
rect 134004 315654 134604 351098
rect 134004 315418 134186 315654
rect 134422 315418 134604 315654
rect 134004 315334 134604 315418
rect 134004 315098 134186 315334
rect 134422 315098 134604 315334
rect 134004 279654 134604 315098
rect 134004 279418 134186 279654
rect 134422 279418 134604 279654
rect 134004 279334 134604 279418
rect 134004 279098 134186 279334
rect 134422 279098 134604 279334
rect 134004 243654 134604 279098
rect 134004 243418 134186 243654
rect 134422 243418 134604 243654
rect 134004 243334 134604 243418
rect 134004 243098 134186 243334
rect 134422 243098 134604 243334
rect 134004 207654 134604 243098
rect 134004 207418 134186 207654
rect 134422 207418 134604 207654
rect 134004 207334 134604 207418
rect 134004 207098 134186 207334
rect 134422 207098 134604 207334
rect 133643 175132 133709 175133
rect 133643 175068 133644 175132
rect 133708 175068 133709 175132
rect 133643 175067 133709 175068
rect 133459 174044 133525 174045
rect 133459 173980 133460 174044
rect 133524 173980 133525 174044
rect 133459 173979 133525 173980
rect 134004 171654 134604 207098
rect 134004 171418 134186 171654
rect 134422 171418 134604 171654
rect 134004 171334 134604 171418
rect 134004 171098 134186 171334
rect 134422 171098 134604 171334
rect 134004 135654 134604 171098
rect 134004 135418 134186 135654
rect 134422 135418 134604 135654
rect 134004 135334 134604 135418
rect 134004 135098 134186 135334
rect 134422 135098 134604 135334
rect 133275 132972 133341 132973
rect 133275 132908 133276 132972
rect 133340 132908 133341 132972
rect 133275 132907 133341 132908
rect 130404 131818 130586 132054
rect 130822 131818 131004 132054
rect 130404 131734 131004 131818
rect 130404 131498 130586 131734
rect 130822 131498 131004 131734
rect 130404 96054 131004 131498
rect 130404 95818 130586 96054
rect 130822 95818 131004 96054
rect 130404 95734 131004 95818
rect 130404 95498 130586 95734
rect 130822 95498 131004 95734
rect 130404 60054 131004 95498
rect 130404 59818 130586 60054
rect 130822 59818 131004 60054
rect 130404 59734 131004 59818
rect 130404 59498 130586 59734
rect 130822 59498 131004 59734
rect 130404 24054 131004 59498
rect 130404 23818 130586 24054
rect 130822 23818 131004 24054
rect 130404 23734 131004 23818
rect 130404 23498 130586 23734
rect 130822 23498 131004 23734
rect 130404 -3166 131004 23498
rect 130404 -3402 130586 -3166
rect 130822 -3402 131004 -3166
rect 130404 -3486 131004 -3402
rect 130404 -3722 130586 -3486
rect 130822 -3722 131004 -3486
rect 130404 -3744 131004 -3722
rect 134004 99654 134604 135098
rect 134004 99418 134186 99654
rect 134422 99418 134604 99654
rect 134004 99334 134604 99418
rect 134004 99098 134186 99334
rect 134422 99098 134604 99334
rect 134004 63654 134604 99098
rect 134004 63418 134186 63654
rect 134422 63418 134604 63654
rect 134004 63334 134604 63418
rect 134004 63098 134186 63334
rect 134422 63098 134604 63334
rect 134004 27654 134604 63098
rect 134004 27418 134186 27654
rect 134422 27418 134604 27654
rect 134004 27334 134604 27418
rect 134004 27098 134186 27334
rect 134422 27098 134604 27334
rect 134004 -5046 134604 27098
rect 134004 -5282 134186 -5046
rect 134422 -5282 134604 -5046
rect 134004 -5366 134604 -5282
rect 134004 -5602 134186 -5366
rect 134422 -5602 134604 -5366
rect 134004 -5624 134604 -5602
rect 137604 679254 138204 710862
rect 155604 710478 156204 711440
rect 155604 710242 155786 710478
rect 156022 710242 156204 710478
rect 155604 710158 156204 710242
rect 155604 709922 155786 710158
rect 156022 709922 156204 710158
rect 152004 708598 152604 709560
rect 152004 708362 152186 708598
rect 152422 708362 152604 708598
rect 152004 708278 152604 708362
rect 152004 708042 152186 708278
rect 152422 708042 152604 708278
rect 148404 706718 149004 707680
rect 148404 706482 148586 706718
rect 148822 706482 149004 706718
rect 148404 706398 149004 706482
rect 148404 706162 148586 706398
rect 148822 706162 149004 706398
rect 137604 679018 137786 679254
rect 138022 679018 138204 679254
rect 137604 678934 138204 679018
rect 137604 678698 137786 678934
rect 138022 678698 138204 678934
rect 137604 643254 138204 678698
rect 137604 643018 137786 643254
rect 138022 643018 138204 643254
rect 137604 642934 138204 643018
rect 137604 642698 137786 642934
rect 138022 642698 138204 642934
rect 137604 607254 138204 642698
rect 137604 607018 137786 607254
rect 138022 607018 138204 607254
rect 137604 606934 138204 607018
rect 137604 606698 137786 606934
rect 138022 606698 138204 606934
rect 137604 571254 138204 606698
rect 137604 571018 137786 571254
rect 138022 571018 138204 571254
rect 137604 570934 138204 571018
rect 137604 570698 137786 570934
rect 138022 570698 138204 570934
rect 137604 535254 138204 570698
rect 137604 535018 137786 535254
rect 138022 535018 138204 535254
rect 137604 534934 138204 535018
rect 137604 534698 137786 534934
rect 138022 534698 138204 534934
rect 137604 499254 138204 534698
rect 137604 499018 137786 499254
rect 138022 499018 138204 499254
rect 137604 498934 138204 499018
rect 137604 498698 137786 498934
rect 138022 498698 138204 498934
rect 137604 463254 138204 498698
rect 137604 463018 137786 463254
rect 138022 463018 138204 463254
rect 137604 462934 138204 463018
rect 137604 462698 137786 462934
rect 138022 462698 138204 462934
rect 137604 427254 138204 462698
rect 137604 427018 137786 427254
rect 138022 427018 138204 427254
rect 137604 426934 138204 427018
rect 137604 426698 137786 426934
rect 138022 426698 138204 426934
rect 137604 391254 138204 426698
rect 137604 391018 137786 391254
rect 138022 391018 138204 391254
rect 137604 390934 138204 391018
rect 137604 390698 137786 390934
rect 138022 390698 138204 390934
rect 137604 355254 138204 390698
rect 137604 355018 137786 355254
rect 138022 355018 138204 355254
rect 137604 354934 138204 355018
rect 137604 354698 137786 354934
rect 138022 354698 138204 354934
rect 137604 319254 138204 354698
rect 137604 319018 137786 319254
rect 138022 319018 138204 319254
rect 137604 318934 138204 319018
rect 137604 318698 137786 318934
rect 138022 318698 138204 318934
rect 137604 283254 138204 318698
rect 137604 283018 137786 283254
rect 138022 283018 138204 283254
rect 137604 282934 138204 283018
rect 137604 282698 137786 282934
rect 138022 282698 138204 282934
rect 137604 247254 138204 282698
rect 137604 247018 137786 247254
rect 138022 247018 138204 247254
rect 137604 246934 138204 247018
rect 137604 246698 137786 246934
rect 138022 246698 138204 246934
rect 137604 211254 138204 246698
rect 137604 211018 137786 211254
rect 138022 211018 138204 211254
rect 137604 210934 138204 211018
rect 137604 210698 137786 210934
rect 138022 210698 138204 210934
rect 137604 175254 138204 210698
rect 137604 175018 137786 175254
rect 138022 175018 138204 175254
rect 137604 174934 138204 175018
rect 137604 174698 137786 174934
rect 138022 174698 138204 174934
rect 137604 139254 138204 174698
rect 137604 139018 137786 139254
rect 138022 139018 138204 139254
rect 137604 138934 138204 139018
rect 137604 138698 137786 138934
rect 138022 138698 138204 138934
rect 137604 103254 138204 138698
rect 137604 103018 137786 103254
rect 138022 103018 138204 103254
rect 137604 102934 138204 103018
rect 137604 102698 137786 102934
rect 138022 102698 138204 102934
rect 137604 67254 138204 102698
rect 137604 67018 137786 67254
rect 138022 67018 138204 67254
rect 137604 66934 138204 67018
rect 137604 66698 137786 66934
rect 138022 66698 138204 66934
rect 137604 31254 138204 66698
rect 137604 31018 137786 31254
rect 138022 31018 138204 31254
rect 137604 30934 138204 31018
rect 137604 30698 137786 30934
rect 138022 30698 138204 30934
rect 119604 -6222 119786 -5986
rect 120022 -6222 120204 -5986
rect 119604 -6306 120204 -6222
rect 119604 -6542 119786 -6306
rect 120022 -6542 120204 -6306
rect 119604 -7504 120204 -6542
rect 137604 -6926 138204 30698
rect 144804 704838 145404 705800
rect 144804 704602 144986 704838
rect 145222 704602 145404 704838
rect 144804 704518 145404 704602
rect 144804 704282 144986 704518
rect 145222 704282 145404 704518
rect 144804 686454 145404 704282
rect 144804 686218 144986 686454
rect 145222 686218 145404 686454
rect 144804 686134 145404 686218
rect 144804 685898 144986 686134
rect 145222 685898 145404 686134
rect 144804 650454 145404 685898
rect 144804 650218 144986 650454
rect 145222 650218 145404 650454
rect 144804 650134 145404 650218
rect 144804 649898 144986 650134
rect 145222 649898 145404 650134
rect 144804 614454 145404 649898
rect 144804 614218 144986 614454
rect 145222 614218 145404 614454
rect 144804 614134 145404 614218
rect 144804 613898 144986 614134
rect 145222 613898 145404 614134
rect 144804 578454 145404 613898
rect 144804 578218 144986 578454
rect 145222 578218 145404 578454
rect 144804 578134 145404 578218
rect 144804 577898 144986 578134
rect 145222 577898 145404 578134
rect 144804 542454 145404 577898
rect 144804 542218 144986 542454
rect 145222 542218 145404 542454
rect 144804 542134 145404 542218
rect 144804 541898 144986 542134
rect 145222 541898 145404 542134
rect 144804 506454 145404 541898
rect 144804 506218 144986 506454
rect 145222 506218 145404 506454
rect 144804 506134 145404 506218
rect 144804 505898 144986 506134
rect 145222 505898 145404 506134
rect 144804 470454 145404 505898
rect 144804 470218 144986 470454
rect 145222 470218 145404 470454
rect 144804 470134 145404 470218
rect 144804 469898 144986 470134
rect 145222 469898 145404 470134
rect 144804 434454 145404 469898
rect 144804 434218 144986 434454
rect 145222 434218 145404 434454
rect 144804 434134 145404 434218
rect 144804 433898 144986 434134
rect 145222 433898 145404 434134
rect 144804 398454 145404 433898
rect 144804 398218 144986 398454
rect 145222 398218 145404 398454
rect 144804 398134 145404 398218
rect 144804 397898 144986 398134
rect 145222 397898 145404 398134
rect 144804 362454 145404 397898
rect 144804 362218 144986 362454
rect 145222 362218 145404 362454
rect 144804 362134 145404 362218
rect 144804 361898 144986 362134
rect 145222 361898 145404 362134
rect 144804 326454 145404 361898
rect 144804 326218 144986 326454
rect 145222 326218 145404 326454
rect 144804 326134 145404 326218
rect 144804 325898 144986 326134
rect 145222 325898 145404 326134
rect 144804 290454 145404 325898
rect 144804 290218 144986 290454
rect 145222 290218 145404 290454
rect 144804 290134 145404 290218
rect 144804 289898 144986 290134
rect 145222 289898 145404 290134
rect 144804 254454 145404 289898
rect 144804 254218 144986 254454
rect 145222 254218 145404 254454
rect 144804 254134 145404 254218
rect 144804 253898 144986 254134
rect 145222 253898 145404 254134
rect 144804 218454 145404 253898
rect 144804 218218 144986 218454
rect 145222 218218 145404 218454
rect 144804 218134 145404 218218
rect 144804 217898 144986 218134
rect 145222 217898 145404 218134
rect 144804 182454 145404 217898
rect 144804 182218 144986 182454
rect 145222 182218 145404 182454
rect 144804 182134 145404 182218
rect 144804 181898 144986 182134
rect 145222 181898 145404 182134
rect 144804 146454 145404 181898
rect 144804 146218 144986 146454
rect 145222 146218 145404 146454
rect 144804 146134 145404 146218
rect 144804 145898 144986 146134
rect 145222 145898 145404 146134
rect 144804 110454 145404 145898
rect 144804 110218 144986 110454
rect 145222 110218 145404 110454
rect 144804 110134 145404 110218
rect 144804 109898 144986 110134
rect 145222 109898 145404 110134
rect 144804 74454 145404 109898
rect 144804 74218 144986 74454
rect 145222 74218 145404 74454
rect 144804 74134 145404 74218
rect 144804 73898 144986 74134
rect 145222 73898 145404 74134
rect 144804 38454 145404 73898
rect 144804 38218 144986 38454
rect 145222 38218 145404 38454
rect 144804 38134 145404 38218
rect 144804 37898 144986 38134
rect 145222 37898 145404 38134
rect 144804 2454 145404 37898
rect 144804 2218 144986 2454
rect 145222 2218 145404 2454
rect 144804 2134 145404 2218
rect 144804 1898 144986 2134
rect 145222 1898 145404 2134
rect 144804 -346 145404 1898
rect 144804 -582 144986 -346
rect 145222 -582 145404 -346
rect 144804 -666 145404 -582
rect 144804 -902 144986 -666
rect 145222 -902 145404 -666
rect 144804 -1864 145404 -902
rect 148404 690054 149004 706162
rect 148404 689818 148586 690054
rect 148822 689818 149004 690054
rect 148404 689734 149004 689818
rect 148404 689498 148586 689734
rect 148822 689498 149004 689734
rect 148404 654054 149004 689498
rect 148404 653818 148586 654054
rect 148822 653818 149004 654054
rect 148404 653734 149004 653818
rect 148404 653498 148586 653734
rect 148822 653498 149004 653734
rect 148404 618054 149004 653498
rect 148404 617818 148586 618054
rect 148822 617818 149004 618054
rect 148404 617734 149004 617818
rect 148404 617498 148586 617734
rect 148822 617498 149004 617734
rect 148404 582054 149004 617498
rect 148404 581818 148586 582054
rect 148822 581818 149004 582054
rect 148404 581734 149004 581818
rect 148404 581498 148586 581734
rect 148822 581498 149004 581734
rect 148404 546054 149004 581498
rect 148404 545818 148586 546054
rect 148822 545818 149004 546054
rect 148404 545734 149004 545818
rect 148404 545498 148586 545734
rect 148822 545498 149004 545734
rect 148404 510054 149004 545498
rect 148404 509818 148586 510054
rect 148822 509818 149004 510054
rect 148404 509734 149004 509818
rect 148404 509498 148586 509734
rect 148822 509498 149004 509734
rect 148404 474054 149004 509498
rect 148404 473818 148586 474054
rect 148822 473818 149004 474054
rect 148404 473734 149004 473818
rect 148404 473498 148586 473734
rect 148822 473498 149004 473734
rect 148404 438054 149004 473498
rect 148404 437818 148586 438054
rect 148822 437818 149004 438054
rect 148404 437734 149004 437818
rect 148404 437498 148586 437734
rect 148822 437498 149004 437734
rect 148404 402054 149004 437498
rect 148404 401818 148586 402054
rect 148822 401818 149004 402054
rect 148404 401734 149004 401818
rect 148404 401498 148586 401734
rect 148822 401498 149004 401734
rect 148404 366054 149004 401498
rect 148404 365818 148586 366054
rect 148822 365818 149004 366054
rect 148404 365734 149004 365818
rect 148404 365498 148586 365734
rect 148822 365498 149004 365734
rect 148404 330054 149004 365498
rect 148404 329818 148586 330054
rect 148822 329818 149004 330054
rect 148404 329734 149004 329818
rect 148404 329498 148586 329734
rect 148822 329498 149004 329734
rect 148404 294054 149004 329498
rect 148404 293818 148586 294054
rect 148822 293818 149004 294054
rect 148404 293734 149004 293818
rect 148404 293498 148586 293734
rect 148822 293498 149004 293734
rect 148404 258054 149004 293498
rect 148404 257818 148586 258054
rect 148822 257818 149004 258054
rect 148404 257734 149004 257818
rect 148404 257498 148586 257734
rect 148822 257498 149004 257734
rect 148404 222054 149004 257498
rect 148404 221818 148586 222054
rect 148822 221818 149004 222054
rect 148404 221734 149004 221818
rect 148404 221498 148586 221734
rect 148822 221498 149004 221734
rect 148404 186054 149004 221498
rect 148404 185818 148586 186054
rect 148822 185818 149004 186054
rect 148404 185734 149004 185818
rect 148404 185498 148586 185734
rect 148822 185498 149004 185734
rect 148404 150054 149004 185498
rect 148404 149818 148586 150054
rect 148822 149818 149004 150054
rect 148404 149734 149004 149818
rect 148404 149498 148586 149734
rect 148822 149498 149004 149734
rect 148404 114054 149004 149498
rect 148404 113818 148586 114054
rect 148822 113818 149004 114054
rect 148404 113734 149004 113818
rect 148404 113498 148586 113734
rect 148822 113498 149004 113734
rect 148404 78054 149004 113498
rect 148404 77818 148586 78054
rect 148822 77818 149004 78054
rect 148404 77734 149004 77818
rect 148404 77498 148586 77734
rect 148822 77498 149004 77734
rect 148404 42054 149004 77498
rect 148404 41818 148586 42054
rect 148822 41818 149004 42054
rect 148404 41734 149004 41818
rect 148404 41498 148586 41734
rect 148822 41498 149004 41734
rect 148404 6054 149004 41498
rect 148404 5818 148586 6054
rect 148822 5818 149004 6054
rect 148404 5734 149004 5818
rect 148404 5498 148586 5734
rect 148822 5498 149004 5734
rect 148404 -2226 149004 5498
rect 148404 -2462 148586 -2226
rect 148822 -2462 149004 -2226
rect 148404 -2546 149004 -2462
rect 148404 -2782 148586 -2546
rect 148822 -2782 149004 -2546
rect 148404 -3744 149004 -2782
rect 152004 693654 152604 708042
rect 152004 693418 152186 693654
rect 152422 693418 152604 693654
rect 152004 693334 152604 693418
rect 152004 693098 152186 693334
rect 152422 693098 152604 693334
rect 152004 657654 152604 693098
rect 152004 657418 152186 657654
rect 152422 657418 152604 657654
rect 152004 657334 152604 657418
rect 152004 657098 152186 657334
rect 152422 657098 152604 657334
rect 152004 621654 152604 657098
rect 152004 621418 152186 621654
rect 152422 621418 152604 621654
rect 152004 621334 152604 621418
rect 152004 621098 152186 621334
rect 152422 621098 152604 621334
rect 152004 585654 152604 621098
rect 152004 585418 152186 585654
rect 152422 585418 152604 585654
rect 152004 585334 152604 585418
rect 152004 585098 152186 585334
rect 152422 585098 152604 585334
rect 152004 549654 152604 585098
rect 152004 549418 152186 549654
rect 152422 549418 152604 549654
rect 152004 549334 152604 549418
rect 152004 549098 152186 549334
rect 152422 549098 152604 549334
rect 152004 513654 152604 549098
rect 152004 513418 152186 513654
rect 152422 513418 152604 513654
rect 152004 513334 152604 513418
rect 152004 513098 152186 513334
rect 152422 513098 152604 513334
rect 152004 477654 152604 513098
rect 152004 477418 152186 477654
rect 152422 477418 152604 477654
rect 152004 477334 152604 477418
rect 152004 477098 152186 477334
rect 152422 477098 152604 477334
rect 152004 441654 152604 477098
rect 155604 697254 156204 709922
rect 173604 711418 174204 711440
rect 173604 711182 173786 711418
rect 174022 711182 174204 711418
rect 173604 711098 174204 711182
rect 173604 710862 173786 711098
rect 174022 710862 174204 711098
rect 170004 709538 170604 709560
rect 170004 709302 170186 709538
rect 170422 709302 170604 709538
rect 170004 709218 170604 709302
rect 170004 708982 170186 709218
rect 170422 708982 170604 709218
rect 166404 707658 167004 707680
rect 166404 707422 166586 707658
rect 166822 707422 167004 707658
rect 166404 707338 167004 707422
rect 166404 707102 166586 707338
rect 166822 707102 167004 707338
rect 155604 697018 155786 697254
rect 156022 697018 156204 697254
rect 155604 696934 156204 697018
rect 155604 696698 155786 696934
rect 156022 696698 156204 696934
rect 155604 661254 156204 696698
rect 155604 661018 155786 661254
rect 156022 661018 156204 661254
rect 155604 660934 156204 661018
rect 155604 660698 155786 660934
rect 156022 660698 156204 660934
rect 155604 625254 156204 660698
rect 155604 625018 155786 625254
rect 156022 625018 156204 625254
rect 155604 624934 156204 625018
rect 155604 624698 155786 624934
rect 156022 624698 156204 624934
rect 155604 589254 156204 624698
rect 155604 589018 155786 589254
rect 156022 589018 156204 589254
rect 155604 588934 156204 589018
rect 155604 588698 155786 588934
rect 156022 588698 156204 588934
rect 155604 553254 156204 588698
rect 155604 553018 155786 553254
rect 156022 553018 156204 553254
rect 155604 552934 156204 553018
rect 155604 552698 155786 552934
rect 156022 552698 156204 552934
rect 155604 517254 156204 552698
rect 155604 517018 155786 517254
rect 156022 517018 156204 517254
rect 155604 516934 156204 517018
rect 155604 516698 155786 516934
rect 156022 516698 156204 516934
rect 155604 481254 156204 516698
rect 155604 481018 155786 481254
rect 156022 481018 156204 481254
rect 155604 480934 156204 481018
rect 155604 480698 155786 480934
rect 156022 480698 156204 480934
rect 153331 447268 153397 447269
rect 153331 447204 153332 447268
rect 153396 447204 153397 447268
rect 153331 447203 153397 447204
rect 153334 444413 153394 447203
rect 155604 445254 156204 480698
rect 155604 445018 155786 445254
rect 156022 445018 156204 445254
rect 155604 444934 156204 445018
rect 155604 444698 155786 444934
rect 156022 444698 156204 444934
rect 153331 444412 153397 444413
rect 153331 444348 153332 444412
rect 153396 444348 153397 444412
rect 153331 444347 153397 444348
rect 152004 441418 152186 441654
rect 152422 441418 152604 441654
rect 152004 441334 152604 441418
rect 152004 441098 152186 441334
rect 152422 441098 152604 441334
rect 152004 405654 152604 441098
rect 152004 405418 152186 405654
rect 152422 405418 152604 405654
rect 152004 405334 152604 405418
rect 152004 405098 152186 405334
rect 152422 405098 152604 405334
rect 152004 369654 152604 405098
rect 152004 369418 152186 369654
rect 152422 369418 152604 369654
rect 152004 369334 152604 369418
rect 152004 369098 152186 369334
rect 152422 369098 152604 369334
rect 152004 333654 152604 369098
rect 152004 333418 152186 333654
rect 152422 333418 152604 333654
rect 152004 333334 152604 333418
rect 152004 333098 152186 333334
rect 152422 333098 152604 333334
rect 152004 297654 152604 333098
rect 152004 297418 152186 297654
rect 152422 297418 152604 297654
rect 152004 297334 152604 297418
rect 152004 297098 152186 297334
rect 152422 297098 152604 297334
rect 152004 261654 152604 297098
rect 152004 261418 152186 261654
rect 152422 261418 152604 261654
rect 152004 261334 152604 261418
rect 152004 261098 152186 261334
rect 152422 261098 152604 261334
rect 152004 225654 152604 261098
rect 152004 225418 152186 225654
rect 152422 225418 152604 225654
rect 152004 225334 152604 225418
rect 152004 225098 152186 225334
rect 152422 225098 152604 225334
rect 152004 189654 152604 225098
rect 152004 189418 152186 189654
rect 152422 189418 152604 189654
rect 152004 189334 152604 189418
rect 152004 189098 152186 189334
rect 152422 189098 152604 189334
rect 152004 153654 152604 189098
rect 152004 153418 152186 153654
rect 152422 153418 152604 153654
rect 152004 153334 152604 153418
rect 152004 153098 152186 153334
rect 152422 153098 152604 153334
rect 152004 117654 152604 153098
rect 152004 117418 152186 117654
rect 152422 117418 152604 117654
rect 152004 117334 152604 117418
rect 152004 117098 152186 117334
rect 152422 117098 152604 117334
rect 152004 81654 152604 117098
rect 152004 81418 152186 81654
rect 152422 81418 152604 81654
rect 152004 81334 152604 81418
rect 152004 81098 152186 81334
rect 152422 81098 152604 81334
rect 152004 45654 152604 81098
rect 152004 45418 152186 45654
rect 152422 45418 152604 45654
rect 152004 45334 152604 45418
rect 152004 45098 152186 45334
rect 152422 45098 152604 45334
rect 152004 9654 152604 45098
rect 152004 9418 152186 9654
rect 152422 9418 152604 9654
rect 152004 9334 152604 9418
rect 152004 9098 152186 9334
rect 152422 9098 152604 9334
rect 152004 -4106 152604 9098
rect 152004 -4342 152186 -4106
rect 152422 -4342 152604 -4106
rect 152004 -4426 152604 -4342
rect 152004 -4662 152186 -4426
rect 152422 -4662 152604 -4426
rect 152004 -5624 152604 -4662
rect 155604 409254 156204 444698
rect 155604 409018 155786 409254
rect 156022 409018 156204 409254
rect 155604 408934 156204 409018
rect 155604 408698 155786 408934
rect 156022 408698 156204 408934
rect 155604 373254 156204 408698
rect 155604 373018 155786 373254
rect 156022 373018 156204 373254
rect 155604 372934 156204 373018
rect 155604 372698 155786 372934
rect 156022 372698 156204 372934
rect 155604 337254 156204 372698
rect 155604 337018 155786 337254
rect 156022 337018 156204 337254
rect 155604 336934 156204 337018
rect 155604 336698 155786 336934
rect 156022 336698 156204 336934
rect 155604 301254 156204 336698
rect 155604 301018 155786 301254
rect 156022 301018 156204 301254
rect 155604 300934 156204 301018
rect 155604 300698 155786 300934
rect 156022 300698 156204 300934
rect 155604 265254 156204 300698
rect 155604 265018 155786 265254
rect 156022 265018 156204 265254
rect 155604 264934 156204 265018
rect 155604 264698 155786 264934
rect 156022 264698 156204 264934
rect 155604 229254 156204 264698
rect 155604 229018 155786 229254
rect 156022 229018 156204 229254
rect 155604 228934 156204 229018
rect 155604 228698 155786 228934
rect 156022 228698 156204 228934
rect 155604 193254 156204 228698
rect 155604 193018 155786 193254
rect 156022 193018 156204 193254
rect 155604 192934 156204 193018
rect 155604 192698 155786 192934
rect 156022 192698 156204 192934
rect 155604 157254 156204 192698
rect 155604 157018 155786 157254
rect 156022 157018 156204 157254
rect 155604 156934 156204 157018
rect 155604 156698 155786 156934
rect 156022 156698 156204 156934
rect 155604 121254 156204 156698
rect 155604 121018 155786 121254
rect 156022 121018 156204 121254
rect 155604 120934 156204 121018
rect 155604 120698 155786 120934
rect 156022 120698 156204 120934
rect 155604 85254 156204 120698
rect 155604 85018 155786 85254
rect 156022 85018 156204 85254
rect 155604 84934 156204 85018
rect 155604 84698 155786 84934
rect 156022 84698 156204 84934
rect 155604 49254 156204 84698
rect 155604 49018 155786 49254
rect 156022 49018 156204 49254
rect 155604 48934 156204 49018
rect 155604 48698 155786 48934
rect 156022 48698 156204 48934
rect 155604 13254 156204 48698
rect 155604 13018 155786 13254
rect 156022 13018 156204 13254
rect 155604 12934 156204 13018
rect 155604 12698 155786 12934
rect 156022 12698 156204 12934
rect 137604 -7162 137786 -6926
rect 138022 -7162 138204 -6926
rect 137604 -7246 138204 -7162
rect 137604 -7482 137786 -7246
rect 138022 -7482 138204 -7246
rect 137604 -7504 138204 -7482
rect 155604 -5986 156204 12698
rect 162804 705778 163404 705800
rect 162804 705542 162986 705778
rect 163222 705542 163404 705778
rect 162804 705458 163404 705542
rect 162804 705222 162986 705458
rect 163222 705222 163404 705458
rect 162804 668454 163404 705222
rect 164187 686492 164253 686493
rect 164187 686428 164188 686492
rect 164252 686428 164253 686492
rect 164187 686427 164253 686428
rect 164190 686221 164250 686427
rect 164187 686220 164253 686221
rect 164187 686156 164188 686220
rect 164252 686156 164253 686220
rect 164187 686155 164253 686156
rect 162804 668218 162986 668454
rect 163222 668218 163404 668454
rect 162804 668134 163404 668218
rect 162804 667898 162986 668134
rect 163222 667898 163404 668134
rect 162804 632454 163404 667898
rect 166404 672054 167004 707102
rect 166404 671818 166586 672054
rect 166822 671818 167004 672054
rect 166404 671734 167004 671818
rect 166404 671498 166586 671734
rect 166822 671498 167004 671734
rect 164187 650588 164253 650589
rect 164187 650524 164188 650588
rect 164252 650524 164253 650588
rect 164187 650523 164253 650524
rect 164190 650317 164250 650523
rect 164187 650316 164253 650317
rect 164187 650252 164188 650316
rect 164252 650252 164253 650316
rect 164187 650251 164253 650252
rect 164187 639164 164253 639165
rect 164187 639100 164188 639164
rect 164252 639100 164253 639164
rect 164187 639099 164253 639100
rect 164190 638893 164250 639099
rect 164187 638892 164253 638893
rect 164187 638828 164188 638892
rect 164252 638828 164253 638892
rect 164187 638827 164253 638828
rect 162804 632218 162986 632454
rect 163222 632218 163404 632454
rect 162804 632134 163404 632218
rect 162804 631898 162986 632134
rect 163222 631898 163404 632134
rect 162804 596454 163404 631898
rect 166404 636054 167004 671498
rect 166404 635818 166586 636054
rect 166822 635818 167004 636054
rect 166404 635734 167004 635818
rect 166404 635498 166586 635734
rect 166822 635498 167004 635734
rect 164187 603260 164253 603261
rect 164187 603196 164188 603260
rect 164252 603196 164253 603260
rect 164187 603195 164253 603196
rect 164190 602989 164250 603195
rect 164187 602988 164253 602989
rect 164187 602924 164188 602988
rect 164252 602924 164253 602988
rect 164187 602923 164253 602924
rect 162804 596218 162986 596454
rect 163222 596218 163404 596454
rect 162804 596134 163404 596218
rect 162804 595898 162986 596134
rect 163222 595898 163404 596134
rect 162804 560454 163404 595898
rect 166404 600054 167004 635498
rect 166404 599818 166586 600054
rect 166822 599818 167004 600054
rect 166404 599734 167004 599818
rect 166404 599498 166586 599734
rect 166822 599498 167004 599734
rect 164187 592652 164253 592653
rect 164187 592588 164188 592652
rect 164252 592588 164253 592652
rect 164187 592587 164253 592588
rect 164190 592381 164250 592587
rect 164187 592380 164253 592381
rect 164187 592316 164188 592380
rect 164252 592316 164253 592380
rect 164187 592315 164253 592316
rect 162804 560218 162986 560454
rect 163222 560218 163404 560454
rect 162804 560134 163404 560218
rect 162804 559898 162986 560134
rect 163222 559898 163404 560134
rect 162804 524454 163404 559898
rect 162804 524218 162986 524454
rect 163222 524218 163404 524454
rect 162804 524134 163404 524218
rect 162804 523898 162986 524134
rect 163222 523898 163404 524134
rect 162804 488454 163404 523898
rect 162804 488218 162986 488454
rect 163222 488218 163404 488454
rect 162804 488134 163404 488218
rect 162804 487898 162986 488134
rect 163222 487898 163404 488134
rect 162804 452454 163404 487898
rect 162804 452218 162986 452454
rect 163222 452218 163404 452454
rect 162804 452134 163404 452218
rect 162804 451898 162986 452134
rect 163222 451898 163404 452134
rect 162804 416454 163404 451898
rect 162804 416218 162986 416454
rect 163222 416218 163404 416454
rect 162804 416134 163404 416218
rect 162804 415898 162986 416134
rect 163222 415898 163404 416134
rect 162804 380454 163404 415898
rect 162804 380218 162986 380454
rect 163222 380218 163404 380454
rect 162804 380134 163404 380218
rect 162804 379898 162986 380134
rect 163222 379898 163404 380134
rect 162804 344454 163404 379898
rect 162804 344218 162986 344454
rect 163222 344218 163404 344454
rect 162804 344134 163404 344218
rect 162804 343898 162986 344134
rect 163222 343898 163404 344134
rect 162804 308454 163404 343898
rect 162804 308218 162986 308454
rect 163222 308218 163404 308454
rect 162804 308134 163404 308218
rect 162804 307898 162986 308134
rect 163222 307898 163404 308134
rect 162804 272454 163404 307898
rect 162804 272218 162986 272454
rect 163222 272218 163404 272454
rect 162804 272134 163404 272218
rect 162804 271898 162986 272134
rect 163222 271898 163404 272134
rect 162804 236454 163404 271898
rect 162804 236218 162986 236454
rect 163222 236218 163404 236454
rect 162804 236134 163404 236218
rect 162804 235898 162986 236134
rect 163222 235898 163404 236134
rect 162804 200454 163404 235898
rect 162804 200218 162986 200454
rect 163222 200218 163404 200454
rect 162804 200134 163404 200218
rect 162804 199898 162986 200134
rect 163222 199898 163404 200134
rect 162804 164454 163404 199898
rect 162804 164218 162986 164454
rect 163222 164218 163404 164454
rect 162804 164134 163404 164218
rect 162804 163898 162986 164134
rect 163222 163898 163404 164134
rect 162804 128454 163404 163898
rect 162804 128218 162986 128454
rect 163222 128218 163404 128454
rect 162804 128134 163404 128218
rect 162804 127898 162986 128134
rect 163222 127898 163404 128134
rect 162804 92454 163404 127898
rect 162804 92218 162986 92454
rect 163222 92218 163404 92454
rect 162804 92134 163404 92218
rect 162804 91898 162986 92134
rect 163222 91898 163404 92134
rect 162804 56454 163404 91898
rect 162804 56218 162986 56454
rect 163222 56218 163404 56454
rect 162804 56134 163404 56218
rect 162804 55898 162986 56134
rect 163222 55898 163404 56134
rect 162804 20454 163404 55898
rect 162804 20218 162986 20454
rect 163222 20218 163404 20454
rect 162804 20134 163404 20218
rect 162804 19898 162986 20134
rect 163222 19898 163404 20134
rect 162804 -1286 163404 19898
rect 162804 -1522 162986 -1286
rect 163222 -1522 163404 -1286
rect 162804 -1606 163404 -1522
rect 162804 -1842 162986 -1606
rect 163222 -1842 163404 -1606
rect 162804 -1864 163404 -1842
rect 166404 564054 167004 599498
rect 166404 563818 166586 564054
rect 166822 563818 167004 564054
rect 166404 563734 167004 563818
rect 166404 563498 166586 563734
rect 166822 563498 167004 563734
rect 166404 528054 167004 563498
rect 166404 527818 166586 528054
rect 166822 527818 167004 528054
rect 166404 527734 167004 527818
rect 166404 527498 166586 527734
rect 166822 527498 167004 527734
rect 166404 492054 167004 527498
rect 166404 491818 166586 492054
rect 166822 491818 167004 492054
rect 166404 491734 167004 491818
rect 166404 491498 166586 491734
rect 166822 491498 167004 491734
rect 166404 456054 167004 491498
rect 166404 455818 166586 456054
rect 166822 455818 167004 456054
rect 166404 455734 167004 455818
rect 166404 455498 166586 455734
rect 166822 455498 167004 455734
rect 166404 420054 167004 455498
rect 166404 419818 166586 420054
rect 166822 419818 167004 420054
rect 166404 419734 167004 419818
rect 166404 419498 166586 419734
rect 166822 419498 167004 419734
rect 166404 384054 167004 419498
rect 166404 383818 166586 384054
rect 166822 383818 167004 384054
rect 166404 383734 167004 383818
rect 166404 383498 166586 383734
rect 166822 383498 167004 383734
rect 166404 348054 167004 383498
rect 166404 347818 166586 348054
rect 166822 347818 167004 348054
rect 166404 347734 167004 347818
rect 166404 347498 166586 347734
rect 166822 347498 167004 347734
rect 166404 312054 167004 347498
rect 166404 311818 166586 312054
rect 166822 311818 167004 312054
rect 166404 311734 167004 311818
rect 166404 311498 166586 311734
rect 166822 311498 167004 311734
rect 166404 276054 167004 311498
rect 166404 275818 166586 276054
rect 166822 275818 167004 276054
rect 166404 275734 167004 275818
rect 166404 275498 166586 275734
rect 166822 275498 167004 275734
rect 166404 240054 167004 275498
rect 166404 239818 166586 240054
rect 166822 239818 167004 240054
rect 166404 239734 167004 239818
rect 166404 239498 166586 239734
rect 166822 239498 167004 239734
rect 166404 204054 167004 239498
rect 166404 203818 166586 204054
rect 166822 203818 167004 204054
rect 166404 203734 167004 203818
rect 166404 203498 166586 203734
rect 166822 203498 167004 203734
rect 166404 168054 167004 203498
rect 166404 167818 166586 168054
rect 166822 167818 167004 168054
rect 166404 167734 167004 167818
rect 166404 167498 166586 167734
rect 166822 167498 167004 167734
rect 166404 132054 167004 167498
rect 166404 131818 166586 132054
rect 166822 131818 167004 132054
rect 166404 131734 167004 131818
rect 166404 131498 166586 131734
rect 166822 131498 167004 131734
rect 166404 96054 167004 131498
rect 166404 95818 166586 96054
rect 166822 95818 167004 96054
rect 166404 95734 167004 95818
rect 166404 95498 166586 95734
rect 166822 95498 167004 95734
rect 166404 60054 167004 95498
rect 166404 59818 166586 60054
rect 166822 59818 167004 60054
rect 166404 59734 167004 59818
rect 166404 59498 166586 59734
rect 166822 59498 167004 59734
rect 166404 24054 167004 59498
rect 166404 23818 166586 24054
rect 166822 23818 167004 24054
rect 166404 23734 167004 23818
rect 166404 23498 166586 23734
rect 166822 23498 167004 23734
rect 166404 -3166 167004 23498
rect 166404 -3402 166586 -3166
rect 166822 -3402 167004 -3166
rect 166404 -3486 167004 -3402
rect 166404 -3722 166586 -3486
rect 166822 -3722 167004 -3486
rect 166404 -3744 167004 -3722
rect 170004 675654 170604 708982
rect 170004 675418 170186 675654
rect 170422 675418 170604 675654
rect 170004 675334 170604 675418
rect 170004 675098 170186 675334
rect 170422 675098 170604 675334
rect 170004 639654 170604 675098
rect 170004 639418 170186 639654
rect 170422 639418 170604 639654
rect 170004 639334 170604 639418
rect 170004 639098 170186 639334
rect 170422 639098 170604 639334
rect 170004 603654 170604 639098
rect 170004 603418 170186 603654
rect 170422 603418 170604 603654
rect 170004 603334 170604 603418
rect 170004 603098 170186 603334
rect 170422 603098 170604 603334
rect 170004 567654 170604 603098
rect 170004 567418 170186 567654
rect 170422 567418 170604 567654
rect 170004 567334 170604 567418
rect 170004 567098 170186 567334
rect 170422 567098 170604 567334
rect 170004 531654 170604 567098
rect 170004 531418 170186 531654
rect 170422 531418 170604 531654
rect 170004 531334 170604 531418
rect 170004 531098 170186 531334
rect 170422 531098 170604 531334
rect 170004 495654 170604 531098
rect 170004 495418 170186 495654
rect 170422 495418 170604 495654
rect 170004 495334 170604 495418
rect 170004 495098 170186 495334
rect 170422 495098 170604 495334
rect 170004 459654 170604 495098
rect 170004 459418 170186 459654
rect 170422 459418 170604 459654
rect 170004 459334 170604 459418
rect 170004 459098 170186 459334
rect 170422 459098 170604 459334
rect 170004 423654 170604 459098
rect 170004 423418 170186 423654
rect 170422 423418 170604 423654
rect 170004 423334 170604 423418
rect 170004 423098 170186 423334
rect 170422 423098 170604 423334
rect 170004 387654 170604 423098
rect 170004 387418 170186 387654
rect 170422 387418 170604 387654
rect 170004 387334 170604 387418
rect 170004 387098 170186 387334
rect 170422 387098 170604 387334
rect 170004 351654 170604 387098
rect 170004 351418 170186 351654
rect 170422 351418 170604 351654
rect 170004 351334 170604 351418
rect 170004 351098 170186 351334
rect 170422 351098 170604 351334
rect 170004 315654 170604 351098
rect 170004 315418 170186 315654
rect 170422 315418 170604 315654
rect 170004 315334 170604 315418
rect 170004 315098 170186 315334
rect 170422 315098 170604 315334
rect 170004 279654 170604 315098
rect 170004 279418 170186 279654
rect 170422 279418 170604 279654
rect 170004 279334 170604 279418
rect 170004 279098 170186 279334
rect 170422 279098 170604 279334
rect 170004 243654 170604 279098
rect 170004 243418 170186 243654
rect 170422 243418 170604 243654
rect 170004 243334 170604 243418
rect 170004 243098 170186 243334
rect 170422 243098 170604 243334
rect 170004 207654 170604 243098
rect 170004 207418 170186 207654
rect 170422 207418 170604 207654
rect 170004 207334 170604 207418
rect 170004 207098 170186 207334
rect 170422 207098 170604 207334
rect 170004 171654 170604 207098
rect 170004 171418 170186 171654
rect 170422 171418 170604 171654
rect 170004 171334 170604 171418
rect 170004 171098 170186 171334
rect 170422 171098 170604 171334
rect 170004 135654 170604 171098
rect 170004 135418 170186 135654
rect 170422 135418 170604 135654
rect 170004 135334 170604 135418
rect 170004 135098 170186 135334
rect 170422 135098 170604 135334
rect 170004 99654 170604 135098
rect 170004 99418 170186 99654
rect 170422 99418 170604 99654
rect 170004 99334 170604 99418
rect 170004 99098 170186 99334
rect 170422 99098 170604 99334
rect 170004 63654 170604 99098
rect 170004 63418 170186 63654
rect 170422 63418 170604 63654
rect 170004 63334 170604 63418
rect 170004 63098 170186 63334
rect 170422 63098 170604 63334
rect 170004 27654 170604 63098
rect 170004 27418 170186 27654
rect 170422 27418 170604 27654
rect 170004 27334 170604 27418
rect 170004 27098 170186 27334
rect 170422 27098 170604 27334
rect 170004 -5046 170604 27098
rect 170004 -5282 170186 -5046
rect 170422 -5282 170604 -5046
rect 170004 -5366 170604 -5282
rect 170004 -5602 170186 -5366
rect 170422 -5602 170604 -5366
rect 170004 -5624 170604 -5602
rect 173604 679254 174204 710862
rect 191604 710478 192204 711440
rect 191604 710242 191786 710478
rect 192022 710242 192204 710478
rect 191604 710158 192204 710242
rect 191604 709922 191786 710158
rect 192022 709922 192204 710158
rect 188004 708598 188604 709560
rect 188004 708362 188186 708598
rect 188422 708362 188604 708598
rect 188004 708278 188604 708362
rect 188004 708042 188186 708278
rect 188422 708042 188604 708278
rect 184404 706718 185004 707680
rect 184404 706482 184586 706718
rect 184822 706482 185004 706718
rect 184404 706398 185004 706482
rect 184404 706162 184586 706398
rect 184822 706162 185004 706398
rect 173604 679018 173786 679254
rect 174022 679018 174204 679254
rect 173604 678934 174204 679018
rect 173604 678698 173786 678934
rect 174022 678698 174204 678934
rect 173604 643254 174204 678698
rect 173604 643018 173786 643254
rect 174022 643018 174204 643254
rect 173604 642934 174204 643018
rect 173604 642698 173786 642934
rect 174022 642698 174204 642934
rect 173604 607254 174204 642698
rect 173604 607018 173786 607254
rect 174022 607018 174204 607254
rect 173604 606934 174204 607018
rect 173604 606698 173786 606934
rect 174022 606698 174204 606934
rect 173604 571254 174204 606698
rect 173604 571018 173786 571254
rect 174022 571018 174204 571254
rect 173604 570934 174204 571018
rect 173604 570698 173786 570934
rect 174022 570698 174204 570934
rect 173604 535254 174204 570698
rect 173604 535018 173786 535254
rect 174022 535018 174204 535254
rect 173604 534934 174204 535018
rect 173604 534698 173786 534934
rect 174022 534698 174204 534934
rect 173604 499254 174204 534698
rect 173604 499018 173786 499254
rect 174022 499018 174204 499254
rect 173604 498934 174204 499018
rect 173604 498698 173786 498934
rect 174022 498698 174204 498934
rect 173604 463254 174204 498698
rect 173604 463018 173786 463254
rect 174022 463018 174204 463254
rect 173604 462934 174204 463018
rect 173604 462698 173786 462934
rect 174022 462698 174204 462934
rect 173604 427254 174204 462698
rect 173604 427018 173786 427254
rect 174022 427018 174204 427254
rect 173604 426934 174204 427018
rect 173604 426698 173786 426934
rect 174022 426698 174204 426934
rect 173604 391254 174204 426698
rect 173604 391018 173786 391254
rect 174022 391018 174204 391254
rect 173604 390934 174204 391018
rect 173604 390698 173786 390934
rect 174022 390698 174204 390934
rect 173604 355254 174204 390698
rect 173604 355018 173786 355254
rect 174022 355018 174204 355254
rect 173604 354934 174204 355018
rect 173604 354698 173786 354934
rect 174022 354698 174204 354934
rect 173604 319254 174204 354698
rect 173604 319018 173786 319254
rect 174022 319018 174204 319254
rect 173604 318934 174204 319018
rect 173604 318698 173786 318934
rect 174022 318698 174204 318934
rect 173604 283254 174204 318698
rect 173604 283018 173786 283254
rect 174022 283018 174204 283254
rect 173604 282934 174204 283018
rect 173604 282698 173786 282934
rect 174022 282698 174204 282934
rect 173604 247254 174204 282698
rect 173604 247018 173786 247254
rect 174022 247018 174204 247254
rect 173604 246934 174204 247018
rect 173604 246698 173786 246934
rect 174022 246698 174204 246934
rect 173604 211254 174204 246698
rect 173604 211018 173786 211254
rect 174022 211018 174204 211254
rect 173604 210934 174204 211018
rect 173604 210698 173786 210934
rect 174022 210698 174204 210934
rect 173604 175254 174204 210698
rect 173604 175018 173786 175254
rect 174022 175018 174204 175254
rect 173604 174934 174204 175018
rect 173604 174698 173786 174934
rect 174022 174698 174204 174934
rect 173604 139254 174204 174698
rect 173604 139018 173786 139254
rect 174022 139018 174204 139254
rect 173604 138934 174204 139018
rect 173604 138698 173786 138934
rect 174022 138698 174204 138934
rect 173604 103254 174204 138698
rect 173604 103018 173786 103254
rect 174022 103018 174204 103254
rect 173604 102934 174204 103018
rect 173604 102698 173786 102934
rect 174022 102698 174204 102934
rect 173604 67254 174204 102698
rect 173604 67018 173786 67254
rect 174022 67018 174204 67254
rect 173604 66934 174204 67018
rect 173604 66698 173786 66934
rect 174022 66698 174204 66934
rect 173604 31254 174204 66698
rect 173604 31018 173786 31254
rect 174022 31018 174204 31254
rect 173604 30934 174204 31018
rect 173604 30698 173786 30934
rect 174022 30698 174204 30934
rect 155604 -6222 155786 -5986
rect 156022 -6222 156204 -5986
rect 155604 -6306 156204 -6222
rect 155604 -6542 155786 -6306
rect 156022 -6542 156204 -6306
rect 155604 -7504 156204 -6542
rect 173604 -6926 174204 30698
rect 180804 704838 181404 705800
rect 180804 704602 180986 704838
rect 181222 704602 181404 704838
rect 180804 704518 181404 704602
rect 180804 704282 180986 704518
rect 181222 704282 181404 704518
rect 180804 686454 181404 704282
rect 180804 686218 180986 686454
rect 181222 686218 181404 686454
rect 180804 686134 181404 686218
rect 180804 685898 180986 686134
rect 181222 685898 181404 686134
rect 180804 650454 181404 685898
rect 180804 650218 180986 650454
rect 181222 650218 181404 650454
rect 180804 650134 181404 650218
rect 180804 649898 180986 650134
rect 181222 649898 181404 650134
rect 180804 614454 181404 649898
rect 180804 614218 180986 614454
rect 181222 614218 181404 614454
rect 180804 614134 181404 614218
rect 180804 613898 180986 614134
rect 181222 613898 181404 614134
rect 180804 578454 181404 613898
rect 180804 578218 180986 578454
rect 181222 578218 181404 578454
rect 180804 578134 181404 578218
rect 180804 577898 180986 578134
rect 181222 577898 181404 578134
rect 180804 542454 181404 577898
rect 180804 542218 180986 542454
rect 181222 542218 181404 542454
rect 180804 542134 181404 542218
rect 180804 541898 180986 542134
rect 181222 541898 181404 542134
rect 180804 506454 181404 541898
rect 180804 506218 180986 506454
rect 181222 506218 181404 506454
rect 180804 506134 181404 506218
rect 180804 505898 180986 506134
rect 181222 505898 181404 506134
rect 180804 470454 181404 505898
rect 180804 470218 180986 470454
rect 181222 470218 181404 470454
rect 180804 470134 181404 470218
rect 180804 469898 180986 470134
rect 181222 469898 181404 470134
rect 180804 434454 181404 469898
rect 180804 434218 180986 434454
rect 181222 434218 181404 434454
rect 180804 434134 181404 434218
rect 180804 433898 180986 434134
rect 181222 433898 181404 434134
rect 180804 398454 181404 433898
rect 180804 398218 180986 398454
rect 181222 398218 181404 398454
rect 180804 398134 181404 398218
rect 180804 397898 180986 398134
rect 181222 397898 181404 398134
rect 180804 362454 181404 397898
rect 180804 362218 180986 362454
rect 181222 362218 181404 362454
rect 180804 362134 181404 362218
rect 180804 361898 180986 362134
rect 181222 361898 181404 362134
rect 180804 326454 181404 361898
rect 180804 326218 180986 326454
rect 181222 326218 181404 326454
rect 180804 326134 181404 326218
rect 180804 325898 180986 326134
rect 181222 325898 181404 326134
rect 180804 290454 181404 325898
rect 180804 290218 180986 290454
rect 181222 290218 181404 290454
rect 180804 290134 181404 290218
rect 180804 289898 180986 290134
rect 181222 289898 181404 290134
rect 180804 254454 181404 289898
rect 180804 254218 180986 254454
rect 181222 254218 181404 254454
rect 180804 254134 181404 254218
rect 180804 253898 180986 254134
rect 181222 253898 181404 254134
rect 180804 218454 181404 253898
rect 180804 218218 180986 218454
rect 181222 218218 181404 218454
rect 180804 218134 181404 218218
rect 180804 217898 180986 218134
rect 181222 217898 181404 218134
rect 180804 182454 181404 217898
rect 180804 182218 180986 182454
rect 181222 182218 181404 182454
rect 180804 182134 181404 182218
rect 180804 181898 180986 182134
rect 181222 181898 181404 182134
rect 180804 146454 181404 181898
rect 180804 146218 180986 146454
rect 181222 146218 181404 146454
rect 180804 146134 181404 146218
rect 180804 145898 180986 146134
rect 181222 145898 181404 146134
rect 180804 110454 181404 145898
rect 180804 110218 180986 110454
rect 181222 110218 181404 110454
rect 180804 110134 181404 110218
rect 180804 109898 180986 110134
rect 181222 109898 181404 110134
rect 180804 74454 181404 109898
rect 180804 74218 180986 74454
rect 181222 74218 181404 74454
rect 180804 74134 181404 74218
rect 180804 73898 180986 74134
rect 181222 73898 181404 74134
rect 180804 38454 181404 73898
rect 184404 690054 185004 706162
rect 184404 689818 184586 690054
rect 184822 689818 185004 690054
rect 184404 689734 185004 689818
rect 184404 689498 184586 689734
rect 184822 689498 185004 689734
rect 184404 654054 185004 689498
rect 184404 653818 184586 654054
rect 184822 653818 185004 654054
rect 184404 653734 185004 653818
rect 184404 653498 184586 653734
rect 184822 653498 185004 653734
rect 184404 618054 185004 653498
rect 184404 617818 184586 618054
rect 184822 617818 185004 618054
rect 184404 617734 185004 617818
rect 184404 617498 184586 617734
rect 184822 617498 185004 617734
rect 184404 582054 185004 617498
rect 184404 581818 184586 582054
rect 184822 581818 185004 582054
rect 184404 581734 185004 581818
rect 184404 581498 184586 581734
rect 184822 581498 185004 581734
rect 184404 546054 185004 581498
rect 184404 545818 184586 546054
rect 184822 545818 185004 546054
rect 184404 545734 185004 545818
rect 184404 545498 184586 545734
rect 184822 545498 185004 545734
rect 184404 510054 185004 545498
rect 184404 509818 184586 510054
rect 184822 509818 185004 510054
rect 184404 509734 185004 509818
rect 184404 509498 184586 509734
rect 184822 509498 185004 509734
rect 184404 474054 185004 509498
rect 184404 473818 184586 474054
rect 184822 473818 185004 474054
rect 184404 473734 185004 473818
rect 184404 473498 184586 473734
rect 184822 473498 185004 473734
rect 184404 438054 185004 473498
rect 184404 437818 184586 438054
rect 184822 437818 185004 438054
rect 184404 437734 185004 437818
rect 184404 437498 184586 437734
rect 184822 437498 185004 437734
rect 184404 402054 185004 437498
rect 184404 401818 184586 402054
rect 184822 401818 185004 402054
rect 184404 401734 185004 401818
rect 184404 401498 184586 401734
rect 184822 401498 185004 401734
rect 184404 366054 185004 401498
rect 184404 365818 184586 366054
rect 184822 365818 185004 366054
rect 184404 365734 185004 365818
rect 184404 365498 184586 365734
rect 184822 365498 185004 365734
rect 184404 330054 185004 365498
rect 184404 329818 184586 330054
rect 184822 329818 185004 330054
rect 184404 329734 185004 329818
rect 184404 329498 184586 329734
rect 184822 329498 185004 329734
rect 184404 294054 185004 329498
rect 184404 293818 184586 294054
rect 184822 293818 185004 294054
rect 184404 293734 185004 293818
rect 184404 293498 184586 293734
rect 184822 293498 185004 293734
rect 184404 258054 185004 293498
rect 184404 257818 184586 258054
rect 184822 257818 185004 258054
rect 184404 257734 185004 257818
rect 184404 257498 184586 257734
rect 184822 257498 185004 257734
rect 184404 222054 185004 257498
rect 184404 221818 184586 222054
rect 184822 221818 185004 222054
rect 184404 221734 185004 221818
rect 184404 221498 184586 221734
rect 184822 221498 185004 221734
rect 184404 186054 185004 221498
rect 184404 185818 184586 186054
rect 184822 185818 185004 186054
rect 184404 185734 185004 185818
rect 184404 185498 184586 185734
rect 184822 185498 185004 185734
rect 184404 150054 185004 185498
rect 184404 149818 184586 150054
rect 184822 149818 185004 150054
rect 184404 149734 185004 149818
rect 184404 149498 184586 149734
rect 184822 149498 185004 149734
rect 184404 114054 185004 149498
rect 184404 113818 184586 114054
rect 184822 113818 185004 114054
rect 184404 113734 185004 113818
rect 184404 113498 184586 113734
rect 184822 113498 185004 113734
rect 184404 78054 185004 113498
rect 184404 77818 184586 78054
rect 184822 77818 185004 78054
rect 184404 77734 185004 77818
rect 184404 77498 184586 77734
rect 184822 77498 185004 77734
rect 183691 48108 183757 48109
rect 183691 48044 183692 48108
rect 183756 48044 183757 48108
rect 183691 48043 183757 48044
rect 183694 38725 183754 48043
rect 184404 42054 185004 77498
rect 184404 41818 184586 42054
rect 184822 41818 185004 42054
rect 184404 41734 185004 41818
rect 184404 41498 184586 41734
rect 184822 41498 185004 41734
rect 183691 38724 183757 38725
rect 183691 38660 183692 38724
rect 183756 38660 183757 38724
rect 183691 38659 183757 38660
rect 180804 38218 180986 38454
rect 181222 38218 181404 38454
rect 180804 38134 181404 38218
rect 180804 37898 180986 38134
rect 181222 37898 181404 38134
rect 180804 2454 181404 37898
rect 180804 2218 180986 2454
rect 181222 2218 181404 2454
rect 180804 2134 181404 2218
rect 180804 1898 180986 2134
rect 181222 1898 181404 2134
rect 180804 -346 181404 1898
rect 180804 -582 180986 -346
rect 181222 -582 181404 -346
rect 180804 -666 181404 -582
rect 180804 -902 180986 -666
rect 181222 -902 181404 -666
rect 180804 -1864 181404 -902
rect 184404 6054 185004 41498
rect 184404 5818 184586 6054
rect 184822 5818 185004 6054
rect 184404 5734 185004 5818
rect 184404 5498 184586 5734
rect 184822 5498 185004 5734
rect 184404 -2226 185004 5498
rect 184404 -2462 184586 -2226
rect 184822 -2462 185004 -2226
rect 184404 -2546 185004 -2462
rect 184404 -2782 184586 -2546
rect 184822 -2782 185004 -2546
rect 184404 -3744 185004 -2782
rect 188004 693654 188604 708042
rect 188004 693418 188186 693654
rect 188422 693418 188604 693654
rect 188004 693334 188604 693418
rect 188004 693098 188186 693334
rect 188422 693098 188604 693334
rect 188004 657654 188604 693098
rect 188004 657418 188186 657654
rect 188422 657418 188604 657654
rect 188004 657334 188604 657418
rect 188004 657098 188186 657334
rect 188422 657098 188604 657334
rect 188004 621654 188604 657098
rect 188004 621418 188186 621654
rect 188422 621418 188604 621654
rect 188004 621334 188604 621418
rect 188004 621098 188186 621334
rect 188422 621098 188604 621334
rect 188004 585654 188604 621098
rect 188004 585418 188186 585654
rect 188422 585418 188604 585654
rect 188004 585334 188604 585418
rect 188004 585098 188186 585334
rect 188422 585098 188604 585334
rect 188004 549654 188604 585098
rect 188004 549418 188186 549654
rect 188422 549418 188604 549654
rect 188004 549334 188604 549418
rect 188004 549098 188186 549334
rect 188422 549098 188604 549334
rect 188004 513654 188604 549098
rect 188004 513418 188186 513654
rect 188422 513418 188604 513654
rect 188004 513334 188604 513418
rect 188004 513098 188186 513334
rect 188422 513098 188604 513334
rect 188004 477654 188604 513098
rect 188004 477418 188186 477654
rect 188422 477418 188604 477654
rect 188004 477334 188604 477418
rect 188004 477098 188186 477334
rect 188422 477098 188604 477334
rect 188004 441654 188604 477098
rect 188004 441418 188186 441654
rect 188422 441418 188604 441654
rect 188004 441334 188604 441418
rect 188004 441098 188186 441334
rect 188422 441098 188604 441334
rect 188004 405654 188604 441098
rect 188004 405418 188186 405654
rect 188422 405418 188604 405654
rect 188004 405334 188604 405418
rect 188004 405098 188186 405334
rect 188422 405098 188604 405334
rect 188004 369654 188604 405098
rect 188004 369418 188186 369654
rect 188422 369418 188604 369654
rect 188004 369334 188604 369418
rect 188004 369098 188186 369334
rect 188422 369098 188604 369334
rect 188004 333654 188604 369098
rect 188004 333418 188186 333654
rect 188422 333418 188604 333654
rect 188004 333334 188604 333418
rect 188004 333098 188186 333334
rect 188422 333098 188604 333334
rect 188004 297654 188604 333098
rect 188004 297418 188186 297654
rect 188422 297418 188604 297654
rect 188004 297334 188604 297418
rect 188004 297098 188186 297334
rect 188422 297098 188604 297334
rect 188004 261654 188604 297098
rect 188004 261418 188186 261654
rect 188422 261418 188604 261654
rect 188004 261334 188604 261418
rect 188004 261098 188186 261334
rect 188422 261098 188604 261334
rect 188004 225654 188604 261098
rect 188004 225418 188186 225654
rect 188422 225418 188604 225654
rect 188004 225334 188604 225418
rect 188004 225098 188186 225334
rect 188422 225098 188604 225334
rect 188004 189654 188604 225098
rect 188004 189418 188186 189654
rect 188422 189418 188604 189654
rect 188004 189334 188604 189418
rect 188004 189098 188186 189334
rect 188422 189098 188604 189334
rect 188004 153654 188604 189098
rect 188004 153418 188186 153654
rect 188422 153418 188604 153654
rect 188004 153334 188604 153418
rect 188004 153098 188186 153334
rect 188422 153098 188604 153334
rect 188004 117654 188604 153098
rect 188004 117418 188186 117654
rect 188422 117418 188604 117654
rect 188004 117334 188604 117418
rect 188004 117098 188186 117334
rect 188422 117098 188604 117334
rect 188004 81654 188604 117098
rect 188004 81418 188186 81654
rect 188422 81418 188604 81654
rect 188004 81334 188604 81418
rect 188004 81098 188186 81334
rect 188422 81098 188604 81334
rect 188004 45654 188604 81098
rect 188004 45418 188186 45654
rect 188422 45418 188604 45654
rect 188004 45334 188604 45418
rect 188004 45098 188186 45334
rect 188422 45098 188604 45334
rect 188004 9654 188604 45098
rect 188004 9418 188186 9654
rect 188422 9418 188604 9654
rect 188004 9334 188604 9418
rect 188004 9098 188186 9334
rect 188422 9098 188604 9334
rect 188004 -4106 188604 9098
rect 188004 -4342 188186 -4106
rect 188422 -4342 188604 -4106
rect 188004 -4426 188604 -4342
rect 188004 -4662 188186 -4426
rect 188422 -4662 188604 -4426
rect 188004 -5624 188604 -4662
rect 191604 697254 192204 709922
rect 209604 711418 210204 711440
rect 209604 711182 209786 711418
rect 210022 711182 210204 711418
rect 209604 711098 210204 711182
rect 209604 710862 209786 711098
rect 210022 710862 210204 711098
rect 206004 709538 206604 709560
rect 206004 709302 206186 709538
rect 206422 709302 206604 709538
rect 206004 709218 206604 709302
rect 206004 708982 206186 709218
rect 206422 708982 206604 709218
rect 202404 707658 203004 707680
rect 202404 707422 202586 707658
rect 202822 707422 203004 707658
rect 202404 707338 203004 707422
rect 202404 707102 202586 707338
rect 202822 707102 203004 707338
rect 191604 697018 191786 697254
rect 192022 697018 192204 697254
rect 191604 696934 192204 697018
rect 191604 696698 191786 696934
rect 192022 696698 192204 696934
rect 191604 661254 192204 696698
rect 191604 661018 191786 661254
rect 192022 661018 192204 661254
rect 191604 660934 192204 661018
rect 191604 660698 191786 660934
rect 192022 660698 192204 660934
rect 191604 625254 192204 660698
rect 191604 625018 191786 625254
rect 192022 625018 192204 625254
rect 191604 624934 192204 625018
rect 191604 624698 191786 624934
rect 192022 624698 192204 624934
rect 191604 589254 192204 624698
rect 191604 589018 191786 589254
rect 192022 589018 192204 589254
rect 191604 588934 192204 589018
rect 191604 588698 191786 588934
rect 192022 588698 192204 588934
rect 191604 553254 192204 588698
rect 198804 705778 199404 705800
rect 198804 705542 198986 705778
rect 199222 705542 199404 705778
rect 198804 705458 199404 705542
rect 198804 705222 198986 705458
rect 199222 705222 199404 705458
rect 198804 668454 199404 705222
rect 198804 668218 198986 668454
rect 199222 668218 199404 668454
rect 198804 668134 199404 668218
rect 198804 667898 198986 668134
rect 199222 667898 199404 668134
rect 198804 632454 199404 667898
rect 198804 632218 198986 632454
rect 199222 632218 199404 632454
rect 198804 632134 199404 632218
rect 198804 631898 198986 632134
rect 199222 631898 199404 632134
rect 198804 596454 199404 631898
rect 198804 596218 198986 596454
rect 199222 596218 199404 596454
rect 198804 596134 199404 596218
rect 198804 595898 198986 596134
rect 199222 595898 199404 596134
rect 198804 560454 199404 595898
rect 202404 672054 203004 707102
rect 202404 671818 202586 672054
rect 202822 671818 203004 672054
rect 202404 671734 203004 671818
rect 202404 671498 202586 671734
rect 202822 671498 203004 671734
rect 202404 636054 203004 671498
rect 202404 635818 202586 636054
rect 202822 635818 203004 636054
rect 202404 635734 203004 635818
rect 202404 635498 202586 635734
rect 202822 635498 203004 635734
rect 202404 600054 203004 635498
rect 202404 599818 202586 600054
rect 202822 599818 203004 600054
rect 202404 599734 203004 599818
rect 202404 599498 202586 599734
rect 202822 599498 203004 599734
rect 202404 564054 203004 599498
rect 202404 563818 202586 564054
rect 202822 563818 203004 564054
rect 202404 563734 203004 563818
rect 202404 563498 202586 563734
rect 202822 563498 203004 563734
rect 199699 561780 199765 561781
rect 199699 561716 199700 561780
rect 199764 561716 199765 561780
rect 199699 561715 199765 561716
rect 198804 560218 198986 560454
rect 199222 560218 199404 560454
rect 198804 560134 199404 560218
rect 198804 559898 198986 560134
rect 199222 559898 199404 560134
rect 198595 556748 198661 556749
rect 198595 556684 198596 556748
rect 198660 556684 198661 556748
rect 198595 556683 198661 556684
rect 191604 553018 191786 553254
rect 192022 553018 192204 553254
rect 191604 552934 192204 553018
rect 191604 552698 191786 552934
rect 192022 552698 192204 552934
rect 191604 517254 192204 552698
rect 198411 552124 198477 552125
rect 198411 552060 198412 552124
rect 198476 552060 198477 552124
rect 198411 552059 198477 552060
rect 198227 547908 198293 547909
rect 198227 547844 198228 547908
rect 198292 547844 198293 547908
rect 198227 547843 198293 547844
rect 198043 543828 198109 543829
rect 198043 543764 198044 543828
rect 198108 543764 198109 543828
rect 198043 543763 198109 543764
rect 197859 538524 197925 538525
rect 197859 538460 197860 538524
rect 197924 538460 197925 538524
rect 197859 538459 197925 538460
rect 191604 517018 191786 517254
rect 192022 517018 192204 517254
rect 191604 516934 192204 517018
rect 191604 516698 191786 516934
rect 192022 516698 192204 516934
rect 191604 481254 192204 516698
rect 191604 481018 191786 481254
rect 192022 481018 192204 481254
rect 191604 480934 192204 481018
rect 191604 480698 191786 480934
rect 192022 480698 192204 480934
rect 191604 445254 192204 480698
rect 191604 445018 191786 445254
rect 192022 445018 192204 445254
rect 191604 444934 192204 445018
rect 191604 444698 191786 444934
rect 192022 444698 192204 444934
rect 191604 409254 192204 444698
rect 191604 409018 191786 409254
rect 192022 409018 192204 409254
rect 191604 408934 192204 409018
rect 191604 408698 191786 408934
rect 192022 408698 192204 408934
rect 191604 373254 192204 408698
rect 191604 373018 191786 373254
rect 192022 373018 192204 373254
rect 191604 372934 192204 373018
rect 191604 372698 191786 372934
rect 192022 372698 192204 372934
rect 191604 337254 192204 372698
rect 191604 337018 191786 337254
rect 192022 337018 192204 337254
rect 191604 336934 192204 337018
rect 191604 336698 191786 336934
rect 192022 336698 192204 336934
rect 191604 301254 192204 336698
rect 191604 301018 191786 301254
rect 192022 301018 192204 301254
rect 191604 300934 192204 301018
rect 191604 300698 191786 300934
rect 192022 300698 192204 300934
rect 191604 265254 192204 300698
rect 191604 265018 191786 265254
rect 192022 265018 192204 265254
rect 191604 264934 192204 265018
rect 191604 264698 191786 264934
rect 192022 264698 192204 264934
rect 191604 229254 192204 264698
rect 191604 229018 191786 229254
rect 192022 229018 192204 229254
rect 191604 228934 192204 229018
rect 191604 228698 191786 228934
rect 192022 228698 192204 228934
rect 191604 193254 192204 228698
rect 197862 202605 197922 538459
rect 197859 202604 197925 202605
rect 197859 202540 197860 202604
rect 197924 202540 197925 202604
rect 197859 202539 197925 202540
rect 198046 201653 198106 543763
rect 198230 202333 198290 547843
rect 198227 202332 198293 202333
rect 198227 202268 198228 202332
rect 198292 202268 198293 202332
rect 198227 202267 198293 202268
rect 198414 201925 198474 552059
rect 198411 201924 198477 201925
rect 198411 201860 198412 201924
rect 198476 201860 198477 201924
rect 198411 201859 198477 201860
rect 198598 201789 198658 556683
rect 198804 524454 199404 559898
rect 198804 524218 198986 524454
rect 199222 524218 199404 524454
rect 198804 524134 199404 524218
rect 198804 523898 198986 524134
rect 199222 523898 199404 524134
rect 198804 488454 199404 523898
rect 198804 488218 198986 488454
rect 199222 488218 199404 488454
rect 198804 488134 199404 488218
rect 198804 487898 198986 488134
rect 199222 487898 199404 488134
rect 198804 452454 199404 487898
rect 198804 452218 198986 452454
rect 199222 452218 199404 452454
rect 198804 452134 199404 452218
rect 198804 451898 198986 452134
rect 199222 451898 199404 452134
rect 198804 416454 199404 451898
rect 198804 416218 198986 416454
rect 199222 416218 199404 416454
rect 198804 416134 199404 416218
rect 198804 415898 198986 416134
rect 199222 415898 199404 416134
rect 198804 380454 199404 415898
rect 198804 380218 198986 380454
rect 199222 380218 199404 380454
rect 198804 380134 199404 380218
rect 198804 379898 198986 380134
rect 199222 379898 199404 380134
rect 198804 344454 199404 379898
rect 198804 344218 198986 344454
rect 199222 344218 199404 344454
rect 198804 344134 199404 344218
rect 198804 343898 198986 344134
rect 199222 343898 199404 344134
rect 198804 308454 199404 343898
rect 198804 308218 198986 308454
rect 199222 308218 199404 308454
rect 198804 308134 199404 308218
rect 198804 307898 198986 308134
rect 199222 307898 199404 308134
rect 198804 272454 199404 307898
rect 198804 272218 198986 272454
rect 199222 272218 199404 272454
rect 198804 272134 199404 272218
rect 198804 271898 198986 272134
rect 199222 271898 199404 272134
rect 198804 236454 199404 271898
rect 198804 236218 198986 236454
rect 199222 236218 199404 236454
rect 198804 236134 199404 236218
rect 198804 235898 198986 236134
rect 199222 235898 199404 236134
rect 198595 201788 198661 201789
rect 198595 201724 198596 201788
rect 198660 201724 198661 201788
rect 198595 201723 198661 201724
rect 198043 201652 198109 201653
rect 198043 201588 198044 201652
rect 198108 201588 198109 201652
rect 198043 201587 198109 201588
rect 191604 193018 191786 193254
rect 192022 193018 192204 193254
rect 191604 192934 192204 193018
rect 191604 192698 191786 192934
rect 192022 192698 192204 192934
rect 191604 157254 192204 192698
rect 191604 157018 191786 157254
rect 192022 157018 192204 157254
rect 191604 156934 192204 157018
rect 191604 156698 191786 156934
rect 192022 156698 192204 156934
rect 191604 121254 192204 156698
rect 191604 121018 191786 121254
rect 192022 121018 192204 121254
rect 191604 120934 192204 121018
rect 191604 120698 191786 120934
rect 192022 120698 192204 120934
rect 191604 85254 192204 120698
rect 191604 85018 191786 85254
rect 192022 85018 192204 85254
rect 191604 84934 192204 85018
rect 191604 84698 191786 84934
rect 192022 84698 192204 84934
rect 191604 49254 192204 84698
rect 191604 49018 191786 49254
rect 192022 49018 192204 49254
rect 191604 48934 192204 49018
rect 191604 48698 191786 48934
rect 192022 48698 192204 48934
rect 191604 13254 192204 48698
rect 191604 13018 191786 13254
rect 192022 13018 192204 13254
rect 191604 12934 192204 13018
rect 191604 12698 191786 12934
rect 192022 12698 192204 12934
rect 173604 -7162 173786 -6926
rect 174022 -7162 174204 -6926
rect 173604 -7246 174204 -7162
rect 173604 -7482 173786 -7246
rect 174022 -7482 174204 -7246
rect 173604 -7504 174204 -7482
rect 191604 -5986 192204 12698
rect 198804 200454 199404 235898
rect 199702 202061 199762 561715
rect 202404 528054 203004 563498
rect 202404 527818 202586 528054
rect 202822 527818 203004 528054
rect 202404 527734 203004 527818
rect 202404 527498 202586 527734
rect 202822 527498 203004 527734
rect 202404 492054 203004 527498
rect 202404 491818 202586 492054
rect 202822 491818 203004 492054
rect 202404 491734 203004 491818
rect 202404 491498 202586 491734
rect 202822 491498 203004 491734
rect 202404 456054 203004 491498
rect 202404 455818 202586 456054
rect 202822 455818 203004 456054
rect 202404 455734 203004 455818
rect 202404 455498 202586 455734
rect 202822 455498 203004 455734
rect 202404 420054 203004 455498
rect 202404 419818 202586 420054
rect 202822 419818 203004 420054
rect 202404 419734 203004 419818
rect 202404 419498 202586 419734
rect 202822 419498 203004 419734
rect 202404 384054 203004 419498
rect 202404 383818 202586 384054
rect 202822 383818 203004 384054
rect 202404 383734 203004 383818
rect 202404 383498 202586 383734
rect 202822 383498 203004 383734
rect 202404 348054 203004 383498
rect 202404 347818 202586 348054
rect 202822 347818 203004 348054
rect 202404 347734 203004 347818
rect 202404 347498 202586 347734
rect 202822 347498 203004 347734
rect 202404 312054 203004 347498
rect 202404 311818 202586 312054
rect 202822 311818 203004 312054
rect 202404 311734 203004 311818
rect 202404 311498 202586 311734
rect 202822 311498 203004 311734
rect 202404 276054 203004 311498
rect 202404 275818 202586 276054
rect 202822 275818 203004 276054
rect 202404 275734 203004 275818
rect 202404 275498 202586 275734
rect 202822 275498 203004 275734
rect 202404 240054 203004 275498
rect 202404 239818 202586 240054
rect 202822 239818 203004 240054
rect 202404 239734 203004 239818
rect 202404 239498 202586 239734
rect 202822 239498 203004 239734
rect 202404 204054 203004 239498
rect 202404 203818 202586 204054
rect 202822 203818 203004 204054
rect 202404 203734 203004 203818
rect 202404 203498 202586 203734
rect 202822 203498 203004 203734
rect 199699 202060 199765 202061
rect 199699 201996 199700 202060
rect 199764 201996 199765 202060
rect 199699 201995 199765 201996
rect 198804 200218 198986 200454
rect 199222 200218 199404 200454
rect 198804 200134 199404 200218
rect 198804 199898 198986 200134
rect 199222 199898 199404 200134
rect 198804 164454 199404 199898
rect 198804 164218 198986 164454
rect 199222 164218 199404 164454
rect 198804 164134 199404 164218
rect 198804 163898 198986 164134
rect 199222 163898 199404 164134
rect 198804 128454 199404 163898
rect 198804 128218 198986 128454
rect 199222 128218 199404 128454
rect 198804 128134 199404 128218
rect 198804 127898 198986 128134
rect 199222 127898 199404 128134
rect 198804 92454 199404 127898
rect 198804 92218 198986 92454
rect 199222 92218 199404 92454
rect 198804 92134 199404 92218
rect 198804 91898 198986 92134
rect 199222 91898 199404 92134
rect 198804 56454 199404 91898
rect 198804 56218 198986 56454
rect 199222 56218 199404 56454
rect 198804 56134 199404 56218
rect 198804 55898 198986 56134
rect 199222 55898 199404 56134
rect 198804 20454 199404 55898
rect 198804 20218 198986 20454
rect 199222 20218 199404 20454
rect 198804 20134 199404 20218
rect 198804 19898 198986 20134
rect 199222 19898 199404 20134
rect 198804 -1286 199404 19898
rect 198804 -1522 198986 -1286
rect 199222 -1522 199404 -1286
rect 198804 -1606 199404 -1522
rect 198804 -1842 198986 -1606
rect 199222 -1842 199404 -1606
rect 198804 -1864 199404 -1842
rect 202404 168054 203004 203498
rect 202404 167818 202586 168054
rect 202822 167818 203004 168054
rect 202404 167734 203004 167818
rect 202404 167498 202586 167734
rect 202822 167498 203004 167734
rect 202404 132054 203004 167498
rect 202404 131818 202586 132054
rect 202822 131818 203004 132054
rect 202404 131734 203004 131818
rect 202404 131498 202586 131734
rect 202822 131498 203004 131734
rect 202404 96054 203004 131498
rect 202404 95818 202586 96054
rect 202822 95818 203004 96054
rect 202404 95734 203004 95818
rect 202404 95498 202586 95734
rect 202822 95498 203004 95734
rect 202404 60054 203004 95498
rect 202404 59818 202586 60054
rect 202822 59818 203004 60054
rect 202404 59734 203004 59818
rect 202404 59498 202586 59734
rect 202822 59498 203004 59734
rect 202404 24054 203004 59498
rect 202404 23818 202586 24054
rect 202822 23818 203004 24054
rect 202404 23734 203004 23818
rect 202404 23498 202586 23734
rect 202822 23498 203004 23734
rect 202404 -3166 203004 23498
rect 202404 -3402 202586 -3166
rect 202822 -3402 203004 -3166
rect 202404 -3486 203004 -3402
rect 202404 -3722 202586 -3486
rect 202822 -3722 203004 -3486
rect 202404 -3744 203004 -3722
rect 206004 675654 206604 708982
rect 206004 675418 206186 675654
rect 206422 675418 206604 675654
rect 206004 675334 206604 675418
rect 206004 675098 206186 675334
rect 206422 675098 206604 675334
rect 206004 639654 206604 675098
rect 206004 639418 206186 639654
rect 206422 639418 206604 639654
rect 206004 639334 206604 639418
rect 206004 639098 206186 639334
rect 206422 639098 206604 639334
rect 206004 603654 206604 639098
rect 206004 603418 206186 603654
rect 206422 603418 206604 603654
rect 206004 603334 206604 603418
rect 206004 603098 206186 603334
rect 206422 603098 206604 603334
rect 206004 567654 206604 603098
rect 206004 567418 206186 567654
rect 206422 567418 206604 567654
rect 206004 567334 206604 567418
rect 206004 567098 206186 567334
rect 206422 567098 206604 567334
rect 206004 531654 206604 567098
rect 206004 531418 206186 531654
rect 206422 531418 206604 531654
rect 206004 531334 206604 531418
rect 206004 531098 206186 531334
rect 206422 531098 206604 531334
rect 206004 495654 206604 531098
rect 206004 495418 206186 495654
rect 206422 495418 206604 495654
rect 206004 495334 206604 495418
rect 206004 495098 206186 495334
rect 206422 495098 206604 495334
rect 206004 459654 206604 495098
rect 206004 459418 206186 459654
rect 206422 459418 206604 459654
rect 206004 459334 206604 459418
rect 206004 459098 206186 459334
rect 206422 459098 206604 459334
rect 206004 423654 206604 459098
rect 206004 423418 206186 423654
rect 206422 423418 206604 423654
rect 206004 423334 206604 423418
rect 206004 423098 206186 423334
rect 206422 423098 206604 423334
rect 206004 387654 206604 423098
rect 206004 387418 206186 387654
rect 206422 387418 206604 387654
rect 206004 387334 206604 387418
rect 206004 387098 206186 387334
rect 206422 387098 206604 387334
rect 206004 351654 206604 387098
rect 206004 351418 206186 351654
rect 206422 351418 206604 351654
rect 206004 351334 206604 351418
rect 206004 351098 206186 351334
rect 206422 351098 206604 351334
rect 206004 315654 206604 351098
rect 206004 315418 206186 315654
rect 206422 315418 206604 315654
rect 206004 315334 206604 315418
rect 206004 315098 206186 315334
rect 206422 315098 206604 315334
rect 206004 279654 206604 315098
rect 206004 279418 206186 279654
rect 206422 279418 206604 279654
rect 206004 279334 206604 279418
rect 206004 279098 206186 279334
rect 206422 279098 206604 279334
rect 206004 243654 206604 279098
rect 206004 243418 206186 243654
rect 206422 243418 206604 243654
rect 206004 243334 206604 243418
rect 206004 243098 206186 243334
rect 206422 243098 206604 243334
rect 206004 207654 206604 243098
rect 206004 207418 206186 207654
rect 206422 207418 206604 207654
rect 206004 207334 206604 207418
rect 206004 207098 206186 207334
rect 206422 207098 206604 207334
rect 206004 171654 206604 207098
rect 206004 171418 206186 171654
rect 206422 171418 206604 171654
rect 206004 171334 206604 171418
rect 206004 171098 206186 171334
rect 206422 171098 206604 171334
rect 206004 135654 206604 171098
rect 206004 135418 206186 135654
rect 206422 135418 206604 135654
rect 206004 135334 206604 135418
rect 206004 135098 206186 135334
rect 206422 135098 206604 135334
rect 206004 99654 206604 135098
rect 206004 99418 206186 99654
rect 206422 99418 206604 99654
rect 206004 99334 206604 99418
rect 206004 99098 206186 99334
rect 206422 99098 206604 99334
rect 206004 63654 206604 99098
rect 206004 63418 206186 63654
rect 206422 63418 206604 63654
rect 206004 63334 206604 63418
rect 206004 63098 206186 63334
rect 206422 63098 206604 63334
rect 206004 27654 206604 63098
rect 206004 27418 206186 27654
rect 206422 27418 206604 27654
rect 206004 27334 206604 27418
rect 206004 27098 206186 27334
rect 206422 27098 206604 27334
rect 206004 -5046 206604 27098
rect 206004 -5282 206186 -5046
rect 206422 -5282 206604 -5046
rect 206004 -5366 206604 -5282
rect 206004 -5602 206186 -5366
rect 206422 -5602 206604 -5366
rect 206004 -5624 206604 -5602
rect 209604 679254 210204 710862
rect 227604 710478 228204 711440
rect 227604 710242 227786 710478
rect 228022 710242 228204 710478
rect 227604 710158 228204 710242
rect 227604 709922 227786 710158
rect 228022 709922 228204 710158
rect 224004 708598 224604 709560
rect 224004 708362 224186 708598
rect 224422 708362 224604 708598
rect 224004 708278 224604 708362
rect 224004 708042 224186 708278
rect 224422 708042 224604 708278
rect 220404 706718 221004 707680
rect 220404 706482 220586 706718
rect 220822 706482 221004 706718
rect 220404 706398 221004 706482
rect 220404 706162 220586 706398
rect 220822 706162 221004 706398
rect 209604 679018 209786 679254
rect 210022 679018 210204 679254
rect 209604 678934 210204 679018
rect 209604 678698 209786 678934
rect 210022 678698 210204 678934
rect 209604 643254 210204 678698
rect 209604 643018 209786 643254
rect 210022 643018 210204 643254
rect 209604 642934 210204 643018
rect 209604 642698 209786 642934
rect 210022 642698 210204 642934
rect 209604 607254 210204 642698
rect 209604 607018 209786 607254
rect 210022 607018 210204 607254
rect 209604 606934 210204 607018
rect 209604 606698 209786 606934
rect 210022 606698 210204 606934
rect 209604 571254 210204 606698
rect 209604 571018 209786 571254
rect 210022 571018 210204 571254
rect 209604 570934 210204 571018
rect 209604 570698 209786 570934
rect 210022 570698 210204 570934
rect 209604 535254 210204 570698
rect 209604 535018 209786 535254
rect 210022 535018 210204 535254
rect 209604 534934 210204 535018
rect 209604 534698 209786 534934
rect 210022 534698 210204 534934
rect 209604 499254 210204 534698
rect 209604 499018 209786 499254
rect 210022 499018 210204 499254
rect 209604 498934 210204 499018
rect 209604 498698 209786 498934
rect 210022 498698 210204 498934
rect 209604 463254 210204 498698
rect 209604 463018 209786 463254
rect 210022 463018 210204 463254
rect 209604 462934 210204 463018
rect 209604 462698 209786 462934
rect 210022 462698 210204 462934
rect 209604 427254 210204 462698
rect 209604 427018 209786 427254
rect 210022 427018 210204 427254
rect 209604 426934 210204 427018
rect 209604 426698 209786 426934
rect 210022 426698 210204 426934
rect 209604 391254 210204 426698
rect 209604 391018 209786 391254
rect 210022 391018 210204 391254
rect 209604 390934 210204 391018
rect 209604 390698 209786 390934
rect 210022 390698 210204 390934
rect 209604 355254 210204 390698
rect 209604 355018 209786 355254
rect 210022 355018 210204 355254
rect 209604 354934 210204 355018
rect 209604 354698 209786 354934
rect 210022 354698 210204 354934
rect 209604 319254 210204 354698
rect 209604 319018 209786 319254
rect 210022 319018 210204 319254
rect 209604 318934 210204 319018
rect 209604 318698 209786 318934
rect 210022 318698 210204 318934
rect 209604 283254 210204 318698
rect 209604 283018 209786 283254
rect 210022 283018 210204 283254
rect 209604 282934 210204 283018
rect 209604 282698 209786 282934
rect 210022 282698 210204 282934
rect 209604 247254 210204 282698
rect 209604 247018 209786 247254
rect 210022 247018 210204 247254
rect 209604 246934 210204 247018
rect 209604 246698 209786 246934
rect 210022 246698 210204 246934
rect 209604 211254 210204 246698
rect 209604 211018 209786 211254
rect 210022 211018 210204 211254
rect 209604 210934 210204 211018
rect 209604 210698 209786 210934
rect 210022 210698 210204 210934
rect 209604 175254 210204 210698
rect 209604 175018 209786 175254
rect 210022 175018 210204 175254
rect 209604 174934 210204 175018
rect 209604 174698 209786 174934
rect 210022 174698 210204 174934
rect 209604 139254 210204 174698
rect 209604 139018 209786 139254
rect 210022 139018 210204 139254
rect 209604 138934 210204 139018
rect 209604 138698 209786 138934
rect 210022 138698 210204 138934
rect 209604 103254 210204 138698
rect 209604 103018 209786 103254
rect 210022 103018 210204 103254
rect 209604 102934 210204 103018
rect 209604 102698 209786 102934
rect 210022 102698 210204 102934
rect 209604 67254 210204 102698
rect 209604 67018 209786 67254
rect 210022 67018 210204 67254
rect 209604 66934 210204 67018
rect 209604 66698 209786 66934
rect 210022 66698 210204 66934
rect 209604 31254 210204 66698
rect 209604 31018 209786 31254
rect 210022 31018 210204 31254
rect 209604 30934 210204 31018
rect 209604 30698 209786 30934
rect 210022 30698 210204 30934
rect 191604 -6222 191786 -5986
rect 192022 -6222 192204 -5986
rect 191604 -6306 192204 -6222
rect 191604 -6542 191786 -6306
rect 192022 -6542 192204 -6306
rect 191604 -7504 192204 -6542
rect 209604 -6926 210204 30698
rect 216804 704838 217404 705800
rect 216804 704602 216986 704838
rect 217222 704602 217404 704838
rect 216804 704518 217404 704602
rect 216804 704282 216986 704518
rect 217222 704282 217404 704518
rect 216804 686454 217404 704282
rect 216804 686218 216986 686454
rect 217222 686218 217404 686454
rect 216804 686134 217404 686218
rect 216804 685898 216986 686134
rect 217222 685898 217404 686134
rect 216804 650454 217404 685898
rect 216804 650218 216986 650454
rect 217222 650218 217404 650454
rect 216804 650134 217404 650218
rect 216804 649898 216986 650134
rect 217222 649898 217404 650134
rect 216804 614454 217404 649898
rect 216804 614218 216986 614454
rect 217222 614218 217404 614454
rect 216804 614134 217404 614218
rect 216804 613898 216986 614134
rect 217222 613898 217404 614134
rect 216804 578454 217404 613898
rect 216804 578218 216986 578454
rect 217222 578218 217404 578454
rect 216804 578134 217404 578218
rect 216804 577898 216986 578134
rect 217222 577898 217404 578134
rect 216804 542454 217404 577898
rect 216804 542218 216986 542454
rect 217222 542218 217404 542454
rect 216804 542134 217404 542218
rect 216804 541898 216986 542134
rect 217222 541898 217404 542134
rect 216804 506454 217404 541898
rect 216804 506218 216986 506454
rect 217222 506218 217404 506454
rect 216804 506134 217404 506218
rect 216804 505898 216986 506134
rect 217222 505898 217404 506134
rect 216804 470454 217404 505898
rect 216804 470218 216986 470454
rect 217222 470218 217404 470454
rect 216804 470134 217404 470218
rect 216804 469898 216986 470134
rect 217222 469898 217404 470134
rect 216804 434454 217404 469898
rect 216804 434218 216986 434454
rect 217222 434218 217404 434454
rect 216804 434134 217404 434218
rect 216804 433898 216986 434134
rect 217222 433898 217404 434134
rect 216804 398454 217404 433898
rect 216804 398218 216986 398454
rect 217222 398218 217404 398454
rect 216804 398134 217404 398218
rect 216804 397898 216986 398134
rect 217222 397898 217404 398134
rect 216804 362454 217404 397898
rect 216804 362218 216986 362454
rect 217222 362218 217404 362454
rect 216804 362134 217404 362218
rect 216804 361898 216986 362134
rect 217222 361898 217404 362134
rect 216804 326454 217404 361898
rect 216804 326218 216986 326454
rect 217222 326218 217404 326454
rect 216804 326134 217404 326218
rect 216804 325898 216986 326134
rect 217222 325898 217404 326134
rect 216804 290454 217404 325898
rect 216804 290218 216986 290454
rect 217222 290218 217404 290454
rect 216804 290134 217404 290218
rect 216804 289898 216986 290134
rect 217222 289898 217404 290134
rect 216804 254454 217404 289898
rect 216804 254218 216986 254454
rect 217222 254218 217404 254454
rect 216804 254134 217404 254218
rect 216804 253898 216986 254134
rect 217222 253898 217404 254134
rect 216804 218454 217404 253898
rect 216804 218218 216986 218454
rect 217222 218218 217404 218454
rect 216804 218134 217404 218218
rect 216804 217898 216986 218134
rect 217222 217898 217404 218134
rect 216804 182454 217404 217898
rect 216804 182218 216986 182454
rect 217222 182218 217404 182454
rect 216804 182134 217404 182218
rect 216804 181898 216986 182134
rect 217222 181898 217404 182134
rect 216804 146454 217404 181898
rect 216804 146218 216986 146454
rect 217222 146218 217404 146454
rect 216804 146134 217404 146218
rect 216804 145898 216986 146134
rect 217222 145898 217404 146134
rect 216804 110454 217404 145898
rect 216804 110218 216986 110454
rect 217222 110218 217404 110454
rect 216804 110134 217404 110218
rect 216804 109898 216986 110134
rect 217222 109898 217404 110134
rect 216804 74454 217404 109898
rect 216804 74218 216986 74454
rect 217222 74218 217404 74454
rect 216804 74134 217404 74218
rect 216804 73898 216986 74134
rect 217222 73898 217404 74134
rect 216804 38454 217404 73898
rect 216804 38218 216986 38454
rect 217222 38218 217404 38454
rect 216804 38134 217404 38218
rect 216804 37898 216986 38134
rect 217222 37898 217404 38134
rect 216804 2454 217404 37898
rect 216804 2218 216986 2454
rect 217222 2218 217404 2454
rect 216804 2134 217404 2218
rect 216804 1898 216986 2134
rect 217222 1898 217404 2134
rect 216804 -346 217404 1898
rect 216804 -582 216986 -346
rect 217222 -582 217404 -346
rect 216804 -666 217404 -582
rect 216804 -902 216986 -666
rect 217222 -902 217404 -666
rect 216804 -1864 217404 -902
rect 220404 690054 221004 706162
rect 220404 689818 220586 690054
rect 220822 689818 221004 690054
rect 220404 689734 221004 689818
rect 220404 689498 220586 689734
rect 220822 689498 221004 689734
rect 220404 654054 221004 689498
rect 220404 653818 220586 654054
rect 220822 653818 221004 654054
rect 220404 653734 221004 653818
rect 220404 653498 220586 653734
rect 220822 653498 221004 653734
rect 220404 618054 221004 653498
rect 220404 617818 220586 618054
rect 220822 617818 221004 618054
rect 220404 617734 221004 617818
rect 220404 617498 220586 617734
rect 220822 617498 221004 617734
rect 220404 582054 221004 617498
rect 220404 581818 220586 582054
rect 220822 581818 221004 582054
rect 220404 581734 221004 581818
rect 220404 581498 220586 581734
rect 220822 581498 221004 581734
rect 220404 546054 221004 581498
rect 220404 545818 220586 546054
rect 220822 545818 221004 546054
rect 220404 545734 221004 545818
rect 220404 545498 220586 545734
rect 220822 545498 221004 545734
rect 220404 510054 221004 545498
rect 220404 509818 220586 510054
rect 220822 509818 221004 510054
rect 220404 509734 221004 509818
rect 220404 509498 220586 509734
rect 220822 509498 221004 509734
rect 220404 474054 221004 509498
rect 220404 473818 220586 474054
rect 220822 473818 221004 474054
rect 220404 473734 221004 473818
rect 220404 473498 220586 473734
rect 220822 473498 221004 473734
rect 220404 438054 221004 473498
rect 220404 437818 220586 438054
rect 220822 437818 221004 438054
rect 220404 437734 221004 437818
rect 220404 437498 220586 437734
rect 220822 437498 221004 437734
rect 220404 402054 221004 437498
rect 220404 401818 220586 402054
rect 220822 401818 221004 402054
rect 220404 401734 221004 401818
rect 220404 401498 220586 401734
rect 220822 401498 221004 401734
rect 220404 366054 221004 401498
rect 220404 365818 220586 366054
rect 220822 365818 221004 366054
rect 220404 365734 221004 365818
rect 220404 365498 220586 365734
rect 220822 365498 221004 365734
rect 220404 330054 221004 365498
rect 220404 329818 220586 330054
rect 220822 329818 221004 330054
rect 220404 329734 221004 329818
rect 220404 329498 220586 329734
rect 220822 329498 221004 329734
rect 220404 294054 221004 329498
rect 220404 293818 220586 294054
rect 220822 293818 221004 294054
rect 220404 293734 221004 293818
rect 220404 293498 220586 293734
rect 220822 293498 221004 293734
rect 220404 258054 221004 293498
rect 220404 257818 220586 258054
rect 220822 257818 221004 258054
rect 220404 257734 221004 257818
rect 220404 257498 220586 257734
rect 220822 257498 221004 257734
rect 220404 222054 221004 257498
rect 220404 221818 220586 222054
rect 220822 221818 221004 222054
rect 220404 221734 221004 221818
rect 220404 221498 220586 221734
rect 220822 221498 221004 221734
rect 220404 186054 221004 221498
rect 220404 185818 220586 186054
rect 220822 185818 221004 186054
rect 220404 185734 221004 185818
rect 220404 185498 220586 185734
rect 220822 185498 221004 185734
rect 220404 150054 221004 185498
rect 220404 149818 220586 150054
rect 220822 149818 221004 150054
rect 220404 149734 221004 149818
rect 220404 149498 220586 149734
rect 220822 149498 221004 149734
rect 220404 114054 221004 149498
rect 220404 113818 220586 114054
rect 220822 113818 221004 114054
rect 220404 113734 221004 113818
rect 220404 113498 220586 113734
rect 220822 113498 221004 113734
rect 220404 78054 221004 113498
rect 220404 77818 220586 78054
rect 220822 77818 221004 78054
rect 220404 77734 221004 77818
rect 220404 77498 220586 77734
rect 220822 77498 221004 77734
rect 220404 42054 221004 77498
rect 220404 41818 220586 42054
rect 220822 41818 221004 42054
rect 220404 41734 221004 41818
rect 220404 41498 220586 41734
rect 220822 41498 221004 41734
rect 220404 6054 221004 41498
rect 220404 5818 220586 6054
rect 220822 5818 221004 6054
rect 220404 5734 221004 5818
rect 220404 5498 220586 5734
rect 220822 5498 221004 5734
rect 220404 -2226 221004 5498
rect 220404 -2462 220586 -2226
rect 220822 -2462 221004 -2226
rect 220404 -2546 221004 -2462
rect 220404 -2782 220586 -2546
rect 220822 -2782 221004 -2546
rect 220404 -3744 221004 -2782
rect 224004 693654 224604 708042
rect 224004 693418 224186 693654
rect 224422 693418 224604 693654
rect 224004 693334 224604 693418
rect 224004 693098 224186 693334
rect 224422 693098 224604 693334
rect 224004 657654 224604 693098
rect 224004 657418 224186 657654
rect 224422 657418 224604 657654
rect 224004 657334 224604 657418
rect 224004 657098 224186 657334
rect 224422 657098 224604 657334
rect 224004 621654 224604 657098
rect 224004 621418 224186 621654
rect 224422 621418 224604 621654
rect 224004 621334 224604 621418
rect 224004 621098 224186 621334
rect 224422 621098 224604 621334
rect 224004 585654 224604 621098
rect 224004 585418 224186 585654
rect 224422 585418 224604 585654
rect 224004 585334 224604 585418
rect 224004 585098 224186 585334
rect 224422 585098 224604 585334
rect 224004 549654 224604 585098
rect 224004 549418 224186 549654
rect 224422 549418 224604 549654
rect 224004 549334 224604 549418
rect 224004 549098 224186 549334
rect 224422 549098 224604 549334
rect 224004 513654 224604 549098
rect 224004 513418 224186 513654
rect 224422 513418 224604 513654
rect 224004 513334 224604 513418
rect 224004 513098 224186 513334
rect 224422 513098 224604 513334
rect 224004 477654 224604 513098
rect 224004 477418 224186 477654
rect 224422 477418 224604 477654
rect 224004 477334 224604 477418
rect 224004 477098 224186 477334
rect 224422 477098 224604 477334
rect 224004 441654 224604 477098
rect 224004 441418 224186 441654
rect 224422 441418 224604 441654
rect 224004 441334 224604 441418
rect 224004 441098 224186 441334
rect 224422 441098 224604 441334
rect 224004 405654 224604 441098
rect 224004 405418 224186 405654
rect 224422 405418 224604 405654
rect 224004 405334 224604 405418
rect 224004 405098 224186 405334
rect 224422 405098 224604 405334
rect 224004 369654 224604 405098
rect 224004 369418 224186 369654
rect 224422 369418 224604 369654
rect 224004 369334 224604 369418
rect 224004 369098 224186 369334
rect 224422 369098 224604 369334
rect 224004 333654 224604 369098
rect 224004 333418 224186 333654
rect 224422 333418 224604 333654
rect 224004 333334 224604 333418
rect 224004 333098 224186 333334
rect 224422 333098 224604 333334
rect 224004 297654 224604 333098
rect 224004 297418 224186 297654
rect 224422 297418 224604 297654
rect 224004 297334 224604 297418
rect 224004 297098 224186 297334
rect 224422 297098 224604 297334
rect 224004 261654 224604 297098
rect 224004 261418 224186 261654
rect 224422 261418 224604 261654
rect 224004 261334 224604 261418
rect 224004 261098 224186 261334
rect 224422 261098 224604 261334
rect 224004 225654 224604 261098
rect 224004 225418 224186 225654
rect 224422 225418 224604 225654
rect 224004 225334 224604 225418
rect 224004 225098 224186 225334
rect 224422 225098 224604 225334
rect 224004 189654 224604 225098
rect 224004 189418 224186 189654
rect 224422 189418 224604 189654
rect 224004 189334 224604 189418
rect 224004 189098 224186 189334
rect 224422 189098 224604 189334
rect 224004 153654 224604 189098
rect 224004 153418 224186 153654
rect 224422 153418 224604 153654
rect 224004 153334 224604 153418
rect 224004 153098 224186 153334
rect 224422 153098 224604 153334
rect 224004 117654 224604 153098
rect 224004 117418 224186 117654
rect 224422 117418 224604 117654
rect 224004 117334 224604 117418
rect 224004 117098 224186 117334
rect 224422 117098 224604 117334
rect 224004 81654 224604 117098
rect 224004 81418 224186 81654
rect 224422 81418 224604 81654
rect 224004 81334 224604 81418
rect 224004 81098 224186 81334
rect 224422 81098 224604 81334
rect 224004 45654 224604 81098
rect 224004 45418 224186 45654
rect 224422 45418 224604 45654
rect 224004 45334 224604 45418
rect 224004 45098 224186 45334
rect 224422 45098 224604 45334
rect 224004 9654 224604 45098
rect 224004 9418 224186 9654
rect 224422 9418 224604 9654
rect 224004 9334 224604 9418
rect 224004 9098 224186 9334
rect 224422 9098 224604 9334
rect 224004 -4106 224604 9098
rect 224004 -4342 224186 -4106
rect 224422 -4342 224604 -4106
rect 224004 -4426 224604 -4342
rect 224004 -4662 224186 -4426
rect 224422 -4662 224604 -4426
rect 224004 -5624 224604 -4662
rect 227604 697254 228204 709922
rect 245604 711418 246204 711440
rect 245604 711182 245786 711418
rect 246022 711182 246204 711418
rect 245604 711098 246204 711182
rect 245604 710862 245786 711098
rect 246022 710862 246204 711098
rect 242004 709538 242604 709560
rect 242004 709302 242186 709538
rect 242422 709302 242604 709538
rect 242004 709218 242604 709302
rect 242004 708982 242186 709218
rect 242422 708982 242604 709218
rect 238404 707658 239004 707680
rect 238404 707422 238586 707658
rect 238822 707422 239004 707658
rect 238404 707338 239004 707422
rect 238404 707102 238586 707338
rect 238822 707102 239004 707338
rect 227604 697018 227786 697254
rect 228022 697018 228204 697254
rect 227604 696934 228204 697018
rect 227604 696698 227786 696934
rect 228022 696698 228204 696934
rect 227604 661254 228204 696698
rect 227604 661018 227786 661254
rect 228022 661018 228204 661254
rect 227604 660934 228204 661018
rect 227604 660698 227786 660934
rect 228022 660698 228204 660934
rect 227604 625254 228204 660698
rect 227604 625018 227786 625254
rect 228022 625018 228204 625254
rect 227604 624934 228204 625018
rect 227604 624698 227786 624934
rect 228022 624698 228204 624934
rect 227604 589254 228204 624698
rect 227604 589018 227786 589254
rect 228022 589018 228204 589254
rect 227604 588934 228204 589018
rect 227604 588698 227786 588934
rect 228022 588698 228204 588934
rect 227604 553254 228204 588698
rect 227604 553018 227786 553254
rect 228022 553018 228204 553254
rect 227604 552934 228204 553018
rect 227604 552698 227786 552934
rect 228022 552698 228204 552934
rect 227604 517254 228204 552698
rect 227604 517018 227786 517254
rect 228022 517018 228204 517254
rect 227604 516934 228204 517018
rect 227604 516698 227786 516934
rect 228022 516698 228204 516934
rect 227604 481254 228204 516698
rect 227604 481018 227786 481254
rect 228022 481018 228204 481254
rect 227604 480934 228204 481018
rect 227604 480698 227786 480934
rect 228022 480698 228204 480934
rect 227604 445254 228204 480698
rect 227604 445018 227786 445254
rect 228022 445018 228204 445254
rect 227604 444934 228204 445018
rect 227604 444698 227786 444934
rect 228022 444698 228204 444934
rect 227604 409254 228204 444698
rect 227604 409018 227786 409254
rect 228022 409018 228204 409254
rect 227604 408934 228204 409018
rect 227604 408698 227786 408934
rect 228022 408698 228204 408934
rect 227604 373254 228204 408698
rect 227604 373018 227786 373254
rect 228022 373018 228204 373254
rect 227604 372934 228204 373018
rect 227604 372698 227786 372934
rect 228022 372698 228204 372934
rect 227604 337254 228204 372698
rect 227604 337018 227786 337254
rect 228022 337018 228204 337254
rect 227604 336934 228204 337018
rect 227604 336698 227786 336934
rect 228022 336698 228204 336934
rect 227604 301254 228204 336698
rect 227604 301018 227786 301254
rect 228022 301018 228204 301254
rect 227604 300934 228204 301018
rect 227604 300698 227786 300934
rect 228022 300698 228204 300934
rect 227604 265254 228204 300698
rect 227604 265018 227786 265254
rect 228022 265018 228204 265254
rect 227604 264934 228204 265018
rect 227604 264698 227786 264934
rect 228022 264698 228204 264934
rect 227604 229254 228204 264698
rect 227604 229018 227786 229254
rect 228022 229018 228204 229254
rect 227604 228934 228204 229018
rect 227604 228698 227786 228934
rect 228022 228698 228204 228934
rect 227604 193254 228204 228698
rect 227604 193018 227786 193254
rect 228022 193018 228204 193254
rect 227604 192934 228204 193018
rect 227604 192698 227786 192934
rect 228022 192698 228204 192934
rect 227604 157254 228204 192698
rect 227604 157018 227786 157254
rect 228022 157018 228204 157254
rect 227604 156934 228204 157018
rect 227604 156698 227786 156934
rect 228022 156698 228204 156934
rect 227604 121254 228204 156698
rect 227604 121018 227786 121254
rect 228022 121018 228204 121254
rect 227604 120934 228204 121018
rect 227604 120698 227786 120934
rect 228022 120698 228204 120934
rect 227604 85254 228204 120698
rect 227604 85018 227786 85254
rect 228022 85018 228204 85254
rect 227604 84934 228204 85018
rect 227604 84698 227786 84934
rect 228022 84698 228204 84934
rect 227604 49254 228204 84698
rect 227604 49018 227786 49254
rect 228022 49018 228204 49254
rect 227604 48934 228204 49018
rect 227604 48698 227786 48934
rect 228022 48698 228204 48934
rect 227604 13254 228204 48698
rect 227604 13018 227786 13254
rect 228022 13018 228204 13254
rect 227604 12934 228204 13018
rect 227604 12698 227786 12934
rect 228022 12698 228204 12934
rect 209604 -7162 209786 -6926
rect 210022 -7162 210204 -6926
rect 209604 -7246 210204 -7162
rect 209604 -7482 209786 -7246
rect 210022 -7482 210204 -7246
rect 209604 -7504 210204 -7482
rect 227604 -5986 228204 12698
rect 234804 705778 235404 705800
rect 234804 705542 234986 705778
rect 235222 705542 235404 705778
rect 234804 705458 235404 705542
rect 234804 705222 234986 705458
rect 235222 705222 235404 705458
rect 234804 668454 235404 705222
rect 234804 668218 234986 668454
rect 235222 668218 235404 668454
rect 234804 668134 235404 668218
rect 234804 667898 234986 668134
rect 235222 667898 235404 668134
rect 234804 632454 235404 667898
rect 234804 632218 234986 632454
rect 235222 632218 235404 632454
rect 234804 632134 235404 632218
rect 234804 631898 234986 632134
rect 235222 631898 235404 632134
rect 234804 596454 235404 631898
rect 234804 596218 234986 596454
rect 235222 596218 235404 596454
rect 234804 596134 235404 596218
rect 234804 595898 234986 596134
rect 235222 595898 235404 596134
rect 234804 560454 235404 595898
rect 234804 560218 234986 560454
rect 235222 560218 235404 560454
rect 234804 560134 235404 560218
rect 234804 559898 234986 560134
rect 235222 559898 235404 560134
rect 234804 524454 235404 559898
rect 234804 524218 234986 524454
rect 235222 524218 235404 524454
rect 234804 524134 235404 524218
rect 234804 523898 234986 524134
rect 235222 523898 235404 524134
rect 234804 488454 235404 523898
rect 234804 488218 234986 488454
rect 235222 488218 235404 488454
rect 234804 488134 235404 488218
rect 234804 487898 234986 488134
rect 235222 487898 235404 488134
rect 234804 452454 235404 487898
rect 234804 452218 234986 452454
rect 235222 452218 235404 452454
rect 234804 452134 235404 452218
rect 234804 451898 234986 452134
rect 235222 451898 235404 452134
rect 234804 416454 235404 451898
rect 234804 416218 234986 416454
rect 235222 416218 235404 416454
rect 234804 416134 235404 416218
rect 234804 415898 234986 416134
rect 235222 415898 235404 416134
rect 234804 380454 235404 415898
rect 234804 380218 234986 380454
rect 235222 380218 235404 380454
rect 234804 380134 235404 380218
rect 234804 379898 234986 380134
rect 235222 379898 235404 380134
rect 234804 344454 235404 379898
rect 234804 344218 234986 344454
rect 235222 344218 235404 344454
rect 234804 344134 235404 344218
rect 234804 343898 234986 344134
rect 235222 343898 235404 344134
rect 234804 308454 235404 343898
rect 234804 308218 234986 308454
rect 235222 308218 235404 308454
rect 234804 308134 235404 308218
rect 234804 307898 234986 308134
rect 235222 307898 235404 308134
rect 234804 272454 235404 307898
rect 234804 272218 234986 272454
rect 235222 272218 235404 272454
rect 234804 272134 235404 272218
rect 234804 271898 234986 272134
rect 235222 271898 235404 272134
rect 234804 236454 235404 271898
rect 234804 236218 234986 236454
rect 235222 236218 235404 236454
rect 234804 236134 235404 236218
rect 234804 235898 234986 236134
rect 235222 235898 235404 236134
rect 234804 200454 235404 235898
rect 234804 200218 234986 200454
rect 235222 200218 235404 200454
rect 234804 200134 235404 200218
rect 234804 199898 234986 200134
rect 235222 199898 235404 200134
rect 234804 164454 235404 199898
rect 234804 164218 234986 164454
rect 235222 164218 235404 164454
rect 234804 164134 235404 164218
rect 234804 163898 234986 164134
rect 235222 163898 235404 164134
rect 234804 128454 235404 163898
rect 234804 128218 234986 128454
rect 235222 128218 235404 128454
rect 234804 128134 235404 128218
rect 234804 127898 234986 128134
rect 235222 127898 235404 128134
rect 234804 92454 235404 127898
rect 234804 92218 234986 92454
rect 235222 92218 235404 92454
rect 234804 92134 235404 92218
rect 234804 91898 234986 92134
rect 235222 91898 235404 92134
rect 234804 56454 235404 91898
rect 234804 56218 234986 56454
rect 235222 56218 235404 56454
rect 234804 56134 235404 56218
rect 234804 55898 234986 56134
rect 235222 55898 235404 56134
rect 234804 20454 235404 55898
rect 234804 20218 234986 20454
rect 235222 20218 235404 20454
rect 234804 20134 235404 20218
rect 234804 19898 234986 20134
rect 235222 19898 235404 20134
rect 234804 -1286 235404 19898
rect 234804 -1522 234986 -1286
rect 235222 -1522 235404 -1286
rect 234804 -1606 235404 -1522
rect 234804 -1842 234986 -1606
rect 235222 -1842 235404 -1606
rect 234804 -1864 235404 -1842
rect 238404 672054 239004 707102
rect 238404 671818 238586 672054
rect 238822 671818 239004 672054
rect 238404 671734 239004 671818
rect 238404 671498 238586 671734
rect 238822 671498 239004 671734
rect 238404 636054 239004 671498
rect 238404 635818 238586 636054
rect 238822 635818 239004 636054
rect 238404 635734 239004 635818
rect 238404 635498 238586 635734
rect 238822 635498 239004 635734
rect 238404 600054 239004 635498
rect 238404 599818 238586 600054
rect 238822 599818 239004 600054
rect 238404 599734 239004 599818
rect 238404 599498 238586 599734
rect 238822 599498 239004 599734
rect 238404 564054 239004 599498
rect 238404 563818 238586 564054
rect 238822 563818 239004 564054
rect 238404 563734 239004 563818
rect 238404 563498 238586 563734
rect 238822 563498 239004 563734
rect 238404 528054 239004 563498
rect 238404 527818 238586 528054
rect 238822 527818 239004 528054
rect 238404 527734 239004 527818
rect 238404 527498 238586 527734
rect 238822 527498 239004 527734
rect 238404 492054 239004 527498
rect 238404 491818 238586 492054
rect 238822 491818 239004 492054
rect 238404 491734 239004 491818
rect 238404 491498 238586 491734
rect 238822 491498 239004 491734
rect 238404 456054 239004 491498
rect 238404 455818 238586 456054
rect 238822 455818 239004 456054
rect 238404 455734 239004 455818
rect 238404 455498 238586 455734
rect 238822 455498 239004 455734
rect 238404 420054 239004 455498
rect 238404 419818 238586 420054
rect 238822 419818 239004 420054
rect 238404 419734 239004 419818
rect 238404 419498 238586 419734
rect 238822 419498 239004 419734
rect 238404 384054 239004 419498
rect 238404 383818 238586 384054
rect 238822 383818 239004 384054
rect 238404 383734 239004 383818
rect 238404 383498 238586 383734
rect 238822 383498 239004 383734
rect 238404 348054 239004 383498
rect 238404 347818 238586 348054
rect 238822 347818 239004 348054
rect 238404 347734 239004 347818
rect 238404 347498 238586 347734
rect 238822 347498 239004 347734
rect 238404 312054 239004 347498
rect 238404 311818 238586 312054
rect 238822 311818 239004 312054
rect 238404 311734 239004 311818
rect 238404 311498 238586 311734
rect 238822 311498 239004 311734
rect 238404 276054 239004 311498
rect 238404 275818 238586 276054
rect 238822 275818 239004 276054
rect 238404 275734 239004 275818
rect 238404 275498 238586 275734
rect 238822 275498 239004 275734
rect 238404 240054 239004 275498
rect 238404 239818 238586 240054
rect 238822 239818 239004 240054
rect 238404 239734 239004 239818
rect 238404 239498 238586 239734
rect 238822 239498 239004 239734
rect 238404 204054 239004 239498
rect 238404 203818 238586 204054
rect 238822 203818 239004 204054
rect 238404 203734 239004 203818
rect 238404 203498 238586 203734
rect 238822 203498 239004 203734
rect 238404 168054 239004 203498
rect 238404 167818 238586 168054
rect 238822 167818 239004 168054
rect 238404 167734 239004 167818
rect 238404 167498 238586 167734
rect 238822 167498 239004 167734
rect 238404 132054 239004 167498
rect 238404 131818 238586 132054
rect 238822 131818 239004 132054
rect 238404 131734 239004 131818
rect 238404 131498 238586 131734
rect 238822 131498 239004 131734
rect 238404 96054 239004 131498
rect 238404 95818 238586 96054
rect 238822 95818 239004 96054
rect 238404 95734 239004 95818
rect 238404 95498 238586 95734
rect 238822 95498 239004 95734
rect 238404 60054 239004 95498
rect 238404 59818 238586 60054
rect 238822 59818 239004 60054
rect 238404 59734 239004 59818
rect 238404 59498 238586 59734
rect 238822 59498 239004 59734
rect 238404 24054 239004 59498
rect 238404 23818 238586 24054
rect 238822 23818 239004 24054
rect 238404 23734 239004 23818
rect 238404 23498 238586 23734
rect 238822 23498 239004 23734
rect 238404 -3166 239004 23498
rect 238404 -3402 238586 -3166
rect 238822 -3402 239004 -3166
rect 238404 -3486 239004 -3402
rect 238404 -3722 238586 -3486
rect 238822 -3722 239004 -3486
rect 238404 -3744 239004 -3722
rect 242004 675654 242604 708982
rect 242004 675418 242186 675654
rect 242422 675418 242604 675654
rect 242004 675334 242604 675418
rect 242004 675098 242186 675334
rect 242422 675098 242604 675334
rect 242004 639654 242604 675098
rect 242004 639418 242186 639654
rect 242422 639418 242604 639654
rect 242004 639334 242604 639418
rect 242004 639098 242186 639334
rect 242422 639098 242604 639334
rect 242004 603654 242604 639098
rect 242004 603418 242186 603654
rect 242422 603418 242604 603654
rect 242004 603334 242604 603418
rect 242004 603098 242186 603334
rect 242422 603098 242604 603334
rect 242004 567654 242604 603098
rect 242004 567418 242186 567654
rect 242422 567418 242604 567654
rect 242004 567334 242604 567418
rect 242004 567098 242186 567334
rect 242422 567098 242604 567334
rect 242004 531654 242604 567098
rect 242004 531418 242186 531654
rect 242422 531418 242604 531654
rect 242004 531334 242604 531418
rect 242004 531098 242186 531334
rect 242422 531098 242604 531334
rect 242004 495654 242604 531098
rect 242004 495418 242186 495654
rect 242422 495418 242604 495654
rect 242004 495334 242604 495418
rect 242004 495098 242186 495334
rect 242422 495098 242604 495334
rect 242004 459654 242604 495098
rect 242004 459418 242186 459654
rect 242422 459418 242604 459654
rect 242004 459334 242604 459418
rect 242004 459098 242186 459334
rect 242422 459098 242604 459334
rect 242004 423654 242604 459098
rect 242004 423418 242186 423654
rect 242422 423418 242604 423654
rect 242004 423334 242604 423418
rect 242004 423098 242186 423334
rect 242422 423098 242604 423334
rect 242004 387654 242604 423098
rect 242004 387418 242186 387654
rect 242422 387418 242604 387654
rect 242004 387334 242604 387418
rect 242004 387098 242186 387334
rect 242422 387098 242604 387334
rect 242004 351654 242604 387098
rect 242004 351418 242186 351654
rect 242422 351418 242604 351654
rect 242004 351334 242604 351418
rect 242004 351098 242186 351334
rect 242422 351098 242604 351334
rect 242004 315654 242604 351098
rect 242004 315418 242186 315654
rect 242422 315418 242604 315654
rect 242004 315334 242604 315418
rect 242004 315098 242186 315334
rect 242422 315098 242604 315334
rect 242004 279654 242604 315098
rect 242004 279418 242186 279654
rect 242422 279418 242604 279654
rect 242004 279334 242604 279418
rect 242004 279098 242186 279334
rect 242422 279098 242604 279334
rect 242004 243654 242604 279098
rect 242004 243418 242186 243654
rect 242422 243418 242604 243654
rect 242004 243334 242604 243418
rect 242004 243098 242186 243334
rect 242422 243098 242604 243334
rect 242004 207654 242604 243098
rect 242004 207418 242186 207654
rect 242422 207418 242604 207654
rect 242004 207334 242604 207418
rect 242004 207098 242186 207334
rect 242422 207098 242604 207334
rect 242004 171654 242604 207098
rect 242004 171418 242186 171654
rect 242422 171418 242604 171654
rect 242004 171334 242604 171418
rect 242004 171098 242186 171334
rect 242422 171098 242604 171334
rect 242004 135654 242604 171098
rect 242004 135418 242186 135654
rect 242422 135418 242604 135654
rect 242004 135334 242604 135418
rect 242004 135098 242186 135334
rect 242422 135098 242604 135334
rect 242004 99654 242604 135098
rect 242004 99418 242186 99654
rect 242422 99418 242604 99654
rect 242004 99334 242604 99418
rect 242004 99098 242186 99334
rect 242422 99098 242604 99334
rect 242004 63654 242604 99098
rect 242004 63418 242186 63654
rect 242422 63418 242604 63654
rect 242004 63334 242604 63418
rect 242004 63098 242186 63334
rect 242422 63098 242604 63334
rect 242004 27654 242604 63098
rect 242004 27418 242186 27654
rect 242422 27418 242604 27654
rect 242004 27334 242604 27418
rect 242004 27098 242186 27334
rect 242422 27098 242604 27334
rect 242004 -5046 242604 27098
rect 242004 -5282 242186 -5046
rect 242422 -5282 242604 -5046
rect 242004 -5366 242604 -5282
rect 242004 -5602 242186 -5366
rect 242422 -5602 242604 -5366
rect 242004 -5624 242604 -5602
rect 245604 679254 246204 710862
rect 263604 710478 264204 711440
rect 263604 710242 263786 710478
rect 264022 710242 264204 710478
rect 263604 710158 264204 710242
rect 263604 709922 263786 710158
rect 264022 709922 264204 710158
rect 260004 708598 260604 709560
rect 260004 708362 260186 708598
rect 260422 708362 260604 708598
rect 260004 708278 260604 708362
rect 260004 708042 260186 708278
rect 260422 708042 260604 708278
rect 256404 706718 257004 707680
rect 256404 706482 256586 706718
rect 256822 706482 257004 706718
rect 256404 706398 257004 706482
rect 256404 706162 256586 706398
rect 256822 706162 257004 706398
rect 245604 679018 245786 679254
rect 246022 679018 246204 679254
rect 245604 678934 246204 679018
rect 245604 678698 245786 678934
rect 246022 678698 246204 678934
rect 245604 643254 246204 678698
rect 245604 643018 245786 643254
rect 246022 643018 246204 643254
rect 245604 642934 246204 643018
rect 245604 642698 245786 642934
rect 246022 642698 246204 642934
rect 245604 607254 246204 642698
rect 245604 607018 245786 607254
rect 246022 607018 246204 607254
rect 245604 606934 246204 607018
rect 245604 606698 245786 606934
rect 246022 606698 246204 606934
rect 245604 571254 246204 606698
rect 245604 571018 245786 571254
rect 246022 571018 246204 571254
rect 245604 570934 246204 571018
rect 245604 570698 245786 570934
rect 246022 570698 246204 570934
rect 245604 535254 246204 570698
rect 245604 535018 245786 535254
rect 246022 535018 246204 535254
rect 245604 534934 246204 535018
rect 245604 534698 245786 534934
rect 246022 534698 246204 534934
rect 245604 499254 246204 534698
rect 245604 499018 245786 499254
rect 246022 499018 246204 499254
rect 245604 498934 246204 499018
rect 245604 498698 245786 498934
rect 246022 498698 246204 498934
rect 245604 463254 246204 498698
rect 245604 463018 245786 463254
rect 246022 463018 246204 463254
rect 245604 462934 246204 463018
rect 245604 462698 245786 462934
rect 246022 462698 246204 462934
rect 245604 427254 246204 462698
rect 245604 427018 245786 427254
rect 246022 427018 246204 427254
rect 245604 426934 246204 427018
rect 245604 426698 245786 426934
rect 246022 426698 246204 426934
rect 245604 391254 246204 426698
rect 245604 391018 245786 391254
rect 246022 391018 246204 391254
rect 245604 390934 246204 391018
rect 245604 390698 245786 390934
rect 246022 390698 246204 390934
rect 245604 355254 246204 390698
rect 245604 355018 245786 355254
rect 246022 355018 246204 355254
rect 245604 354934 246204 355018
rect 245604 354698 245786 354934
rect 246022 354698 246204 354934
rect 245604 319254 246204 354698
rect 245604 319018 245786 319254
rect 246022 319018 246204 319254
rect 245604 318934 246204 319018
rect 245604 318698 245786 318934
rect 246022 318698 246204 318934
rect 245604 283254 246204 318698
rect 245604 283018 245786 283254
rect 246022 283018 246204 283254
rect 245604 282934 246204 283018
rect 245604 282698 245786 282934
rect 246022 282698 246204 282934
rect 245604 247254 246204 282698
rect 245604 247018 245786 247254
rect 246022 247018 246204 247254
rect 245604 246934 246204 247018
rect 245604 246698 245786 246934
rect 246022 246698 246204 246934
rect 245604 211254 246204 246698
rect 245604 211018 245786 211254
rect 246022 211018 246204 211254
rect 245604 210934 246204 211018
rect 245604 210698 245786 210934
rect 246022 210698 246204 210934
rect 245604 175254 246204 210698
rect 245604 175018 245786 175254
rect 246022 175018 246204 175254
rect 245604 174934 246204 175018
rect 245604 174698 245786 174934
rect 246022 174698 246204 174934
rect 245604 139254 246204 174698
rect 245604 139018 245786 139254
rect 246022 139018 246204 139254
rect 245604 138934 246204 139018
rect 245604 138698 245786 138934
rect 246022 138698 246204 138934
rect 245604 103254 246204 138698
rect 245604 103018 245786 103254
rect 246022 103018 246204 103254
rect 245604 102934 246204 103018
rect 245604 102698 245786 102934
rect 246022 102698 246204 102934
rect 245604 67254 246204 102698
rect 245604 67018 245786 67254
rect 246022 67018 246204 67254
rect 245604 66934 246204 67018
rect 245604 66698 245786 66934
rect 246022 66698 246204 66934
rect 245604 31254 246204 66698
rect 245604 31018 245786 31254
rect 246022 31018 246204 31254
rect 245604 30934 246204 31018
rect 245604 30698 245786 30934
rect 246022 30698 246204 30934
rect 227604 -6222 227786 -5986
rect 228022 -6222 228204 -5986
rect 227604 -6306 228204 -6222
rect 227604 -6542 227786 -6306
rect 228022 -6542 228204 -6306
rect 227604 -7504 228204 -6542
rect 245604 -6926 246204 30698
rect 252804 704838 253404 705800
rect 252804 704602 252986 704838
rect 253222 704602 253404 704838
rect 252804 704518 253404 704602
rect 252804 704282 252986 704518
rect 253222 704282 253404 704518
rect 252804 686454 253404 704282
rect 252804 686218 252986 686454
rect 253222 686218 253404 686454
rect 252804 686134 253404 686218
rect 252804 685898 252986 686134
rect 253222 685898 253404 686134
rect 252804 650454 253404 685898
rect 252804 650218 252986 650454
rect 253222 650218 253404 650454
rect 252804 650134 253404 650218
rect 252804 649898 252986 650134
rect 253222 649898 253404 650134
rect 252804 614454 253404 649898
rect 252804 614218 252986 614454
rect 253222 614218 253404 614454
rect 252804 614134 253404 614218
rect 252804 613898 252986 614134
rect 253222 613898 253404 614134
rect 252804 578454 253404 613898
rect 252804 578218 252986 578454
rect 253222 578218 253404 578454
rect 252804 578134 253404 578218
rect 252804 577898 252986 578134
rect 253222 577898 253404 578134
rect 252804 542454 253404 577898
rect 252804 542218 252986 542454
rect 253222 542218 253404 542454
rect 252804 542134 253404 542218
rect 252804 541898 252986 542134
rect 253222 541898 253404 542134
rect 252804 506454 253404 541898
rect 252804 506218 252986 506454
rect 253222 506218 253404 506454
rect 252804 506134 253404 506218
rect 252804 505898 252986 506134
rect 253222 505898 253404 506134
rect 252804 470454 253404 505898
rect 252804 470218 252986 470454
rect 253222 470218 253404 470454
rect 252804 470134 253404 470218
rect 252804 469898 252986 470134
rect 253222 469898 253404 470134
rect 252804 434454 253404 469898
rect 252804 434218 252986 434454
rect 253222 434218 253404 434454
rect 252804 434134 253404 434218
rect 252804 433898 252986 434134
rect 253222 433898 253404 434134
rect 252804 398454 253404 433898
rect 252804 398218 252986 398454
rect 253222 398218 253404 398454
rect 252804 398134 253404 398218
rect 252804 397898 252986 398134
rect 253222 397898 253404 398134
rect 252804 362454 253404 397898
rect 252804 362218 252986 362454
rect 253222 362218 253404 362454
rect 252804 362134 253404 362218
rect 252804 361898 252986 362134
rect 253222 361898 253404 362134
rect 252804 326454 253404 361898
rect 252804 326218 252986 326454
rect 253222 326218 253404 326454
rect 252804 326134 253404 326218
rect 252804 325898 252986 326134
rect 253222 325898 253404 326134
rect 252804 290454 253404 325898
rect 252804 290218 252986 290454
rect 253222 290218 253404 290454
rect 252804 290134 253404 290218
rect 252804 289898 252986 290134
rect 253222 289898 253404 290134
rect 252804 254454 253404 289898
rect 252804 254218 252986 254454
rect 253222 254218 253404 254454
rect 252804 254134 253404 254218
rect 252804 253898 252986 254134
rect 253222 253898 253404 254134
rect 252804 218454 253404 253898
rect 252804 218218 252986 218454
rect 253222 218218 253404 218454
rect 252804 218134 253404 218218
rect 252804 217898 252986 218134
rect 253222 217898 253404 218134
rect 252804 182454 253404 217898
rect 252804 182218 252986 182454
rect 253222 182218 253404 182454
rect 252804 182134 253404 182218
rect 252804 181898 252986 182134
rect 253222 181898 253404 182134
rect 252804 146454 253404 181898
rect 252804 146218 252986 146454
rect 253222 146218 253404 146454
rect 252804 146134 253404 146218
rect 252804 145898 252986 146134
rect 253222 145898 253404 146134
rect 252804 110454 253404 145898
rect 252804 110218 252986 110454
rect 253222 110218 253404 110454
rect 252804 110134 253404 110218
rect 252804 109898 252986 110134
rect 253222 109898 253404 110134
rect 252804 74454 253404 109898
rect 252804 74218 252986 74454
rect 253222 74218 253404 74454
rect 252804 74134 253404 74218
rect 252804 73898 252986 74134
rect 253222 73898 253404 74134
rect 252804 38454 253404 73898
rect 252804 38218 252986 38454
rect 253222 38218 253404 38454
rect 252804 38134 253404 38218
rect 252804 37898 252986 38134
rect 253222 37898 253404 38134
rect 252804 2454 253404 37898
rect 252804 2218 252986 2454
rect 253222 2218 253404 2454
rect 252804 2134 253404 2218
rect 252804 1898 252986 2134
rect 253222 1898 253404 2134
rect 252804 -346 253404 1898
rect 252804 -582 252986 -346
rect 253222 -582 253404 -346
rect 252804 -666 253404 -582
rect 252804 -902 252986 -666
rect 253222 -902 253404 -666
rect 252804 -1864 253404 -902
rect 256404 690054 257004 706162
rect 256404 689818 256586 690054
rect 256822 689818 257004 690054
rect 256404 689734 257004 689818
rect 256404 689498 256586 689734
rect 256822 689498 257004 689734
rect 256404 654054 257004 689498
rect 256404 653818 256586 654054
rect 256822 653818 257004 654054
rect 256404 653734 257004 653818
rect 256404 653498 256586 653734
rect 256822 653498 257004 653734
rect 256404 618054 257004 653498
rect 256404 617818 256586 618054
rect 256822 617818 257004 618054
rect 256404 617734 257004 617818
rect 256404 617498 256586 617734
rect 256822 617498 257004 617734
rect 256404 582054 257004 617498
rect 256404 581818 256586 582054
rect 256822 581818 257004 582054
rect 256404 581734 257004 581818
rect 256404 581498 256586 581734
rect 256822 581498 257004 581734
rect 256404 546054 257004 581498
rect 256404 545818 256586 546054
rect 256822 545818 257004 546054
rect 256404 545734 257004 545818
rect 256404 545498 256586 545734
rect 256822 545498 257004 545734
rect 256404 510054 257004 545498
rect 256404 509818 256586 510054
rect 256822 509818 257004 510054
rect 256404 509734 257004 509818
rect 256404 509498 256586 509734
rect 256822 509498 257004 509734
rect 256404 474054 257004 509498
rect 256404 473818 256586 474054
rect 256822 473818 257004 474054
rect 256404 473734 257004 473818
rect 256404 473498 256586 473734
rect 256822 473498 257004 473734
rect 256404 438054 257004 473498
rect 256404 437818 256586 438054
rect 256822 437818 257004 438054
rect 256404 437734 257004 437818
rect 256404 437498 256586 437734
rect 256822 437498 257004 437734
rect 256404 402054 257004 437498
rect 256404 401818 256586 402054
rect 256822 401818 257004 402054
rect 256404 401734 257004 401818
rect 256404 401498 256586 401734
rect 256822 401498 257004 401734
rect 256404 366054 257004 401498
rect 256404 365818 256586 366054
rect 256822 365818 257004 366054
rect 256404 365734 257004 365818
rect 256404 365498 256586 365734
rect 256822 365498 257004 365734
rect 256404 330054 257004 365498
rect 256404 329818 256586 330054
rect 256822 329818 257004 330054
rect 256404 329734 257004 329818
rect 256404 329498 256586 329734
rect 256822 329498 257004 329734
rect 256404 294054 257004 329498
rect 260004 693654 260604 708042
rect 260004 693418 260186 693654
rect 260422 693418 260604 693654
rect 260004 693334 260604 693418
rect 260004 693098 260186 693334
rect 260422 693098 260604 693334
rect 260004 657654 260604 693098
rect 260004 657418 260186 657654
rect 260422 657418 260604 657654
rect 260004 657334 260604 657418
rect 260004 657098 260186 657334
rect 260422 657098 260604 657334
rect 260004 621654 260604 657098
rect 260004 621418 260186 621654
rect 260422 621418 260604 621654
rect 260004 621334 260604 621418
rect 260004 621098 260186 621334
rect 260422 621098 260604 621334
rect 260004 585654 260604 621098
rect 260004 585418 260186 585654
rect 260422 585418 260604 585654
rect 260004 585334 260604 585418
rect 260004 585098 260186 585334
rect 260422 585098 260604 585334
rect 260004 549654 260604 585098
rect 260004 549418 260186 549654
rect 260422 549418 260604 549654
rect 260004 549334 260604 549418
rect 260004 549098 260186 549334
rect 260422 549098 260604 549334
rect 260004 513654 260604 549098
rect 260004 513418 260186 513654
rect 260422 513418 260604 513654
rect 260004 513334 260604 513418
rect 260004 513098 260186 513334
rect 260422 513098 260604 513334
rect 260004 477654 260604 513098
rect 260004 477418 260186 477654
rect 260422 477418 260604 477654
rect 260004 477334 260604 477418
rect 260004 477098 260186 477334
rect 260422 477098 260604 477334
rect 260004 441654 260604 477098
rect 260004 441418 260186 441654
rect 260422 441418 260604 441654
rect 260004 441334 260604 441418
rect 260004 441098 260186 441334
rect 260422 441098 260604 441334
rect 260004 405654 260604 441098
rect 260004 405418 260186 405654
rect 260422 405418 260604 405654
rect 260004 405334 260604 405418
rect 260004 405098 260186 405334
rect 260422 405098 260604 405334
rect 260004 369654 260604 405098
rect 260004 369418 260186 369654
rect 260422 369418 260604 369654
rect 260004 369334 260604 369418
rect 260004 369098 260186 369334
rect 260422 369098 260604 369334
rect 260004 333654 260604 369098
rect 260004 333418 260186 333654
rect 260422 333418 260604 333654
rect 260004 333334 260604 333418
rect 260004 333098 260186 333334
rect 260422 333098 260604 333334
rect 257659 317388 257725 317389
rect 257659 317324 257660 317388
rect 257724 317324 257725 317388
rect 257659 317323 257725 317324
rect 257662 311813 257722 317323
rect 257659 311812 257725 311813
rect 257659 311748 257660 311812
rect 257724 311748 257725 311812
rect 257659 311747 257725 311748
rect 256404 293818 256586 294054
rect 256822 293818 257004 294054
rect 256404 293734 257004 293818
rect 256404 293498 256586 293734
rect 256822 293498 257004 293734
rect 256404 258054 257004 293498
rect 256404 257818 256586 258054
rect 256822 257818 257004 258054
rect 256404 257734 257004 257818
rect 256404 257498 256586 257734
rect 256822 257498 257004 257734
rect 256404 222054 257004 257498
rect 256404 221818 256586 222054
rect 256822 221818 257004 222054
rect 256404 221734 257004 221818
rect 256404 221498 256586 221734
rect 256822 221498 257004 221734
rect 256404 186054 257004 221498
rect 256404 185818 256586 186054
rect 256822 185818 257004 186054
rect 256404 185734 257004 185818
rect 256404 185498 256586 185734
rect 256822 185498 257004 185734
rect 256404 150054 257004 185498
rect 256404 149818 256586 150054
rect 256822 149818 257004 150054
rect 256404 149734 257004 149818
rect 256404 149498 256586 149734
rect 256822 149498 257004 149734
rect 256404 114054 257004 149498
rect 256404 113818 256586 114054
rect 256822 113818 257004 114054
rect 256404 113734 257004 113818
rect 256404 113498 256586 113734
rect 256822 113498 257004 113734
rect 256404 78054 257004 113498
rect 256404 77818 256586 78054
rect 256822 77818 257004 78054
rect 256404 77734 257004 77818
rect 256404 77498 256586 77734
rect 256822 77498 257004 77734
rect 256404 42054 257004 77498
rect 256404 41818 256586 42054
rect 256822 41818 257004 42054
rect 256404 41734 257004 41818
rect 256404 41498 256586 41734
rect 256822 41498 257004 41734
rect 256404 6054 257004 41498
rect 256404 5818 256586 6054
rect 256822 5818 257004 6054
rect 256404 5734 257004 5818
rect 256404 5498 256586 5734
rect 256822 5498 257004 5734
rect 256404 -2226 257004 5498
rect 256404 -2462 256586 -2226
rect 256822 -2462 257004 -2226
rect 256404 -2546 257004 -2462
rect 256404 -2782 256586 -2546
rect 256822 -2782 257004 -2546
rect 256404 -3744 257004 -2782
rect 260004 297654 260604 333098
rect 260004 297418 260186 297654
rect 260422 297418 260604 297654
rect 260004 297334 260604 297418
rect 260004 297098 260186 297334
rect 260422 297098 260604 297334
rect 260004 261654 260604 297098
rect 260004 261418 260186 261654
rect 260422 261418 260604 261654
rect 260004 261334 260604 261418
rect 260004 261098 260186 261334
rect 260422 261098 260604 261334
rect 260004 225654 260604 261098
rect 260004 225418 260186 225654
rect 260422 225418 260604 225654
rect 260004 225334 260604 225418
rect 260004 225098 260186 225334
rect 260422 225098 260604 225334
rect 260004 189654 260604 225098
rect 260004 189418 260186 189654
rect 260422 189418 260604 189654
rect 260004 189334 260604 189418
rect 260004 189098 260186 189334
rect 260422 189098 260604 189334
rect 260004 153654 260604 189098
rect 260004 153418 260186 153654
rect 260422 153418 260604 153654
rect 260004 153334 260604 153418
rect 260004 153098 260186 153334
rect 260422 153098 260604 153334
rect 260004 117654 260604 153098
rect 260004 117418 260186 117654
rect 260422 117418 260604 117654
rect 260004 117334 260604 117418
rect 260004 117098 260186 117334
rect 260422 117098 260604 117334
rect 260004 81654 260604 117098
rect 260004 81418 260186 81654
rect 260422 81418 260604 81654
rect 260004 81334 260604 81418
rect 260004 81098 260186 81334
rect 260422 81098 260604 81334
rect 260004 45654 260604 81098
rect 260004 45418 260186 45654
rect 260422 45418 260604 45654
rect 260004 45334 260604 45418
rect 260004 45098 260186 45334
rect 260422 45098 260604 45334
rect 260004 9654 260604 45098
rect 260004 9418 260186 9654
rect 260422 9418 260604 9654
rect 260004 9334 260604 9418
rect 260004 9098 260186 9334
rect 260422 9098 260604 9334
rect 260004 -4106 260604 9098
rect 260004 -4342 260186 -4106
rect 260422 -4342 260604 -4106
rect 260004 -4426 260604 -4342
rect 260004 -4662 260186 -4426
rect 260422 -4662 260604 -4426
rect 260004 -5624 260604 -4662
rect 263604 697254 264204 709922
rect 281604 711418 282204 711440
rect 281604 711182 281786 711418
rect 282022 711182 282204 711418
rect 281604 711098 282204 711182
rect 281604 710862 281786 711098
rect 282022 710862 282204 711098
rect 278004 709538 278604 709560
rect 278004 709302 278186 709538
rect 278422 709302 278604 709538
rect 278004 709218 278604 709302
rect 278004 708982 278186 709218
rect 278422 708982 278604 709218
rect 274404 707658 275004 707680
rect 274404 707422 274586 707658
rect 274822 707422 275004 707658
rect 274404 707338 275004 707422
rect 274404 707102 274586 707338
rect 274822 707102 275004 707338
rect 263604 697018 263786 697254
rect 264022 697018 264204 697254
rect 263604 696934 264204 697018
rect 263604 696698 263786 696934
rect 264022 696698 264204 696934
rect 263604 661254 264204 696698
rect 263604 661018 263786 661254
rect 264022 661018 264204 661254
rect 263604 660934 264204 661018
rect 263604 660698 263786 660934
rect 264022 660698 264204 660934
rect 263604 625254 264204 660698
rect 263604 625018 263786 625254
rect 264022 625018 264204 625254
rect 263604 624934 264204 625018
rect 263604 624698 263786 624934
rect 264022 624698 264204 624934
rect 263604 589254 264204 624698
rect 263604 589018 263786 589254
rect 264022 589018 264204 589254
rect 263604 588934 264204 589018
rect 263604 588698 263786 588934
rect 264022 588698 264204 588934
rect 263604 553254 264204 588698
rect 263604 553018 263786 553254
rect 264022 553018 264204 553254
rect 263604 552934 264204 553018
rect 263604 552698 263786 552934
rect 264022 552698 264204 552934
rect 263604 517254 264204 552698
rect 263604 517018 263786 517254
rect 264022 517018 264204 517254
rect 263604 516934 264204 517018
rect 263604 516698 263786 516934
rect 264022 516698 264204 516934
rect 263604 481254 264204 516698
rect 263604 481018 263786 481254
rect 264022 481018 264204 481254
rect 263604 480934 264204 481018
rect 263604 480698 263786 480934
rect 264022 480698 264204 480934
rect 263604 445254 264204 480698
rect 263604 445018 263786 445254
rect 264022 445018 264204 445254
rect 263604 444934 264204 445018
rect 263604 444698 263786 444934
rect 264022 444698 264204 444934
rect 263604 409254 264204 444698
rect 270804 705778 271404 705800
rect 270804 705542 270986 705778
rect 271222 705542 271404 705778
rect 270804 705458 271404 705542
rect 270804 705222 270986 705458
rect 271222 705222 271404 705458
rect 270804 668454 271404 705222
rect 270804 668218 270986 668454
rect 271222 668218 271404 668454
rect 270804 668134 271404 668218
rect 270804 667898 270986 668134
rect 271222 667898 271404 668134
rect 270804 632454 271404 667898
rect 270804 632218 270986 632454
rect 271222 632218 271404 632454
rect 270804 632134 271404 632218
rect 270804 631898 270986 632134
rect 271222 631898 271404 632134
rect 270804 596454 271404 631898
rect 270804 596218 270986 596454
rect 271222 596218 271404 596454
rect 270804 596134 271404 596218
rect 270804 595898 270986 596134
rect 271222 595898 271404 596134
rect 270804 560454 271404 595898
rect 270804 560218 270986 560454
rect 271222 560218 271404 560454
rect 270804 560134 271404 560218
rect 270804 559898 270986 560134
rect 271222 559898 271404 560134
rect 270804 524454 271404 559898
rect 270804 524218 270986 524454
rect 271222 524218 271404 524454
rect 270804 524134 271404 524218
rect 270804 523898 270986 524134
rect 271222 523898 271404 524134
rect 270804 488454 271404 523898
rect 270804 488218 270986 488454
rect 271222 488218 271404 488454
rect 270804 488134 271404 488218
rect 270804 487898 270986 488134
rect 271222 487898 271404 488134
rect 270804 452454 271404 487898
rect 270804 452218 270986 452454
rect 271222 452218 271404 452454
rect 270804 452134 271404 452218
rect 270804 451898 270986 452134
rect 271222 451898 271404 452134
rect 270804 416454 271404 451898
rect 270804 416218 270986 416454
rect 271222 416218 271404 416454
rect 270804 416134 271404 416218
rect 270804 415898 270986 416134
rect 271222 415898 271404 416134
rect 266859 410412 266925 410413
rect 266859 410348 266860 410412
rect 266924 410348 266925 410412
rect 266859 410347 266925 410348
rect 263604 409018 263786 409254
rect 264022 409018 264204 409254
rect 263604 408934 264204 409018
rect 263604 408698 263786 408934
rect 264022 408698 264204 408934
rect 263604 373254 264204 408698
rect 263604 373018 263786 373254
rect 264022 373018 264204 373254
rect 263604 372934 264204 373018
rect 263604 372698 263786 372934
rect 264022 372698 264204 372934
rect 263604 337254 264204 372698
rect 263604 337018 263786 337254
rect 264022 337018 264204 337254
rect 263604 336934 264204 337018
rect 263604 336698 263786 336934
rect 264022 336698 264204 336934
rect 263604 301254 264204 336698
rect 263604 301018 263786 301254
rect 264022 301018 264204 301254
rect 263604 300934 264204 301018
rect 263604 300698 263786 300934
rect 264022 300698 264204 300934
rect 263604 265254 264204 300698
rect 263604 265018 263786 265254
rect 264022 265018 264204 265254
rect 263604 264934 264204 265018
rect 263604 264698 263786 264934
rect 264022 264698 264204 264934
rect 263604 229254 264204 264698
rect 263604 229018 263786 229254
rect 264022 229018 264204 229254
rect 263604 228934 264204 229018
rect 263604 228698 263786 228934
rect 264022 228698 264204 228934
rect 263604 193254 264204 228698
rect 266862 202877 266922 410347
rect 267779 410276 267845 410277
rect 267779 410212 267780 410276
rect 267844 410212 267845 410276
rect 267779 410211 267845 410212
rect 266859 202876 266925 202877
rect 266859 202812 266860 202876
rect 266924 202812 266925 202876
rect 266859 202811 266925 202812
rect 267782 202197 267842 410211
rect 267963 410140 268029 410141
rect 267963 410076 267964 410140
rect 268028 410076 268029 410140
rect 267963 410075 268029 410076
rect 267779 202196 267845 202197
rect 267779 202132 267780 202196
rect 267844 202132 267845 202196
rect 267779 202131 267845 202132
rect 267966 201653 268026 410075
rect 268147 410004 268213 410005
rect 268147 409940 268148 410004
rect 268212 409940 268213 410004
rect 268147 409939 268213 409940
rect 268150 338741 268210 409939
rect 270804 380454 271404 415898
rect 270804 380218 270986 380454
rect 271222 380218 271404 380454
rect 270804 380134 271404 380218
rect 270804 379898 270986 380134
rect 271222 379898 271404 380134
rect 270804 344454 271404 379898
rect 270804 344218 270986 344454
rect 271222 344218 271404 344454
rect 270804 344134 271404 344218
rect 270804 343898 270986 344134
rect 271222 343898 271404 344134
rect 268147 338740 268213 338741
rect 268147 338676 268148 338740
rect 268212 338676 268213 338740
rect 268147 338675 268213 338676
rect 270804 308454 271404 343898
rect 270804 308218 270986 308454
rect 271222 308218 271404 308454
rect 270804 308134 271404 308218
rect 270804 307898 270986 308134
rect 271222 307898 271404 308134
rect 270804 272454 271404 307898
rect 270804 272218 270986 272454
rect 271222 272218 271404 272454
rect 270804 272134 271404 272218
rect 270804 271898 270986 272134
rect 271222 271898 271404 272134
rect 270804 236454 271404 271898
rect 270804 236218 270986 236454
rect 271222 236218 271404 236454
rect 270804 236134 271404 236218
rect 270804 235898 270986 236134
rect 271222 235898 271404 236134
rect 267963 201652 268029 201653
rect 267963 201588 267964 201652
rect 268028 201588 268029 201652
rect 267963 201587 268029 201588
rect 263604 193018 263786 193254
rect 264022 193018 264204 193254
rect 263604 192934 264204 193018
rect 263604 192698 263786 192934
rect 264022 192698 264204 192934
rect 263604 157254 264204 192698
rect 263604 157018 263786 157254
rect 264022 157018 264204 157254
rect 263604 156934 264204 157018
rect 263604 156698 263786 156934
rect 264022 156698 264204 156934
rect 263604 121254 264204 156698
rect 263604 121018 263786 121254
rect 264022 121018 264204 121254
rect 263604 120934 264204 121018
rect 263604 120698 263786 120934
rect 264022 120698 264204 120934
rect 263604 85254 264204 120698
rect 263604 85018 263786 85254
rect 264022 85018 264204 85254
rect 263604 84934 264204 85018
rect 263604 84698 263786 84934
rect 264022 84698 264204 84934
rect 263604 49254 264204 84698
rect 263604 49018 263786 49254
rect 264022 49018 264204 49254
rect 263604 48934 264204 49018
rect 263604 48698 263786 48934
rect 264022 48698 264204 48934
rect 263604 13254 264204 48698
rect 263604 13018 263786 13254
rect 264022 13018 264204 13254
rect 263604 12934 264204 13018
rect 263604 12698 263786 12934
rect 264022 12698 264204 12934
rect 245604 -7162 245786 -6926
rect 246022 -7162 246204 -6926
rect 245604 -7246 246204 -7162
rect 245604 -7482 245786 -7246
rect 246022 -7482 246204 -7246
rect 245604 -7504 246204 -7482
rect 263604 -5986 264204 12698
rect 270804 200454 271404 235898
rect 270804 200218 270986 200454
rect 271222 200218 271404 200454
rect 270804 200134 271404 200218
rect 270804 199898 270986 200134
rect 271222 199898 271404 200134
rect 270804 164454 271404 199898
rect 270804 164218 270986 164454
rect 271222 164218 271404 164454
rect 270804 164134 271404 164218
rect 270804 163898 270986 164134
rect 271222 163898 271404 164134
rect 270804 128454 271404 163898
rect 270804 128218 270986 128454
rect 271222 128218 271404 128454
rect 270804 128134 271404 128218
rect 270804 127898 270986 128134
rect 271222 127898 271404 128134
rect 270804 92454 271404 127898
rect 270804 92218 270986 92454
rect 271222 92218 271404 92454
rect 270804 92134 271404 92218
rect 270804 91898 270986 92134
rect 271222 91898 271404 92134
rect 270804 56454 271404 91898
rect 270804 56218 270986 56454
rect 271222 56218 271404 56454
rect 270804 56134 271404 56218
rect 270804 55898 270986 56134
rect 271222 55898 271404 56134
rect 270804 20454 271404 55898
rect 270804 20218 270986 20454
rect 271222 20218 271404 20454
rect 270804 20134 271404 20218
rect 270804 19898 270986 20134
rect 271222 19898 271404 20134
rect 270804 -1286 271404 19898
rect 270804 -1522 270986 -1286
rect 271222 -1522 271404 -1286
rect 270804 -1606 271404 -1522
rect 270804 -1842 270986 -1606
rect 271222 -1842 271404 -1606
rect 270804 -1864 271404 -1842
rect 274404 672054 275004 707102
rect 274404 671818 274586 672054
rect 274822 671818 275004 672054
rect 274404 671734 275004 671818
rect 274404 671498 274586 671734
rect 274822 671498 275004 671734
rect 274404 636054 275004 671498
rect 274404 635818 274586 636054
rect 274822 635818 275004 636054
rect 274404 635734 275004 635818
rect 274404 635498 274586 635734
rect 274822 635498 275004 635734
rect 274404 600054 275004 635498
rect 274404 599818 274586 600054
rect 274822 599818 275004 600054
rect 274404 599734 275004 599818
rect 274404 599498 274586 599734
rect 274822 599498 275004 599734
rect 274404 564054 275004 599498
rect 274404 563818 274586 564054
rect 274822 563818 275004 564054
rect 274404 563734 275004 563818
rect 274404 563498 274586 563734
rect 274822 563498 275004 563734
rect 274404 528054 275004 563498
rect 274404 527818 274586 528054
rect 274822 527818 275004 528054
rect 274404 527734 275004 527818
rect 274404 527498 274586 527734
rect 274822 527498 275004 527734
rect 274404 492054 275004 527498
rect 274404 491818 274586 492054
rect 274822 491818 275004 492054
rect 274404 491734 275004 491818
rect 274404 491498 274586 491734
rect 274822 491498 275004 491734
rect 274404 456054 275004 491498
rect 274404 455818 274586 456054
rect 274822 455818 275004 456054
rect 274404 455734 275004 455818
rect 274404 455498 274586 455734
rect 274822 455498 275004 455734
rect 274404 420054 275004 455498
rect 274404 419818 274586 420054
rect 274822 419818 275004 420054
rect 274404 419734 275004 419818
rect 274404 419498 274586 419734
rect 274822 419498 275004 419734
rect 274404 384054 275004 419498
rect 274404 383818 274586 384054
rect 274822 383818 275004 384054
rect 274404 383734 275004 383818
rect 274404 383498 274586 383734
rect 274822 383498 275004 383734
rect 274404 348054 275004 383498
rect 274404 347818 274586 348054
rect 274822 347818 275004 348054
rect 274404 347734 275004 347818
rect 274404 347498 274586 347734
rect 274822 347498 275004 347734
rect 274404 312054 275004 347498
rect 274404 311818 274586 312054
rect 274822 311818 275004 312054
rect 274404 311734 275004 311818
rect 274404 311498 274586 311734
rect 274822 311498 275004 311734
rect 274404 276054 275004 311498
rect 274404 275818 274586 276054
rect 274822 275818 275004 276054
rect 274404 275734 275004 275818
rect 274404 275498 274586 275734
rect 274822 275498 275004 275734
rect 274404 240054 275004 275498
rect 274404 239818 274586 240054
rect 274822 239818 275004 240054
rect 274404 239734 275004 239818
rect 274404 239498 274586 239734
rect 274822 239498 275004 239734
rect 274404 204054 275004 239498
rect 274404 203818 274586 204054
rect 274822 203818 275004 204054
rect 274404 203734 275004 203818
rect 274404 203498 274586 203734
rect 274822 203498 275004 203734
rect 274404 168054 275004 203498
rect 274404 167818 274586 168054
rect 274822 167818 275004 168054
rect 274404 167734 275004 167818
rect 274404 167498 274586 167734
rect 274822 167498 275004 167734
rect 274404 132054 275004 167498
rect 274404 131818 274586 132054
rect 274822 131818 275004 132054
rect 274404 131734 275004 131818
rect 274404 131498 274586 131734
rect 274822 131498 275004 131734
rect 274404 96054 275004 131498
rect 274404 95818 274586 96054
rect 274822 95818 275004 96054
rect 274404 95734 275004 95818
rect 274404 95498 274586 95734
rect 274822 95498 275004 95734
rect 274404 60054 275004 95498
rect 274404 59818 274586 60054
rect 274822 59818 275004 60054
rect 274404 59734 275004 59818
rect 274404 59498 274586 59734
rect 274822 59498 275004 59734
rect 274404 24054 275004 59498
rect 274404 23818 274586 24054
rect 274822 23818 275004 24054
rect 274404 23734 275004 23818
rect 274404 23498 274586 23734
rect 274822 23498 275004 23734
rect 274404 -3166 275004 23498
rect 274404 -3402 274586 -3166
rect 274822 -3402 275004 -3166
rect 274404 -3486 275004 -3402
rect 274404 -3722 274586 -3486
rect 274822 -3722 275004 -3486
rect 274404 -3744 275004 -3722
rect 278004 675654 278604 708982
rect 278004 675418 278186 675654
rect 278422 675418 278604 675654
rect 278004 675334 278604 675418
rect 278004 675098 278186 675334
rect 278422 675098 278604 675334
rect 278004 639654 278604 675098
rect 278004 639418 278186 639654
rect 278422 639418 278604 639654
rect 278004 639334 278604 639418
rect 278004 639098 278186 639334
rect 278422 639098 278604 639334
rect 278004 603654 278604 639098
rect 278004 603418 278186 603654
rect 278422 603418 278604 603654
rect 278004 603334 278604 603418
rect 278004 603098 278186 603334
rect 278422 603098 278604 603334
rect 278004 567654 278604 603098
rect 278004 567418 278186 567654
rect 278422 567418 278604 567654
rect 278004 567334 278604 567418
rect 278004 567098 278186 567334
rect 278422 567098 278604 567334
rect 278004 531654 278604 567098
rect 278004 531418 278186 531654
rect 278422 531418 278604 531654
rect 278004 531334 278604 531418
rect 278004 531098 278186 531334
rect 278422 531098 278604 531334
rect 278004 495654 278604 531098
rect 278004 495418 278186 495654
rect 278422 495418 278604 495654
rect 278004 495334 278604 495418
rect 278004 495098 278186 495334
rect 278422 495098 278604 495334
rect 278004 459654 278604 495098
rect 278004 459418 278186 459654
rect 278422 459418 278604 459654
rect 278004 459334 278604 459418
rect 278004 459098 278186 459334
rect 278422 459098 278604 459334
rect 278004 423654 278604 459098
rect 278004 423418 278186 423654
rect 278422 423418 278604 423654
rect 278004 423334 278604 423418
rect 278004 423098 278186 423334
rect 278422 423098 278604 423334
rect 278004 387654 278604 423098
rect 278004 387418 278186 387654
rect 278422 387418 278604 387654
rect 278004 387334 278604 387418
rect 278004 387098 278186 387334
rect 278422 387098 278604 387334
rect 278004 351654 278604 387098
rect 278004 351418 278186 351654
rect 278422 351418 278604 351654
rect 278004 351334 278604 351418
rect 278004 351098 278186 351334
rect 278422 351098 278604 351334
rect 278004 315654 278604 351098
rect 278004 315418 278186 315654
rect 278422 315418 278604 315654
rect 278004 315334 278604 315418
rect 278004 315098 278186 315334
rect 278422 315098 278604 315334
rect 278004 279654 278604 315098
rect 278004 279418 278186 279654
rect 278422 279418 278604 279654
rect 278004 279334 278604 279418
rect 278004 279098 278186 279334
rect 278422 279098 278604 279334
rect 278004 243654 278604 279098
rect 278004 243418 278186 243654
rect 278422 243418 278604 243654
rect 278004 243334 278604 243418
rect 278004 243098 278186 243334
rect 278422 243098 278604 243334
rect 278004 207654 278604 243098
rect 278004 207418 278186 207654
rect 278422 207418 278604 207654
rect 278004 207334 278604 207418
rect 278004 207098 278186 207334
rect 278422 207098 278604 207334
rect 278004 171654 278604 207098
rect 278004 171418 278186 171654
rect 278422 171418 278604 171654
rect 278004 171334 278604 171418
rect 278004 171098 278186 171334
rect 278422 171098 278604 171334
rect 278004 135654 278604 171098
rect 278004 135418 278186 135654
rect 278422 135418 278604 135654
rect 278004 135334 278604 135418
rect 278004 135098 278186 135334
rect 278422 135098 278604 135334
rect 278004 99654 278604 135098
rect 278004 99418 278186 99654
rect 278422 99418 278604 99654
rect 278004 99334 278604 99418
rect 278004 99098 278186 99334
rect 278422 99098 278604 99334
rect 278004 63654 278604 99098
rect 278004 63418 278186 63654
rect 278422 63418 278604 63654
rect 278004 63334 278604 63418
rect 278004 63098 278186 63334
rect 278422 63098 278604 63334
rect 278004 27654 278604 63098
rect 278004 27418 278186 27654
rect 278422 27418 278604 27654
rect 278004 27334 278604 27418
rect 278004 27098 278186 27334
rect 278422 27098 278604 27334
rect 278004 -5046 278604 27098
rect 278004 -5282 278186 -5046
rect 278422 -5282 278604 -5046
rect 278004 -5366 278604 -5282
rect 278004 -5602 278186 -5366
rect 278422 -5602 278604 -5366
rect 278004 -5624 278604 -5602
rect 281604 679254 282204 710862
rect 299604 710478 300204 711440
rect 299604 710242 299786 710478
rect 300022 710242 300204 710478
rect 299604 710158 300204 710242
rect 299604 709922 299786 710158
rect 300022 709922 300204 710158
rect 296004 708598 296604 709560
rect 296004 708362 296186 708598
rect 296422 708362 296604 708598
rect 296004 708278 296604 708362
rect 296004 708042 296186 708278
rect 296422 708042 296604 708278
rect 292404 706718 293004 707680
rect 292404 706482 292586 706718
rect 292822 706482 293004 706718
rect 292404 706398 293004 706482
rect 292404 706162 292586 706398
rect 292822 706162 293004 706398
rect 281604 679018 281786 679254
rect 282022 679018 282204 679254
rect 281604 678934 282204 679018
rect 281604 678698 281786 678934
rect 282022 678698 282204 678934
rect 281604 643254 282204 678698
rect 281604 643018 281786 643254
rect 282022 643018 282204 643254
rect 281604 642934 282204 643018
rect 281604 642698 281786 642934
rect 282022 642698 282204 642934
rect 281604 607254 282204 642698
rect 281604 607018 281786 607254
rect 282022 607018 282204 607254
rect 281604 606934 282204 607018
rect 281604 606698 281786 606934
rect 282022 606698 282204 606934
rect 281604 571254 282204 606698
rect 281604 571018 281786 571254
rect 282022 571018 282204 571254
rect 281604 570934 282204 571018
rect 281604 570698 281786 570934
rect 282022 570698 282204 570934
rect 281604 535254 282204 570698
rect 281604 535018 281786 535254
rect 282022 535018 282204 535254
rect 281604 534934 282204 535018
rect 281604 534698 281786 534934
rect 282022 534698 282204 534934
rect 281604 499254 282204 534698
rect 281604 499018 281786 499254
rect 282022 499018 282204 499254
rect 281604 498934 282204 499018
rect 281604 498698 281786 498934
rect 282022 498698 282204 498934
rect 281604 463254 282204 498698
rect 281604 463018 281786 463254
rect 282022 463018 282204 463254
rect 281604 462934 282204 463018
rect 281604 462698 281786 462934
rect 282022 462698 282204 462934
rect 281604 427254 282204 462698
rect 281604 427018 281786 427254
rect 282022 427018 282204 427254
rect 281604 426934 282204 427018
rect 281604 426698 281786 426934
rect 282022 426698 282204 426934
rect 281604 391254 282204 426698
rect 281604 391018 281786 391254
rect 282022 391018 282204 391254
rect 281604 390934 282204 391018
rect 281604 390698 281786 390934
rect 282022 390698 282204 390934
rect 281604 355254 282204 390698
rect 288804 704838 289404 705800
rect 288804 704602 288986 704838
rect 289222 704602 289404 704838
rect 288804 704518 289404 704602
rect 288804 704282 288986 704518
rect 289222 704282 289404 704518
rect 288804 686454 289404 704282
rect 288804 686218 288986 686454
rect 289222 686218 289404 686454
rect 288804 686134 289404 686218
rect 288804 685898 288986 686134
rect 289222 685898 289404 686134
rect 288804 650454 289404 685898
rect 288804 650218 288986 650454
rect 289222 650218 289404 650454
rect 288804 650134 289404 650218
rect 288804 649898 288986 650134
rect 289222 649898 289404 650134
rect 288804 614454 289404 649898
rect 288804 614218 288986 614454
rect 289222 614218 289404 614454
rect 288804 614134 289404 614218
rect 288804 613898 288986 614134
rect 289222 613898 289404 614134
rect 288804 578454 289404 613898
rect 288804 578218 288986 578454
rect 289222 578218 289404 578454
rect 288804 578134 289404 578218
rect 288804 577898 288986 578134
rect 289222 577898 289404 578134
rect 288804 542454 289404 577898
rect 288804 542218 288986 542454
rect 289222 542218 289404 542454
rect 288804 542134 289404 542218
rect 288804 541898 288986 542134
rect 289222 541898 289404 542134
rect 288804 506454 289404 541898
rect 288804 506218 288986 506454
rect 289222 506218 289404 506454
rect 288804 506134 289404 506218
rect 288804 505898 288986 506134
rect 289222 505898 289404 506134
rect 288804 470454 289404 505898
rect 288804 470218 288986 470454
rect 289222 470218 289404 470454
rect 288804 470134 289404 470218
rect 288804 469898 288986 470134
rect 289222 469898 289404 470134
rect 288804 434454 289404 469898
rect 288804 434218 288986 434454
rect 289222 434218 289404 434454
rect 288804 434134 289404 434218
rect 288804 433898 288986 434134
rect 289222 433898 289404 434134
rect 288804 398454 289404 433898
rect 288804 398218 288986 398454
rect 289222 398218 289404 398454
rect 288804 398134 289404 398218
rect 288804 397898 288986 398134
rect 289222 397898 289404 398134
rect 283971 380220 284037 380221
rect 283971 380156 283972 380220
rect 284036 380156 284037 380220
rect 283971 380155 284037 380156
rect 283974 367301 284034 380155
rect 283971 367300 284037 367301
rect 283971 367236 283972 367300
rect 284036 367236 284037 367300
rect 283971 367235 284037 367236
rect 281604 355018 281786 355254
rect 282022 355018 282204 355254
rect 281604 354934 282204 355018
rect 281604 354698 281786 354934
rect 282022 354698 282204 354934
rect 281604 319254 282204 354698
rect 281604 319018 281786 319254
rect 282022 319018 282204 319254
rect 281604 318934 282204 319018
rect 281604 318698 281786 318934
rect 282022 318698 282204 318934
rect 281604 283254 282204 318698
rect 281604 283018 281786 283254
rect 282022 283018 282204 283254
rect 281604 282934 282204 283018
rect 281604 282698 281786 282934
rect 282022 282698 282204 282934
rect 281604 247254 282204 282698
rect 281604 247018 281786 247254
rect 282022 247018 282204 247254
rect 281604 246934 282204 247018
rect 281604 246698 281786 246934
rect 282022 246698 282204 246934
rect 281604 211254 282204 246698
rect 281604 211018 281786 211254
rect 282022 211018 282204 211254
rect 281604 210934 282204 211018
rect 281604 210698 281786 210934
rect 282022 210698 282204 210934
rect 281604 175254 282204 210698
rect 281604 175018 281786 175254
rect 282022 175018 282204 175254
rect 281604 174934 282204 175018
rect 281604 174698 281786 174934
rect 282022 174698 282204 174934
rect 281604 139254 282204 174698
rect 281604 139018 281786 139254
rect 282022 139018 282204 139254
rect 281604 138934 282204 139018
rect 281604 138698 281786 138934
rect 282022 138698 282204 138934
rect 281604 103254 282204 138698
rect 281604 103018 281786 103254
rect 282022 103018 282204 103254
rect 281604 102934 282204 103018
rect 281604 102698 281786 102934
rect 282022 102698 282204 102934
rect 281604 67254 282204 102698
rect 281604 67018 281786 67254
rect 282022 67018 282204 67254
rect 281604 66934 282204 67018
rect 281604 66698 281786 66934
rect 282022 66698 282204 66934
rect 281604 31254 282204 66698
rect 281604 31018 281786 31254
rect 282022 31018 282204 31254
rect 281604 30934 282204 31018
rect 281604 30698 281786 30934
rect 282022 30698 282204 30934
rect 263604 -6222 263786 -5986
rect 264022 -6222 264204 -5986
rect 263604 -6306 264204 -6222
rect 263604 -6542 263786 -6306
rect 264022 -6542 264204 -6306
rect 263604 -7504 264204 -6542
rect 281604 -6926 282204 30698
rect 288804 362454 289404 397898
rect 288804 362218 288986 362454
rect 289222 362218 289404 362454
rect 288804 362134 289404 362218
rect 288804 361898 288986 362134
rect 289222 361898 289404 362134
rect 288804 326454 289404 361898
rect 288804 326218 288986 326454
rect 289222 326218 289404 326454
rect 288804 326134 289404 326218
rect 288804 325898 288986 326134
rect 289222 325898 289404 326134
rect 288804 290454 289404 325898
rect 288804 290218 288986 290454
rect 289222 290218 289404 290454
rect 288804 290134 289404 290218
rect 288804 289898 288986 290134
rect 289222 289898 289404 290134
rect 288804 254454 289404 289898
rect 288804 254218 288986 254454
rect 289222 254218 289404 254454
rect 288804 254134 289404 254218
rect 288804 253898 288986 254134
rect 289222 253898 289404 254134
rect 288804 218454 289404 253898
rect 288804 218218 288986 218454
rect 289222 218218 289404 218454
rect 288804 218134 289404 218218
rect 288804 217898 288986 218134
rect 289222 217898 289404 218134
rect 288804 182454 289404 217898
rect 288804 182218 288986 182454
rect 289222 182218 289404 182454
rect 288804 182134 289404 182218
rect 288804 181898 288986 182134
rect 289222 181898 289404 182134
rect 288804 146454 289404 181898
rect 288804 146218 288986 146454
rect 289222 146218 289404 146454
rect 288804 146134 289404 146218
rect 288804 145898 288986 146134
rect 289222 145898 289404 146134
rect 288804 110454 289404 145898
rect 288804 110218 288986 110454
rect 289222 110218 289404 110454
rect 288804 110134 289404 110218
rect 288804 109898 288986 110134
rect 289222 109898 289404 110134
rect 288804 74454 289404 109898
rect 288804 74218 288986 74454
rect 289222 74218 289404 74454
rect 288804 74134 289404 74218
rect 288804 73898 288986 74134
rect 289222 73898 289404 74134
rect 288804 38454 289404 73898
rect 288804 38218 288986 38454
rect 289222 38218 289404 38454
rect 288804 38134 289404 38218
rect 288804 37898 288986 38134
rect 289222 37898 289404 38134
rect 288804 2454 289404 37898
rect 288804 2218 288986 2454
rect 289222 2218 289404 2454
rect 288804 2134 289404 2218
rect 288804 1898 288986 2134
rect 289222 1898 289404 2134
rect 288804 -346 289404 1898
rect 288804 -582 288986 -346
rect 289222 -582 289404 -346
rect 288804 -666 289404 -582
rect 288804 -902 288986 -666
rect 289222 -902 289404 -666
rect 288804 -1864 289404 -902
rect 292404 690054 293004 706162
rect 292404 689818 292586 690054
rect 292822 689818 293004 690054
rect 292404 689734 293004 689818
rect 292404 689498 292586 689734
rect 292822 689498 293004 689734
rect 292404 654054 293004 689498
rect 292404 653818 292586 654054
rect 292822 653818 293004 654054
rect 292404 653734 293004 653818
rect 292404 653498 292586 653734
rect 292822 653498 293004 653734
rect 292404 618054 293004 653498
rect 292404 617818 292586 618054
rect 292822 617818 293004 618054
rect 292404 617734 293004 617818
rect 292404 617498 292586 617734
rect 292822 617498 293004 617734
rect 292404 582054 293004 617498
rect 292404 581818 292586 582054
rect 292822 581818 293004 582054
rect 292404 581734 293004 581818
rect 292404 581498 292586 581734
rect 292822 581498 293004 581734
rect 292404 546054 293004 581498
rect 292404 545818 292586 546054
rect 292822 545818 293004 546054
rect 292404 545734 293004 545818
rect 292404 545498 292586 545734
rect 292822 545498 293004 545734
rect 292404 510054 293004 545498
rect 292404 509818 292586 510054
rect 292822 509818 293004 510054
rect 292404 509734 293004 509818
rect 292404 509498 292586 509734
rect 292822 509498 293004 509734
rect 292404 474054 293004 509498
rect 292404 473818 292586 474054
rect 292822 473818 293004 474054
rect 292404 473734 293004 473818
rect 292404 473498 292586 473734
rect 292822 473498 293004 473734
rect 292404 438054 293004 473498
rect 292404 437818 292586 438054
rect 292822 437818 293004 438054
rect 292404 437734 293004 437818
rect 292404 437498 292586 437734
rect 292822 437498 293004 437734
rect 292404 402054 293004 437498
rect 292404 401818 292586 402054
rect 292822 401818 293004 402054
rect 292404 401734 293004 401818
rect 292404 401498 292586 401734
rect 292822 401498 293004 401734
rect 292404 366054 293004 401498
rect 292404 365818 292586 366054
rect 292822 365818 293004 366054
rect 292404 365734 293004 365818
rect 292404 365498 292586 365734
rect 292822 365498 293004 365734
rect 292404 330054 293004 365498
rect 292404 329818 292586 330054
rect 292822 329818 293004 330054
rect 292404 329734 293004 329818
rect 292404 329498 292586 329734
rect 292822 329498 293004 329734
rect 292404 294054 293004 329498
rect 292404 293818 292586 294054
rect 292822 293818 293004 294054
rect 292404 293734 293004 293818
rect 292404 293498 292586 293734
rect 292822 293498 293004 293734
rect 292404 258054 293004 293498
rect 292404 257818 292586 258054
rect 292822 257818 293004 258054
rect 292404 257734 293004 257818
rect 292404 257498 292586 257734
rect 292822 257498 293004 257734
rect 292404 222054 293004 257498
rect 292404 221818 292586 222054
rect 292822 221818 293004 222054
rect 292404 221734 293004 221818
rect 292404 221498 292586 221734
rect 292822 221498 293004 221734
rect 292404 186054 293004 221498
rect 292404 185818 292586 186054
rect 292822 185818 293004 186054
rect 292404 185734 293004 185818
rect 292404 185498 292586 185734
rect 292822 185498 293004 185734
rect 292404 150054 293004 185498
rect 292404 149818 292586 150054
rect 292822 149818 293004 150054
rect 292404 149734 293004 149818
rect 292404 149498 292586 149734
rect 292822 149498 293004 149734
rect 292404 114054 293004 149498
rect 292404 113818 292586 114054
rect 292822 113818 293004 114054
rect 292404 113734 293004 113818
rect 292404 113498 292586 113734
rect 292822 113498 293004 113734
rect 292404 78054 293004 113498
rect 292404 77818 292586 78054
rect 292822 77818 293004 78054
rect 292404 77734 293004 77818
rect 292404 77498 292586 77734
rect 292822 77498 293004 77734
rect 292404 42054 293004 77498
rect 292404 41818 292586 42054
rect 292822 41818 293004 42054
rect 292404 41734 293004 41818
rect 292404 41498 292586 41734
rect 292822 41498 293004 41734
rect 292404 6054 293004 41498
rect 292404 5818 292586 6054
rect 292822 5818 293004 6054
rect 292404 5734 293004 5818
rect 292404 5498 292586 5734
rect 292822 5498 293004 5734
rect 292404 -2226 293004 5498
rect 292404 -2462 292586 -2226
rect 292822 -2462 293004 -2226
rect 292404 -2546 293004 -2462
rect 292404 -2782 292586 -2546
rect 292822 -2782 293004 -2546
rect 292404 -3744 293004 -2782
rect 296004 693654 296604 708042
rect 296004 693418 296186 693654
rect 296422 693418 296604 693654
rect 296004 693334 296604 693418
rect 296004 693098 296186 693334
rect 296422 693098 296604 693334
rect 296004 657654 296604 693098
rect 296004 657418 296186 657654
rect 296422 657418 296604 657654
rect 296004 657334 296604 657418
rect 296004 657098 296186 657334
rect 296422 657098 296604 657334
rect 296004 621654 296604 657098
rect 296004 621418 296186 621654
rect 296422 621418 296604 621654
rect 296004 621334 296604 621418
rect 296004 621098 296186 621334
rect 296422 621098 296604 621334
rect 296004 585654 296604 621098
rect 296004 585418 296186 585654
rect 296422 585418 296604 585654
rect 296004 585334 296604 585418
rect 296004 585098 296186 585334
rect 296422 585098 296604 585334
rect 296004 549654 296604 585098
rect 296004 549418 296186 549654
rect 296422 549418 296604 549654
rect 296004 549334 296604 549418
rect 296004 549098 296186 549334
rect 296422 549098 296604 549334
rect 296004 513654 296604 549098
rect 296004 513418 296186 513654
rect 296422 513418 296604 513654
rect 296004 513334 296604 513418
rect 296004 513098 296186 513334
rect 296422 513098 296604 513334
rect 296004 477654 296604 513098
rect 296004 477418 296186 477654
rect 296422 477418 296604 477654
rect 296004 477334 296604 477418
rect 296004 477098 296186 477334
rect 296422 477098 296604 477334
rect 296004 441654 296604 477098
rect 296004 441418 296186 441654
rect 296422 441418 296604 441654
rect 296004 441334 296604 441418
rect 296004 441098 296186 441334
rect 296422 441098 296604 441334
rect 296004 405654 296604 441098
rect 296004 405418 296186 405654
rect 296422 405418 296604 405654
rect 296004 405334 296604 405418
rect 296004 405098 296186 405334
rect 296422 405098 296604 405334
rect 296004 369654 296604 405098
rect 296004 369418 296186 369654
rect 296422 369418 296604 369654
rect 296004 369334 296604 369418
rect 296004 369098 296186 369334
rect 296422 369098 296604 369334
rect 296004 333654 296604 369098
rect 296004 333418 296186 333654
rect 296422 333418 296604 333654
rect 296004 333334 296604 333418
rect 296004 333098 296186 333334
rect 296422 333098 296604 333334
rect 296004 297654 296604 333098
rect 299604 697254 300204 709922
rect 317604 711418 318204 711440
rect 317604 711182 317786 711418
rect 318022 711182 318204 711418
rect 317604 711098 318204 711182
rect 317604 710862 317786 711098
rect 318022 710862 318204 711098
rect 314004 709538 314604 709560
rect 314004 709302 314186 709538
rect 314422 709302 314604 709538
rect 314004 709218 314604 709302
rect 314004 708982 314186 709218
rect 314422 708982 314604 709218
rect 310404 707658 311004 707680
rect 310404 707422 310586 707658
rect 310822 707422 311004 707658
rect 310404 707338 311004 707422
rect 310404 707102 310586 707338
rect 310822 707102 311004 707338
rect 299604 697018 299786 697254
rect 300022 697018 300204 697254
rect 299604 696934 300204 697018
rect 299604 696698 299786 696934
rect 300022 696698 300204 696934
rect 299604 661254 300204 696698
rect 299604 661018 299786 661254
rect 300022 661018 300204 661254
rect 299604 660934 300204 661018
rect 299604 660698 299786 660934
rect 300022 660698 300204 660934
rect 299604 625254 300204 660698
rect 299604 625018 299786 625254
rect 300022 625018 300204 625254
rect 299604 624934 300204 625018
rect 299604 624698 299786 624934
rect 300022 624698 300204 624934
rect 299604 589254 300204 624698
rect 299604 589018 299786 589254
rect 300022 589018 300204 589254
rect 299604 588934 300204 589018
rect 299604 588698 299786 588934
rect 300022 588698 300204 588934
rect 299604 553254 300204 588698
rect 299604 553018 299786 553254
rect 300022 553018 300204 553254
rect 299604 552934 300204 553018
rect 299604 552698 299786 552934
rect 300022 552698 300204 552934
rect 299604 517254 300204 552698
rect 299604 517018 299786 517254
rect 300022 517018 300204 517254
rect 299604 516934 300204 517018
rect 299604 516698 299786 516934
rect 300022 516698 300204 516934
rect 299604 481254 300204 516698
rect 299604 481018 299786 481254
rect 300022 481018 300204 481254
rect 299604 480934 300204 481018
rect 299604 480698 299786 480934
rect 300022 480698 300204 480934
rect 299604 445254 300204 480698
rect 299604 445018 299786 445254
rect 300022 445018 300204 445254
rect 299604 444934 300204 445018
rect 299604 444698 299786 444934
rect 300022 444698 300204 444934
rect 299604 409254 300204 444698
rect 299604 409018 299786 409254
rect 300022 409018 300204 409254
rect 299604 408934 300204 409018
rect 299604 408698 299786 408934
rect 300022 408698 300204 408934
rect 299604 373254 300204 408698
rect 299604 373018 299786 373254
rect 300022 373018 300204 373254
rect 299604 372934 300204 373018
rect 299604 372698 299786 372934
rect 300022 372698 300204 372934
rect 299604 337254 300204 372698
rect 299604 337018 299786 337254
rect 300022 337018 300204 337254
rect 299604 336934 300204 337018
rect 299604 336698 299786 336934
rect 300022 336698 300204 336934
rect 299604 301254 300204 336698
rect 299604 301018 299786 301254
rect 300022 301018 300204 301254
rect 299604 300934 300204 301018
rect 299604 300698 299786 300934
rect 300022 300698 300204 300934
rect 297771 298076 297837 298077
rect 297771 298012 297772 298076
rect 297836 298012 297837 298076
rect 297771 298011 297837 298012
rect 296004 297418 296186 297654
rect 296422 297418 296604 297654
rect 296004 297334 296604 297418
rect 296004 297098 296186 297334
rect 296422 297098 296604 297334
rect 296004 261654 296604 297098
rect 297774 288557 297834 298011
rect 297771 288556 297837 288557
rect 297771 288492 297772 288556
rect 297836 288492 297837 288556
rect 297771 288491 297837 288492
rect 296004 261418 296186 261654
rect 296422 261418 296604 261654
rect 296004 261334 296604 261418
rect 296004 261098 296186 261334
rect 296422 261098 296604 261334
rect 296004 225654 296604 261098
rect 296004 225418 296186 225654
rect 296422 225418 296604 225654
rect 296004 225334 296604 225418
rect 296004 225098 296186 225334
rect 296422 225098 296604 225334
rect 296004 189654 296604 225098
rect 296004 189418 296186 189654
rect 296422 189418 296604 189654
rect 296004 189334 296604 189418
rect 296004 189098 296186 189334
rect 296422 189098 296604 189334
rect 296004 153654 296604 189098
rect 296004 153418 296186 153654
rect 296422 153418 296604 153654
rect 296004 153334 296604 153418
rect 296004 153098 296186 153334
rect 296422 153098 296604 153334
rect 296004 117654 296604 153098
rect 296004 117418 296186 117654
rect 296422 117418 296604 117654
rect 296004 117334 296604 117418
rect 296004 117098 296186 117334
rect 296422 117098 296604 117334
rect 296004 81654 296604 117098
rect 296004 81418 296186 81654
rect 296422 81418 296604 81654
rect 296004 81334 296604 81418
rect 296004 81098 296186 81334
rect 296422 81098 296604 81334
rect 296004 45654 296604 81098
rect 296004 45418 296186 45654
rect 296422 45418 296604 45654
rect 296004 45334 296604 45418
rect 296004 45098 296186 45334
rect 296422 45098 296604 45334
rect 296004 9654 296604 45098
rect 296004 9418 296186 9654
rect 296422 9418 296604 9654
rect 296004 9334 296604 9418
rect 296004 9098 296186 9334
rect 296422 9098 296604 9334
rect 296004 -4106 296604 9098
rect 296004 -4342 296186 -4106
rect 296422 -4342 296604 -4106
rect 296004 -4426 296604 -4342
rect 296004 -4662 296186 -4426
rect 296422 -4662 296604 -4426
rect 296004 -5624 296604 -4662
rect 299604 265254 300204 300698
rect 299604 265018 299786 265254
rect 300022 265018 300204 265254
rect 299604 264934 300204 265018
rect 299604 264698 299786 264934
rect 300022 264698 300204 264934
rect 299604 229254 300204 264698
rect 299604 229018 299786 229254
rect 300022 229018 300204 229254
rect 299604 228934 300204 229018
rect 299604 228698 299786 228934
rect 300022 228698 300204 228934
rect 299604 193254 300204 228698
rect 299604 193018 299786 193254
rect 300022 193018 300204 193254
rect 299604 192934 300204 193018
rect 299604 192698 299786 192934
rect 300022 192698 300204 192934
rect 299604 157254 300204 192698
rect 299604 157018 299786 157254
rect 300022 157018 300204 157254
rect 299604 156934 300204 157018
rect 299604 156698 299786 156934
rect 300022 156698 300204 156934
rect 299604 121254 300204 156698
rect 299604 121018 299786 121254
rect 300022 121018 300204 121254
rect 299604 120934 300204 121018
rect 299604 120698 299786 120934
rect 300022 120698 300204 120934
rect 299604 85254 300204 120698
rect 299604 85018 299786 85254
rect 300022 85018 300204 85254
rect 299604 84934 300204 85018
rect 299604 84698 299786 84934
rect 300022 84698 300204 84934
rect 299604 49254 300204 84698
rect 299604 49018 299786 49254
rect 300022 49018 300204 49254
rect 299604 48934 300204 49018
rect 299604 48698 299786 48934
rect 300022 48698 300204 48934
rect 299604 13254 300204 48698
rect 299604 13018 299786 13254
rect 300022 13018 300204 13254
rect 299604 12934 300204 13018
rect 299604 12698 299786 12934
rect 300022 12698 300204 12934
rect 281604 -7162 281786 -6926
rect 282022 -7162 282204 -6926
rect 281604 -7246 282204 -7162
rect 281604 -7482 281786 -7246
rect 282022 -7482 282204 -7246
rect 281604 -7504 282204 -7482
rect 299604 -5986 300204 12698
rect 306804 705778 307404 705800
rect 306804 705542 306986 705778
rect 307222 705542 307404 705778
rect 306804 705458 307404 705542
rect 306804 705222 306986 705458
rect 307222 705222 307404 705458
rect 306804 668454 307404 705222
rect 306804 668218 306986 668454
rect 307222 668218 307404 668454
rect 306804 668134 307404 668218
rect 306804 667898 306986 668134
rect 307222 667898 307404 668134
rect 306804 632454 307404 667898
rect 306804 632218 306986 632454
rect 307222 632218 307404 632454
rect 306804 632134 307404 632218
rect 306804 631898 306986 632134
rect 307222 631898 307404 632134
rect 306804 596454 307404 631898
rect 306804 596218 306986 596454
rect 307222 596218 307404 596454
rect 306804 596134 307404 596218
rect 306804 595898 306986 596134
rect 307222 595898 307404 596134
rect 306804 560454 307404 595898
rect 306804 560218 306986 560454
rect 307222 560218 307404 560454
rect 306804 560134 307404 560218
rect 306804 559898 306986 560134
rect 307222 559898 307404 560134
rect 306804 524454 307404 559898
rect 306804 524218 306986 524454
rect 307222 524218 307404 524454
rect 306804 524134 307404 524218
rect 306804 523898 306986 524134
rect 307222 523898 307404 524134
rect 306804 488454 307404 523898
rect 306804 488218 306986 488454
rect 307222 488218 307404 488454
rect 306804 488134 307404 488218
rect 306804 487898 306986 488134
rect 307222 487898 307404 488134
rect 306804 452454 307404 487898
rect 306804 452218 306986 452454
rect 307222 452218 307404 452454
rect 306804 452134 307404 452218
rect 306804 451898 306986 452134
rect 307222 451898 307404 452134
rect 306804 416454 307404 451898
rect 306804 416218 306986 416454
rect 307222 416218 307404 416454
rect 306804 416134 307404 416218
rect 306804 415898 306986 416134
rect 307222 415898 307404 416134
rect 306804 380454 307404 415898
rect 306804 380218 306986 380454
rect 307222 380218 307404 380454
rect 306804 380134 307404 380218
rect 306804 379898 306986 380134
rect 307222 379898 307404 380134
rect 306804 344454 307404 379898
rect 306804 344218 306986 344454
rect 307222 344218 307404 344454
rect 306804 344134 307404 344218
rect 306804 343898 306986 344134
rect 307222 343898 307404 344134
rect 306804 308454 307404 343898
rect 306804 308218 306986 308454
rect 307222 308218 307404 308454
rect 306804 308134 307404 308218
rect 306804 307898 306986 308134
rect 307222 307898 307404 308134
rect 306804 272454 307404 307898
rect 306804 272218 306986 272454
rect 307222 272218 307404 272454
rect 306804 272134 307404 272218
rect 306804 271898 306986 272134
rect 307222 271898 307404 272134
rect 306804 236454 307404 271898
rect 306804 236218 306986 236454
rect 307222 236218 307404 236454
rect 306804 236134 307404 236218
rect 306804 235898 306986 236134
rect 307222 235898 307404 236134
rect 306804 200454 307404 235898
rect 306804 200218 306986 200454
rect 307222 200218 307404 200454
rect 306804 200134 307404 200218
rect 306804 199898 306986 200134
rect 307222 199898 307404 200134
rect 306804 164454 307404 199898
rect 306804 164218 306986 164454
rect 307222 164218 307404 164454
rect 306804 164134 307404 164218
rect 306804 163898 306986 164134
rect 307222 163898 307404 164134
rect 306804 128454 307404 163898
rect 306804 128218 306986 128454
rect 307222 128218 307404 128454
rect 306804 128134 307404 128218
rect 306804 127898 306986 128134
rect 307222 127898 307404 128134
rect 306804 92454 307404 127898
rect 306804 92218 306986 92454
rect 307222 92218 307404 92454
rect 306804 92134 307404 92218
rect 306804 91898 306986 92134
rect 307222 91898 307404 92134
rect 306804 56454 307404 91898
rect 306804 56218 306986 56454
rect 307222 56218 307404 56454
rect 306804 56134 307404 56218
rect 306804 55898 306986 56134
rect 307222 55898 307404 56134
rect 306804 20454 307404 55898
rect 306804 20218 306986 20454
rect 307222 20218 307404 20454
rect 306804 20134 307404 20218
rect 306804 19898 306986 20134
rect 307222 19898 307404 20134
rect 306804 -1286 307404 19898
rect 306804 -1522 306986 -1286
rect 307222 -1522 307404 -1286
rect 306804 -1606 307404 -1522
rect 306804 -1842 306986 -1606
rect 307222 -1842 307404 -1606
rect 306804 -1864 307404 -1842
rect 310404 672054 311004 707102
rect 310404 671818 310586 672054
rect 310822 671818 311004 672054
rect 310404 671734 311004 671818
rect 310404 671498 310586 671734
rect 310822 671498 311004 671734
rect 310404 636054 311004 671498
rect 310404 635818 310586 636054
rect 310822 635818 311004 636054
rect 310404 635734 311004 635818
rect 310404 635498 310586 635734
rect 310822 635498 311004 635734
rect 310404 600054 311004 635498
rect 310404 599818 310586 600054
rect 310822 599818 311004 600054
rect 310404 599734 311004 599818
rect 310404 599498 310586 599734
rect 310822 599498 311004 599734
rect 310404 564054 311004 599498
rect 310404 563818 310586 564054
rect 310822 563818 311004 564054
rect 310404 563734 311004 563818
rect 310404 563498 310586 563734
rect 310822 563498 311004 563734
rect 310404 528054 311004 563498
rect 310404 527818 310586 528054
rect 310822 527818 311004 528054
rect 310404 527734 311004 527818
rect 310404 527498 310586 527734
rect 310822 527498 311004 527734
rect 310404 492054 311004 527498
rect 310404 491818 310586 492054
rect 310822 491818 311004 492054
rect 310404 491734 311004 491818
rect 310404 491498 310586 491734
rect 310822 491498 311004 491734
rect 310404 456054 311004 491498
rect 310404 455818 310586 456054
rect 310822 455818 311004 456054
rect 310404 455734 311004 455818
rect 310404 455498 310586 455734
rect 310822 455498 311004 455734
rect 310404 420054 311004 455498
rect 310404 419818 310586 420054
rect 310822 419818 311004 420054
rect 310404 419734 311004 419818
rect 310404 419498 310586 419734
rect 310822 419498 311004 419734
rect 310404 384054 311004 419498
rect 310404 383818 310586 384054
rect 310822 383818 311004 384054
rect 310404 383734 311004 383818
rect 310404 383498 310586 383734
rect 310822 383498 311004 383734
rect 310404 348054 311004 383498
rect 310404 347818 310586 348054
rect 310822 347818 311004 348054
rect 310404 347734 311004 347818
rect 310404 347498 310586 347734
rect 310822 347498 311004 347734
rect 310404 312054 311004 347498
rect 310404 311818 310586 312054
rect 310822 311818 311004 312054
rect 310404 311734 311004 311818
rect 310404 311498 310586 311734
rect 310822 311498 311004 311734
rect 310404 276054 311004 311498
rect 310404 275818 310586 276054
rect 310822 275818 311004 276054
rect 310404 275734 311004 275818
rect 310404 275498 310586 275734
rect 310822 275498 311004 275734
rect 310404 240054 311004 275498
rect 310404 239818 310586 240054
rect 310822 239818 311004 240054
rect 310404 239734 311004 239818
rect 310404 239498 310586 239734
rect 310822 239498 311004 239734
rect 310404 204054 311004 239498
rect 310404 203818 310586 204054
rect 310822 203818 311004 204054
rect 310404 203734 311004 203818
rect 310404 203498 310586 203734
rect 310822 203498 311004 203734
rect 310404 168054 311004 203498
rect 310404 167818 310586 168054
rect 310822 167818 311004 168054
rect 310404 167734 311004 167818
rect 310404 167498 310586 167734
rect 310822 167498 311004 167734
rect 310404 132054 311004 167498
rect 310404 131818 310586 132054
rect 310822 131818 311004 132054
rect 310404 131734 311004 131818
rect 310404 131498 310586 131734
rect 310822 131498 311004 131734
rect 310404 96054 311004 131498
rect 310404 95818 310586 96054
rect 310822 95818 311004 96054
rect 310404 95734 311004 95818
rect 310404 95498 310586 95734
rect 310822 95498 311004 95734
rect 310404 60054 311004 95498
rect 310404 59818 310586 60054
rect 310822 59818 311004 60054
rect 310404 59734 311004 59818
rect 310404 59498 310586 59734
rect 310822 59498 311004 59734
rect 310404 24054 311004 59498
rect 310404 23818 310586 24054
rect 310822 23818 311004 24054
rect 310404 23734 311004 23818
rect 310404 23498 310586 23734
rect 310822 23498 311004 23734
rect 310404 -3166 311004 23498
rect 310404 -3402 310586 -3166
rect 310822 -3402 311004 -3166
rect 310404 -3486 311004 -3402
rect 310404 -3722 310586 -3486
rect 310822 -3722 311004 -3486
rect 310404 -3744 311004 -3722
rect 314004 675654 314604 708982
rect 314004 675418 314186 675654
rect 314422 675418 314604 675654
rect 314004 675334 314604 675418
rect 314004 675098 314186 675334
rect 314422 675098 314604 675334
rect 314004 639654 314604 675098
rect 314004 639418 314186 639654
rect 314422 639418 314604 639654
rect 314004 639334 314604 639418
rect 314004 639098 314186 639334
rect 314422 639098 314604 639334
rect 314004 603654 314604 639098
rect 314004 603418 314186 603654
rect 314422 603418 314604 603654
rect 314004 603334 314604 603418
rect 314004 603098 314186 603334
rect 314422 603098 314604 603334
rect 314004 567654 314604 603098
rect 314004 567418 314186 567654
rect 314422 567418 314604 567654
rect 314004 567334 314604 567418
rect 314004 567098 314186 567334
rect 314422 567098 314604 567334
rect 314004 531654 314604 567098
rect 314004 531418 314186 531654
rect 314422 531418 314604 531654
rect 314004 531334 314604 531418
rect 314004 531098 314186 531334
rect 314422 531098 314604 531334
rect 314004 495654 314604 531098
rect 314004 495418 314186 495654
rect 314422 495418 314604 495654
rect 314004 495334 314604 495418
rect 314004 495098 314186 495334
rect 314422 495098 314604 495334
rect 314004 459654 314604 495098
rect 314004 459418 314186 459654
rect 314422 459418 314604 459654
rect 314004 459334 314604 459418
rect 314004 459098 314186 459334
rect 314422 459098 314604 459334
rect 314004 423654 314604 459098
rect 314004 423418 314186 423654
rect 314422 423418 314604 423654
rect 314004 423334 314604 423418
rect 314004 423098 314186 423334
rect 314422 423098 314604 423334
rect 314004 387654 314604 423098
rect 314004 387418 314186 387654
rect 314422 387418 314604 387654
rect 314004 387334 314604 387418
rect 314004 387098 314186 387334
rect 314422 387098 314604 387334
rect 314004 351654 314604 387098
rect 314004 351418 314186 351654
rect 314422 351418 314604 351654
rect 314004 351334 314604 351418
rect 314004 351098 314186 351334
rect 314422 351098 314604 351334
rect 314004 315654 314604 351098
rect 314004 315418 314186 315654
rect 314422 315418 314604 315654
rect 314004 315334 314604 315418
rect 314004 315098 314186 315334
rect 314422 315098 314604 315334
rect 314004 279654 314604 315098
rect 314004 279418 314186 279654
rect 314422 279418 314604 279654
rect 314004 279334 314604 279418
rect 314004 279098 314186 279334
rect 314422 279098 314604 279334
rect 314004 243654 314604 279098
rect 314004 243418 314186 243654
rect 314422 243418 314604 243654
rect 314004 243334 314604 243418
rect 314004 243098 314186 243334
rect 314422 243098 314604 243334
rect 314004 207654 314604 243098
rect 314004 207418 314186 207654
rect 314422 207418 314604 207654
rect 314004 207334 314604 207418
rect 314004 207098 314186 207334
rect 314422 207098 314604 207334
rect 314004 171654 314604 207098
rect 314004 171418 314186 171654
rect 314422 171418 314604 171654
rect 314004 171334 314604 171418
rect 314004 171098 314186 171334
rect 314422 171098 314604 171334
rect 314004 135654 314604 171098
rect 314004 135418 314186 135654
rect 314422 135418 314604 135654
rect 314004 135334 314604 135418
rect 314004 135098 314186 135334
rect 314422 135098 314604 135334
rect 314004 99654 314604 135098
rect 314004 99418 314186 99654
rect 314422 99418 314604 99654
rect 314004 99334 314604 99418
rect 314004 99098 314186 99334
rect 314422 99098 314604 99334
rect 314004 63654 314604 99098
rect 314004 63418 314186 63654
rect 314422 63418 314604 63654
rect 314004 63334 314604 63418
rect 314004 63098 314186 63334
rect 314422 63098 314604 63334
rect 314004 27654 314604 63098
rect 314004 27418 314186 27654
rect 314422 27418 314604 27654
rect 314004 27334 314604 27418
rect 314004 27098 314186 27334
rect 314422 27098 314604 27334
rect 314004 -5046 314604 27098
rect 314004 -5282 314186 -5046
rect 314422 -5282 314604 -5046
rect 314004 -5366 314604 -5282
rect 314004 -5602 314186 -5366
rect 314422 -5602 314604 -5366
rect 314004 -5624 314604 -5602
rect 317604 679254 318204 710862
rect 335604 710478 336204 711440
rect 335604 710242 335786 710478
rect 336022 710242 336204 710478
rect 335604 710158 336204 710242
rect 335604 709922 335786 710158
rect 336022 709922 336204 710158
rect 332004 708598 332604 709560
rect 332004 708362 332186 708598
rect 332422 708362 332604 708598
rect 332004 708278 332604 708362
rect 332004 708042 332186 708278
rect 332422 708042 332604 708278
rect 328404 706718 329004 707680
rect 328404 706482 328586 706718
rect 328822 706482 329004 706718
rect 328404 706398 329004 706482
rect 328404 706162 328586 706398
rect 328822 706162 329004 706398
rect 317604 679018 317786 679254
rect 318022 679018 318204 679254
rect 317604 678934 318204 679018
rect 317604 678698 317786 678934
rect 318022 678698 318204 678934
rect 317604 643254 318204 678698
rect 317604 643018 317786 643254
rect 318022 643018 318204 643254
rect 317604 642934 318204 643018
rect 317604 642698 317786 642934
rect 318022 642698 318204 642934
rect 317604 607254 318204 642698
rect 317604 607018 317786 607254
rect 318022 607018 318204 607254
rect 317604 606934 318204 607018
rect 317604 606698 317786 606934
rect 318022 606698 318204 606934
rect 317604 571254 318204 606698
rect 317604 571018 317786 571254
rect 318022 571018 318204 571254
rect 317604 570934 318204 571018
rect 317604 570698 317786 570934
rect 318022 570698 318204 570934
rect 317604 535254 318204 570698
rect 317604 535018 317786 535254
rect 318022 535018 318204 535254
rect 317604 534934 318204 535018
rect 317604 534698 317786 534934
rect 318022 534698 318204 534934
rect 317604 499254 318204 534698
rect 317604 499018 317786 499254
rect 318022 499018 318204 499254
rect 317604 498934 318204 499018
rect 317604 498698 317786 498934
rect 318022 498698 318204 498934
rect 317604 463254 318204 498698
rect 317604 463018 317786 463254
rect 318022 463018 318204 463254
rect 317604 462934 318204 463018
rect 317604 462698 317786 462934
rect 318022 462698 318204 462934
rect 317604 427254 318204 462698
rect 317604 427018 317786 427254
rect 318022 427018 318204 427254
rect 317604 426934 318204 427018
rect 317604 426698 317786 426934
rect 318022 426698 318204 426934
rect 317604 391254 318204 426698
rect 317604 391018 317786 391254
rect 318022 391018 318204 391254
rect 317604 390934 318204 391018
rect 317604 390698 317786 390934
rect 318022 390698 318204 390934
rect 317604 355254 318204 390698
rect 317604 355018 317786 355254
rect 318022 355018 318204 355254
rect 317604 354934 318204 355018
rect 317604 354698 317786 354934
rect 318022 354698 318204 354934
rect 317604 319254 318204 354698
rect 317604 319018 317786 319254
rect 318022 319018 318204 319254
rect 317604 318934 318204 319018
rect 317604 318698 317786 318934
rect 318022 318698 318204 318934
rect 317604 283254 318204 318698
rect 317604 283018 317786 283254
rect 318022 283018 318204 283254
rect 317604 282934 318204 283018
rect 317604 282698 317786 282934
rect 318022 282698 318204 282934
rect 317604 247254 318204 282698
rect 317604 247018 317786 247254
rect 318022 247018 318204 247254
rect 317604 246934 318204 247018
rect 317604 246698 317786 246934
rect 318022 246698 318204 246934
rect 317604 211254 318204 246698
rect 317604 211018 317786 211254
rect 318022 211018 318204 211254
rect 317604 210934 318204 211018
rect 317604 210698 317786 210934
rect 318022 210698 318204 210934
rect 317604 175254 318204 210698
rect 317604 175018 317786 175254
rect 318022 175018 318204 175254
rect 317604 174934 318204 175018
rect 317604 174698 317786 174934
rect 318022 174698 318204 174934
rect 317604 139254 318204 174698
rect 317604 139018 317786 139254
rect 318022 139018 318204 139254
rect 317604 138934 318204 139018
rect 317604 138698 317786 138934
rect 318022 138698 318204 138934
rect 317604 103254 318204 138698
rect 317604 103018 317786 103254
rect 318022 103018 318204 103254
rect 317604 102934 318204 103018
rect 317604 102698 317786 102934
rect 318022 102698 318204 102934
rect 317604 67254 318204 102698
rect 317604 67018 317786 67254
rect 318022 67018 318204 67254
rect 317604 66934 318204 67018
rect 317604 66698 317786 66934
rect 318022 66698 318204 66934
rect 317604 31254 318204 66698
rect 317604 31018 317786 31254
rect 318022 31018 318204 31254
rect 317604 30934 318204 31018
rect 317604 30698 317786 30934
rect 318022 30698 318204 30934
rect 299604 -6222 299786 -5986
rect 300022 -6222 300204 -5986
rect 299604 -6306 300204 -6222
rect 299604 -6542 299786 -6306
rect 300022 -6542 300204 -6306
rect 299604 -7504 300204 -6542
rect 317604 -6926 318204 30698
rect 324804 704838 325404 705800
rect 324804 704602 324986 704838
rect 325222 704602 325404 704838
rect 324804 704518 325404 704602
rect 324804 704282 324986 704518
rect 325222 704282 325404 704518
rect 324804 686454 325404 704282
rect 324804 686218 324986 686454
rect 325222 686218 325404 686454
rect 324804 686134 325404 686218
rect 324804 685898 324986 686134
rect 325222 685898 325404 686134
rect 324804 650454 325404 685898
rect 324804 650218 324986 650454
rect 325222 650218 325404 650454
rect 324804 650134 325404 650218
rect 324804 649898 324986 650134
rect 325222 649898 325404 650134
rect 324804 614454 325404 649898
rect 324804 614218 324986 614454
rect 325222 614218 325404 614454
rect 324804 614134 325404 614218
rect 324804 613898 324986 614134
rect 325222 613898 325404 614134
rect 324804 578454 325404 613898
rect 324804 578218 324986 578454
rect 325222 578218 325404 578454
rect 324804 578134 325404 578218
rect 324804 577898 324986 578134
rect 325222 577898 325404 578134
rect 324804 542454 325404 577898
rect 324804 542218 324986 542454
rect 325222 542218 325404 542454
rect 324804 542134 325404 542218
rect 324804 541898 324986 542134
rect 325222 541898 325404 542134
rect 324804 506454 325404 541898
rect 324804 506218 324986 506454
rect 325222 506218 325404 506454
rect 324804 506134 325404 506218
rect 324804 505898 324986 506134
rect 325222 505898 325404 506134
rect 324804 470454 325404 505898
rect 324804 470218 324986 470454
rect 325222 470218 325404 470454
rect 324804 470134 325404 470218
rect 324804 469898 324986 470134
rect 325222 469898 325404 470134
rect 324804 434454 325404 469898
rect 324804 434218 324986 434454
rect 325222 434218 325404 434454
rect 324804 434134 325404 434218
rect 324804 433898 324986 434134
rect 325222 433898 325404 434134
rect 324804 398454 325404 433898
rect 324804 398218 324986 398454
rect 325222 398218 325404 398454
rect 324804 398134 325404 398218
rect 324804 397898 324986 398134
rect 325222 397898 325404 398134
rect 324804 362454 325404 397898
rect 324804 362218 324986 362454
rect 325222 362218 325404 362454
rect 324804 362134 325404 362218
rect 324804 361898 324986 362134
rect 325222 361898 325404 362134
rect 324804 326454 325404 361898
rect 324804 326218 324986 326454
rect 325222 326218 325404 326454
rect 324804 326134 325404 326218
rect 324804 325898 324986 326134
rect 325222 325898 325404 326134
rect 324804 290454 325404 325898
rect 324804 290218 324986 290454
rect 325222 290218 325404 290454
rect 324804 290134 325404 290218
rect 324804 289898 324986 290134
rect 325222 289898 325404 290134
rect 324804 254454 325404 289898
rect 324804 254218 324986 254454
rect 325222 254218 325404 254454
rect 324804 254134 325404 254218
rect 324804 253898 324986 254134
rect 325222 253898 325404 254134
rect 324804 218454 325404 253898
rect 324804 218218 324986 218454
rect 325222 218218 325404 218454
rect 324804 218134 325404 218218
rect 324804 217898 324986 218134
rect 325222 217898 325404 218134
rect 324804 182454 325404 217898
rect 324804 182218 324986 182454
rect 325222 182218 325404 182454
rect 324804 182134 325404 182218
rect 324804 181898 324986 182134
rect 325222 181898 325404 182134
rect 324804 146454 325404 181898
rect 324804 146218 324986 146454
rect 325222 146218 325404 146454
rect 324804 146134 325404 146218
rect 324804 145898 324986 146134
rect 325222 145898 325404 146134
rect 324804 110454 325404 145898
rect 324804 110218 324986 110454
rect 325222 110218 325404 110454
rect 324804 110134 325404 110218
rect 324804 109898 324986 110134
rect 325222 109898 325404 110134
rect 324804 74454 325404 109898
rect 324804 74218 324986 74454
rect 325222 74218 325404 74454
rect 324804 74134 325404 74218
rect 324804 73898 324986 74134
rect 325222 73898 325404 74134
rect 324804 38454 325404 73898
rect 324804 38218 324986 38454
rect 325222 38218 325404 38454
rect 324804 38134 325404 38218
rect 324804 37898 324986 38134
rect 325222 37898 325404 38134
rect 324804 2454 325404 37898
rect 324804 2218 324986 2454
rect 325222 2218 325404 2454
rect 324804 2134 325404 2218
rect 324804 1898 324986 2134
rect 325222 1898 325404 2134
rect 324804 -346 325404 1898
rect 324804 -582 324986 -346
rect 325222 -582 325404 -346
rect 324804 -666 325404 -582
rect 324804 -902 324986 -666
rect 325222 -902 325404 -666
rect 324804 -1864 325404 -902
rect 328404 690054 329004 706162
rect 328404 689818 328586 690054
rect 328822 689818 329004 690054
rect 328404 689734 329004 689818
rect 328404 689498 328586 689734
rect 328822 689498 329004 689734
rect 328404 654054 329004 689498
rect 328404 653818 328586 654054
rect 328822 653818 329004 654054
rect 328404 653734 329004 653818
rect 328404 653498 328586 653734
rect 328822 653498 329004 653734
rect 328404 618054 329004 653498
rect 328404 617818 328586 618054
rect 328822 617818 329004 618054
rect 328404 617734 329004 617818
rect 328404 617498 328586 617734
rect 328822 617498 329004 617734
rect 328404 582054 329004 617498
rect 328404 581818 328586 582054
rect 328822 581818 329004 582054
rect 328404 581734 329004 581818
rect 328404 581498 328586 581734
rect 328822 581498 329004 581734
rect 328404 546054 329004 581498
rect 328404 545818 328586 546054
rect 328822 545818 329004 546054
rect 328404 545734 329004 545818
rect 328404 545498 328586 545734
rect 328822 545498 329004 545734
rect 328404 510054 329004 545498
rect 328404 509818 328586 510054
rect 328822 509818 329004 510054
rect 328404 509734 329004 509818
rect 328404 509498 328586 509734
rect 328822 509498 329004 509734
rect 328404 474054 329004 509498
rect 328404 473818 328586 474054
rect 328822 473818 329004 474054
rect 328404 473734 329004 473818
rect 328404 473498 328586 473734
rect 328822 473498 329004 473734
rect 328404 438054 329004 473498
rect 328404 437818 328586 438054
rect 328822 437818 329004 438054
rect 328404 437734 329004 437818
rect 328404 437498 328586 437734
rect 328822 437498 329004 437734
rect 328404 402054 329004 437498
rect 328404 401818 328586 402054
rect 328822 401818 329004 402054
rect 328404 401734 329004 401818
rect 328404 401498 328586 401734
rect 328822 401498 329004 401734
rect 328404 366054 329004 401498
rect 328404 365818 328586 366054
rect 328822 365818 329004 366054
rect 328404 365734 329004 365818
rect 328404 365498 328586 365734
rect 328822 365498 329004 365734
rect 328404 330054 329004 365498
rect 328404 329818 328586 330054
rect 328822 329818 329004 330054
rect 328404 329734 329004 329818
rect 328404 329498 328586 329734
rect 328822 329498 329004 329734
rect 328404 294054 329004 329498
rect 328404 293818 328586 294054
rect 328822 293818 329004 294054
rect 328404 293734 329004 293818
rect 328404 293498 328586 293734
rect 328822 293498 329004 293734
rect 328404 258054 329004 293498
rect 328404 257818 328586 258054
rect 328822 257818 329004 258054
rect 328404 257734 329004 257818
rect 328404 257498 328586 257734
rect 328822 257498 329004 257734
rect 328404 222054 329004 257498
rect 328404 221818 328586 222054
rect 328822 221818 329004 222054
rect 328404 221734 329004 221818
rect 328404 221498 328586 221734
rect 328822 221498 329004 221734
rect 328404 186054 329004 221498
rect 328404 185818 328586 186054
rect 328822 185818 329004 186054
rect 328404 185734 329004 185818
rect 328404 185498 328586 185734
rect 328822 185498 329004 185734
rect 328404 150054 329004 185498
rect 328404 149818 328586 150054
rect 328822 149818 329004 150054
rect 328404 149734 329004 149818
rect 328404 149498 328586 149734
rect 328822 149498 329004 149734
rect 328404 114054 329004 149498
rect 328404 113818 328586 114054
rect 328822 113818 329004 114054
rect 328404 113734 329004 113818
rect 328404 113498 328586 113734
rect 328822 113498 329004 113734
rect 328404 78054 329004 113498
rect 328404 77818 328586 78054
rect 328822 77818 329004 78054
rect 328404 77734 329004 77818
rect 328404 77498 328586 77734
rect 328822 77498 329004 77734
rect 328404 42054 329004 77498
rect 328404 41818 328586 42054
rect 328822 41818 329004 42054
rect 328404 41734 329004 41818
rect 328404 41498 328586 41734
rect 328822 41498 329004 41734
rect 328404 6054 329004 41498
rect 328404 5818 328586 6054
rect 328822 5818 329004 6054
rect 328404 5734 329004 5818
rect 328404 5498 328586 5734
rect 328822 5498 329004 5734
rect 328404 -2226 329004 5498
rect 328404 -2462 328586 -2226
rect 328822 -2462 329004 -2226
rect 328404 -2546 329004 -2462
rect 328404 -2782 328586 -2546
rect 328822 -2782 329004 -2546
rect 328404 -3744 329004 -2782
rect 332004 693654 332604 708042
rect 332004 693418 332186 693654
rect 332422 693418 332604 693654
rect 332004 693334 332604 693418
rect 332004 693098 332186 693334
rect 332422 693098 332604 693334
rect 332004 657654 332604 693098
rect 332004 657418 332186 657654
rect 332422 657418 332604 657654
rect 332004 657334 332604 657418
rect 332004 657098 332186 657334
rect 332422 657098 332604 657334
rect 332004 621654 332604 657098
rect 332004 621418 332186 621654
rect 332422 621418 332604 621654
rect 332004 621334 332604 621418
rect 332004 621098 332186 621334
rect 332422 621098 332604 621334
rect 332004 585654 332604 621098
rect 332004 585418 332186 585654
rect 332422 585418 332604 585654
rect 332004 585334 332604 585418
rect 332004 585098 332186 585334
rect 332422 585098 332604 585334
rect 332004 549654 332604 585098
rect 332004 549418 332186 549654
rect 332422 549418 332604 549654
rect 332004 549334 332604 549418
rect 332004 549098 332186 549334
rect 332422 549098 332604 549334
rect 332004 513654 332604 549098
rect 332004 513418 332186 513654
rect 332422 513418 332604 513654
rect 332004 513334 332604 513418
rect 332004 513098 332186 513334
rect 332422 513098 332604 513334
rect 332004 477654 332604 513098
rect 332004 477418 332186 477654
rect 332422 477418 332604 477654
rect 332004 477334 332604 477418
rect 332004 477098 332186 477334
rect 332422 477098 332604 477334
rect 332004 441654 332604 477098
rect 332004 441418 332186 441654
rect 332422 441418 332604 441654
rect 332004 441334 332604 441418
rect 332004 441098 332186 441334
rect 332422 441098 332604 441334
rect 332004 405654 332604 441098
rect 332004 405418 332186 405654
rect 332422 405418 332604 405654
rect 332004 405334 332604 405418
rect 332004 405098 332186 405334
rect 332422 405098 332604 405334
rect 332004 369654 332604 405098
rect 332004 369418 332186 369654
rect 332422 369418 332604 369654
rect 332004 369334 332604 369418
rect 332004 369098 332186 369334
rect 332422 369098 332604 369334
rect 332004 333654 332604 369098
rect 332004 333418 332186 333654
rect 332422 333418 332604 333654
rect 332004 333334 332604 333418
rect 332004 333098 332186 333334
rect 332422 333098 332604 333334
rect 332004 297654 332604 333098
rect 332004 297418 332186 297654
rect 332422 297418 332604 297654
rect 332004 297334 332604 297418
rect 332004 297098 332186 297334
rect 332422 297098 332604 297334
rect 332004 261654 332604 297098
rect 332004 261418 332186 261654
rect 332422 261418 332604 261654
rect 332004 261334 332604 261418
rect 332004 261098 332186 261334
rect 332422 261098 332604 261334
rect 332004 225654 332604 261098
rect 332004 225418 332186 225654
rect 332422 225418 332604 225654
rect 332004 225334 332604 225418
rect 332004 225098 332186 225334
rect 332422 225098 332604 225334
rect 332004 189654 332604 225098
rect 332004 189418 332186 189654
rect 332422 189418 332604 189654
rect 332004 189334 332604 189418
rect 332004 189098 332186 189334
rect 332422 189098 332604 189334
rect 332004 153654 332604 189098
rect 332004 153418 332186 153654
rect 332422 153418 332604 153654
rect 332004 153334 332604 153418
rect 332004 153098 332186 153334
rect 332422 153098 332604 153334
rect 332004 117654 332604 153098
rect 332004 117418 332186 117654
rect 332422 117418 332604 117654
rect 332004 117334 332604 117418
rect 332004 117098 332186 117334
rect 332422 117098 332604 117334
rect 332004 81654 332604 117098
rect 332004 81418 332186 81654
rect 332422 81418 332604 81654
rect 332004 81334 332604 81418
rect 332004 81098 332186 81334
rect 332422 81098 332604 81334
rect 332004 45654 332604 81098
rect 332004 45418 332186 45654
rect 332422 45418 332604 45654
rect 332004 45334 332604 45418
rect 332004 45098 332186 45334
rect 332422 45098 332604 45334
rect 332004 9654 332604 45098
rect 332004 9418 332186 9654
rect 332422 9418 332604 9654
rect 332004 9334 332604 9418
rect 332004 9098 332186 9334
rect 332422 9098 332604 9334
rect 332004 -4106 332604 9098
rect 332004 -4342 332186 -4106
rect 332422 -4342 332604 -4106
rect 332004 -4426 332604 -4342
rect 332004 -4662 332186 -4426
rect 332422 -4662 332604 -4426
rect 332004 -5624 332604 -4662
rect 335604 697254 336204 709922
rect 353604 711418 354204 711440
rect 353604 711182 353786 711418
rect 354022 711182 354204 711418
rect 353604 711098 354204 711182
rect 353604 710862 353786 711098
rect 354022 710862 354204 711098
rect 350004 709538 350604 709560
rect 350004 709302 350186 709538
rect 350422 709302 350604 709538
rect 350004 709218 350604 709302
rect 350004 708982 350186 709218
rect 350422 708982 350604 709218
rect 346404 707658 347004 707680
rect 346404 707422 346586 707658
rect 346822 707422 347004 707658
rect 346404 707338 347004 707422
rect 346404 707102 346586 707338
rect 346822 707102 347004 707338
rect 335604 697018 335786 697254
rect 336022 697018 336204 697254
rect 335604 696934 336204 697018
rect 335604 696698 335786 696934
rect 336022 696698 336204 696934
rect 335604 661254 336204 696698
rect 335604 661018 335786 661254
rect 336022 661018 336204 661254
rect 335604 660934 336204 661018
rect 335604 660698 335786 660934
rect 336022 660698 336204 660934
rect 335604 625254 336204 660698
rect 335604 625018 335786 625254
rect 336022 625018 336204 625254
rect 335604 624934 336204 625018
rect 335604 624698 335786 624934
rect 336022 624698 336204 624934
rect 335604 589254 336204 624698
rect 335604 589018 335786 589254
rect 336022 589018 336204 589254
rect 335604 588934 336204 589018
rect 335604 588698 335786 588934
rect 336022 588698 336204 588934
rect 335604 553254 336204 588698
rect 335604 553018 335786 553254
rect 336022 553018 336204 553254
rect 335604 552934 336204 553018
rect 335604 552698 335786 552934
rect 336022 552698 336204 552934
rect 335604 517254 336204 552698
rect 335604 517018 335786 517254
rect 336022 517018 336204 517254
rect 335604 516934 336204 517018
rect 335604 516698 335786 516934
rect 336022 516698 336204 516934
rect 335604 481254 336204 516698
rect 335604 481018 335786 481254
rect 336022 481018 336204 481254
rect 335604 480934 336204 481018
rect 335604 480698 335786 480934
rect 336022 480698 336204 480934
rect 335604 445254 336204 480698
rect 335604 445018 335786 445254
rect 336022 445018 336204 445254
rect 335604 444934 336204 445018
rect 335604 444698 335786 444934
rect 336022 444698 336204 444934
rect 335604 409254 336204 444698
rect 335604 409018 335786 409254
rect 336022 409018 336204 409254
rect 335604 408934 336204 409018
rect 335604 408698 335786 408934
rect 336022 408698 336204 408934
rect 335604 373254 336204 408698
rect 335604 373018 335786 373254
rect 336022 373018 336204 373254
rect 335604 372934 336204 373018
rect 335604 372698 335786 372934
rect 336022 372698 336204 372934
rect 335604 337254 336204 372698
rect 335604 337018 335786 337254
rect 336022 337018 336204 337254
rect 335604 336934 336204 337018
rect 335604 336698 335786 336934
rect 336022 336698 336204 336934
rect 335604 301254 336204 336698
rect 335604 301018 335786 301254
rect 336022 301018 336204 301254
rect 335604 300934 336204 301018
rect 335604 300698 335786 300934
rect 336022 300698 336204 300934
rect 335604 265254 336204 300698
rect 335604 265018 335786 265254
rect 336022 265018 336204 265254
rect 335604 264934 336204 265018
rect 335604 264698 335786 264934
rect 336022 264698 336204 264934
rect 335604 229254 336204 264698
rect 335604 229018 335786 229254
rect 336022 229018 336204 229254
rect 335604 228934 336204 229018
rect 335604 228698 335786 228934
rect 336022 228698 336204 228934
rect 335604 193254 336204 228698
rect 335604 193018 335786 193254
rect 336022 193018 336204 193254
rect 335604 192934 336204 193018
rect 335604 192698 335786 192934
rect 336022 192698 336204 192934
rect 335604 157254 336204 192698
rect 335604 157018 335786 157254
rect 336022 157018 336204 157254
rect 335604 156934 336204 157018
rect 335604 156698 335786 156934
rect 336022 156698 336204 156934
rect 335604 121254 336204 156698
rect 335604 121018 335786 121254
rect 336022 121018 336204 121254
rect 335604 120934 336204 121018
rect 335604 120698 335786 120934
rect 336022 120698 336204 120934
rect 335604 85254 336204 120698
rect 335604 85018 335786 85254
rect 336022 85018 336204 85254
rect 335604 84934 336204 85018
rect 335604 84698 335786 84934
rect 336022 84698 336204 84934
rect 335604 49254 336204 84698
rect 335604 49018 335786 49254
rect 336022 49018 336204 49254
rect 335604 48934 336204 49018
rect 335604 48698 335786 48934
rect 336022 48698 336204 48934
rect 335604 13254 336204 48698
rect 335604 13018 335786 13254
rect 336022 13018 336204 13254
rect 335604 12934 336204 13018
rect 335604 12698 335786 12934
rect 336022 12698 336204 12934
rect 317604 -7162 317786 -6926
rect 318022 -7162 318204 -6926
rect 317604 -7246 318204 -7162
rect 317604 -7482 317786 -7246
rect 318022 -7482 318204 -7246
rect 317604 -7504 318204 -7482
rect 335604 -5986 336204 12698
rect 342804 705778 343404 705800
rect 342804 705542 342986 705778
rect 343222 705542 343404 705778
rect 342804 705458 343404 705542
rect 342804 705222 342986 705458
rect 343222 705222 343404 705458
rect 342804 668454 343404 705222
rect 342804 668218 342986 668454
rect 343222 668218 343404 668454
rect 342804 668134 343404 668218
rect 342804 667898 342986 668134
rect 343222 667898 343404 668134
rect 342804 632454 343404 667898
rect 342804 632218 342986 632454
rect 343222 632218 343404 632454
rect 342804 632134 343404 632218
rect 342804 631898 342986 632134
rect 343222 631898 343404 632134
rect 342804 596454 343404 631898
rect 342804 596218 342986 596454
rect 343222 596218 343404 596454
rect 342804 596134 343404 596218
rect 342804 595898 342986 596134
rect 343222 595898 343404 596134
rect 342804 560454 343404 595898
rect 342804 560218 342986 560454
rect 343222 560218 343404 560454
rect 342804 560134 343404 560218
rect 342804 559898 342986 560134
rect 343222 559898 343404 560134
rect 342804 524454 343404 559898
rect 342804 524218 342986 524454
rect 343222 524218 343404 524454
rect 342804 524134 343404 524218
rect 342804 523898 342986 524134
rect 343222 523898 343404 524134
rect 342804 488454 343404 523898
rect 342804 488218 342986 488454
rect 343222 488218 343404 488454
rect 342804 488134 343404 488218
rect 342804 487898 342986 488134
rect 343222 487898 343404 488134
rect 342804 452454 343404 487898
rect 342804 452218 342986 452454
rect 343222 452218 343404 452454
rect 342804 452134 343404 452218
rect 342804 451898 342986 452134
rect 343222 451898 343404 452134
rect 342804 416454 343404 451898
rect 342804 416218 342986 416454
rect 343222 416218 343404 416454
rect 342804 416134 343404 416218
rect 342804 415898 342986 416134
rect 343222 415898 343404 416134
rect 342804 380454 343404 415898
rect 342804 380218 342986 380454
rect 343222 380218 343404 380454
rect 342804 380134 343404 380218
rect 342804 379898 342986 380134
rect 343222 379898 343404 380134
rect 342804 344454 343404 379898
rect 342804 344218 342986 344454
rect 343222 344218 343404 344454
rect 342804 344134 343404 344218
rect 342804 343898 342986 344134
rect 343222 343898 343404 344134
rect 342804 308454 343404 343898
rect 342804 308218 342986 308454
rect 343222 308218 343404 308454
rect 342804 308134 343404 308218
rect 342804 307898 342986 308134
rect 343222 307898 343404 308134
rect 342804 272454 343404 307898
rect 342804 272218 342986 272454
rect 343222 272218 343404 272454
rect 342804 272134 343404 272218
rect 342804 271898 342986 272134
rect 343222 271898 343404 272134
rect 342804 236454 343404 271898
rect 342804 236218 342986 236454
rect 343222 236218 343404 236454
rect 342804 236134 343404 236218
rect 342804 235898 342986 236134
rect 343222 235898 343404 236134
rect 342804 200454 343404 235898
rect 342804 200218 342986 200454
rect 343222 200218 343404 200454
rect 342804 200134 343404 200218
rect 342804 199898 342986 200134
rect 343222 199898 343404 200134
rect 342804 164454 343404 199898
rect 342804 164218 342986 164454
rect 343222 164218 343404 164454
rect 342804 164134 343404 164218
rect 342804 163898 342986 164134
rect 343222 163898 343404 164134
rect 342804 128454 343404 163898
rect 342804 128218 342986 128454
rect 343222 128218 343404 128454
rect 342804 128134 343404 128218
rect 342804 127898 342986 128134
rect 343222 127898 343404 128134
rect 342804 92454 343404 127898
rect 342804 92218 342986 92454
rect 343222 92218 343404 92454
rect 342804 92134 343404 92218
rect 342804 91898 342986 92134
rect 343222 91898 343404 92134
rect 342804 56454 343404 91898
rect 342804 56218 342986 56454
rect 343222 56218 343404 56454
rect 342804 56134 343404 56218
rect 342804 55898 342986 56134
rect 343222 55898 343404 56134
rect 342804 20454 343404 55898
rect 342804 20218 342986 20454
rect 343222 20218 343404 20454
rect 342804 20134 343404 20218
rect 342804 19898 342986 20134
rect 343222 19898 343404 20134
rect 342804 -1286 343404 19898
rect 342804 -1522 342986 -1286
rect 343222 -1522 343404 -1286
rect 342804 -1606 343404 -1522
rect 342804 -1842 342986 -1606
rect 343222 -1842 343404 -1606
rect 342804 -1864 343404 -1842
rect 346404 672054 347004 707102
rect 346404 671818 346586 672054
rect 346822 671818 347004 672054
rect 346404 671734 347004 671818
rect 346404 671498 346586 671734
rect 346822 671498 347004 671734
rect 346404 636054 347004 671498
rect 346404 635818 346586 636054
rect 346822 635818 347004 636054
rect 346404 635734 347004 635818
rect 346404 635498 346586 635734
rect 346822 635498 347004 635734
rect 346404 600054 347004 635498
rect 346404 599818 346586 600054
rect 346822 599818 347004 600054
rect 346404 599734 347004 599818
rect 346404 599498 346586 599734
rect 346822 599498 347004 599734
rect 346404 564054 347004 599498
rect 346404 563818 346586 564054
rect 346822 563818 347004 564054
rect 346404 563734 347004 563818
rect 346404 563498 346586 563734
rect 346822 563498 347004 563734
rect 346404 528054 347004 563498
rect 346404 527818 346586 528054
rect 346822 527818 347004 528054
rect 346404 527734 347004 527818
rect 346404 527498 346586 527734
rect 346822 527498 347004 527734
rect 346404 492054 347004 527498
rect 346404 491818 346586 492054
rect 346822 491818 347004 492054
rect 346404 491734 347004 491818
rect 346404 491498 346586 491734
rect 346822 491498 347004 491734
rect 346404 456054 347004 491498
rect 346404 455818 346586 456054
rect 346822 455818 347004 456054
rect 346404 455734 347004 455818
rect 346404 455498 346586 455734
rect 346822 455498 347004 455734
rect 346404 420054 347004 455498
rect 346404 419818 346586 420054
rect 346822 419818 347004 420054
rect 346404 419734 347004 419818
rect 346404 419498 346586 419734
rect 346822 419498 347004 419734
rect 346404 384054 347004 419498
rect 346404 383818 346586 384054
rect 346822 383818 347004 384054
rect 346404 383734 347004 383818
rect 346404 383498 346586 383734
rect 346822 383498 347004 383734
rect 346404 348054 347004 383498
rect 346404 347818 346586 348054
rect 346822 347818 347004 348054
rect 346404 347734 347004 347818
rect 346404 347498 346586 347734
rect 346822 347498 347004 347734
rect 346404 312054 347004 347498
rect 346404 311818 346586 312054
rect 346822 311818 347004 312054
rect 346404 311734 347004 311818
rect 346404 311498 346586 311734
rect 346822 311498 347004 311734
rect 346404 276054 347004 311498
rect 346404 275818 346586 276054
rect 346822 275818 347004 276054
rect 346404 275734 347004 275818
rect 346404 275498 346586 275734
rect 346822 275498 347004 275734
rect 346404 240054 347004 275498
rect 346404 239818 346586 240054
rect 346822 239818 347004 240054
rect 346404 239734 347004 239818
rect 346404 239498 346586 239734
rect 346822 239498 347004 239734
rect 346404 204054 347004 239498
rect 346404 203818 346586 204054
rect 346822 203818 347004 204054
rect 346404 203734 347004 203818
rect 346404 203498 346586 203734
rect 346822 203498 347004 203734
rect 346404 168054 347004 203498
rect 346404 167818 346586 168054
rect 346822 167818 347004 168054
rect 346404 167734 347004 167818
rect 346404 167498 346586 167734
rect 346822 167498 347004 167734
rect 346404 132054 347004 167498
rect 346404 131818 346586 132054
rect 346822 131818 347004 132054
rect 346404 131734 347004 131818
rect 346404 131498 346586 131734
rect 346822 131498 347004 131734
rect 346404 96054 347004 131498
rect 346404 95818 346586 96054
rect 346822 95818 347004 96054
rect 346404 95734 347004 95818
rect 346404 95498 346586 95734
rect 346822 95498 347004 95734
rect 346404 60054 347004 95498
rect 346404 59818 346586 60054
rect 346822 59818 347004 60054
rect 346404 59734 347004 59818
rect 346404 59498 346586 59734
rect 346822 59498 347004 59734
rect 346404 24054 347004 59498
rect 346404 23818 346586 24054
rect 346822 23818 347004 24054
rect 346404 23734 347004 23818
rect 346404 23498 346586 23734
rect 346822 23498 347004 23734
rect 346404 -3166 347004 23498
rect 346404 -3402 346586 -3166
rect 346822 -3402 347004 -3166
rect 346404 -3486 347004 -3402
rect 346404 -3722 346586 -3486
rect 346822 -3722 347004 -3486
rect 346404 -3744 347004 -3722
rect 350004 675654 350604 708982
rect 350004 675418 350186 675654
rect 350422 675418 350604 675654
rect 350004 675334 350604 675418
rect 350004 675098 350186 675334
rect 350422 675098 350604 675334
rect 350004 639654 350604 675098
rect 350004 639418 350186 639654
rect 350422 639418 350604 639654
rect 350004 639334 350604 639418
rect 350004 639098 350186 639334
rect 350422 639098 350604 639334
rect 350004 603654 350604 639098
rect 350004 603418 350186 603654
rect 350422 603418 350604 603654
rect 350004 603334 350604 603418
rect 350004 603098 350186 603334
rect 350422 603098 350604 603334
rect 350004 567654 350604 603098
rect 350004 567418 350186 567654
rect 350422 567418 350604 567654
rect 350004 567334 350604 567418
rect 350004 567098 350186 567334
rect 350422 567098 350604 567334
rect 350004 531654 350604 567098
rect 350004 531418 350186 531654
rect 350422 531418 350604 531654
rect 350004 531334 350604 531418
rect 350004 531098 350186 531334
rect 350422 531098 350604 531334
rect 350004 495654 350604 531098
rect 350004 495418 350186 495654
rect 350422 495418 350604 495654
rect 350004 495334 350604 495418
rect 350004 495098 350186 495334
rect 350422 495098 350604 495334
rect 350004 459654 350604 495098
rect 350004 459418 350186 459654
rect 350422 459418 350604 459654
rect 350004 459334 350604 459418
rect 350004 459098 350186 459334
rect 350422 459098 350604 459334
rect 350004 423654 350604 459098
rect 350004 423418 350186 423654
rect 350422 423418 350604 423654
rect 350004 423334 350604 423418
rect 350004 423098 350186 423334
rect 350422 423098 350604 423334
rect 350004 387654 350604 423098
rect 350004 387418 350186 387654
rect 350422 387418 350604 387654
rect 350004 387334 350604 387418
rect 350004 387098 350186 387334
rect 350422 387098 350604 387334
rect 350004 351654 350604 387098
rect 350004 351418 350186 351654
rect 350422 351418 350604 351654
rect 350004 351334 350604 351418
rect 350004 351098 350186 351334
rect 350422 351098 350604 351334
rect 350004 315654 350604 351098
rect 350004 315418 350186 315654
rect 350422 315418 350604 315654
rect 350004 315334 350604 315418
rect 350004 315098 350186 315334
rect 350422 315098 350604 315334
rect 350004 279654 350604 315098
rect 350004 279418 350186 279654
rect 350422 279418 350604 279654
rect 350004 279334 350604 279418
rect 350004 279098 350186 279334
rect 350422 279098 350604 279334
rect 350004 243654 350604 279098
rect 350004 243418 350186 243654
rect 350422 243418 350604 243654
rect 350004 243334 350604 243418
rect 350004 243098 350186 243334
rect 350422 243098 350604 243334
rect 350004 207654 350604 243098
rect 350004 207418 350186 207654
rect 350422 207418 350604 207654
rect 350004 207334 350604 207418
rect 350004 207098 350186 207334
rect 350422 207098 350604 207334
rect 350004 171654 350604 207098
rect 350004 171418 350186 171654
rect 350422 171418 350604 171654
rect 350004 171334 350604 171418
rect 350004 171098 350186 171334
rect 350422 171098 350604 171334
rect 350004 135654 350604 171098
rect 350004 135418 350186 135654
rect 350422 135418 350604 135654
rect 350004 135334 350604 135418
rect 350004 135098 350186 135334
rect 350422 135098 350604 135334
rect 350004 99654 350604 135098
rect 350004 99418 350186 99654
rect 350422 99418 350604 99654
rect 350004 99334 350604 99418
rect 350004 99098 350186 99334
rect 350422 99098 350604 99334
rect 350004 63654 350604 99098
rect 350004 63418 350186 63654
rect 350422 63418 350604 63654
rect 350004 63334 350604 63418
rect 350004 63098 350186 63334
rect 350422 63098 350604 63334
rect 350004 27654 350604 63098
rect 350004 27418 350186 27654
rect 350422 27418 350604 27654
rect 350004 27334 350604 27418
rect 350004 27098 350186 27334
rect 350422 27098 350604 27334
rect 350004 -5046 350604 27098
rect 350004 -5282 350186 -5046
rect 350422 -5282 350604 -5046
rect 350004 -5366 350604 -5282
rect 350004 -5602 350186 -5366
rect 350422 -5602 350604 -5366
rect 350004 -5624 350604 -5602
rect 353604 679254 354204 710862
rect 371604 710478 372204 711440
rect 371604 710242 371786 710478
rect 372022 710242 372204 710478
rect 371604 710158 372204 710242
rect 371604 709922 371786 710158
rect 372022 709922 372204 710158
rect 368004 708598 368604 709560
rect 368004 708362 368186 708598
rect 368422 708362 368604 708598
rect 368004 708278 368604 708362
rect 368004 708042 368186 708278
rect 368422 708042 368604 708278
rect 364404 706718 365004 707680
rect 364404 706482 364586 706718
rect 364822 706482 365004 706718
rect 364404 706398 365004 706482
rect 364404 706162 364586 706398
rect 364822 706162 365004 706398
rect 353604 679018 353786 679254
rect 354022 679018 354204 679254
rect 353604 678934 354204 679018
rect 353604 678698 353786 678934
rect 354022 678698 354204 678934
rect 353604 643254 354204 678698
rect 353604 643018 353786 643254
rect 354022 643018 354204 643254
rect 353604 642934 354204 643018
rect 353604 642698 353786 642934
rect 354022 642698 354204 642934
rect 353604 607254 354204 642698
rect 353604 607018 353786 607254
rect 354022 607018 354204 607254
rect 353604 606934 354204 607018
rect 353604 606698 353786 606934
rect 354022 606698 354204 606934
rect 353604 571254 354204 606698
rect 353604 571018 353786 571254
rect 354022 571018 354204 571254
rect 353604 570934 354204 571018
rect 353604 570698 353786 570934
rect 354022 570698 354204 570934
rect 353604 535254 354204 570698
rect 353604 535018 353786 535254
rect 354022 535018 354204 535254
rect 353604 534934 354204 535018
rect 353604 534698 353786 534934
rect 354022 534698 354204 534934
rect 353604 499254 354204 534698
rect 353604 499018 353786 499254
rect 354022 499018 354204 499254
rect 353604 498934 354204 499018
rect 353604 498698 353786 498934
rect 354022 498698 354204 498934
rect 353604 463254 354204 498698
rect 353604 463018 353786 463254
rect 354022 463018 354204 463254
rect 353604 462934 354204 463018
rect 353604 462698 353786 462934
rect 354022 462698 354204 462934
rect 353604 427254 354204 462698
rect 353604 427018 353786 427254
rect 354022 427018 354204 427254
rect 353604 426934 354204 427018
rect 353604 426698 353786 426934
rect 354022 426698 354204 426934
rect 353604 391254 354204 426698
rect 353604 391018 353786 391254
rect 354022 391018 354204 391254
rect 353604 390934 354204 391018
rect 353604 390698 353786 390934
rect 354022 390698 354204 390934
rect 353604 355254 354204 390698
rect 353604 355018 353786 355254
rect 354022 355018 354204 355254
rect 353604 354934 354204 355018
rect 353604 354698 353786 354934
rect 354022 354698 354204 354934
rect 353604 319254 354204 354698
rect 353604 319018 353786 319254
rect 354022 319018 354204 319254
rect 353604 318934 354204 319018
rect 353604 318698 353786 318934
rect 354022 318698 354204 318934
rect 353604 283254 354204 318698
rect 353604 283018 353786 283254
rect 354022 283018 354204 283254
rect 353604 282934 354204 283018
rect 353604 282698 353786 282934
rect 354022 282698 354204 282934
rect 353604 247254 354204 282698
rect 353604 247018 353786 247254
rect 354022 247018 354204 247254
rect 353604 246934 354204 247018
rect 353604 246698 353786 246934
rect 354022 246698 354204 246934
rect 353604 211254 354204 246698
rect 353604 211018 353786 211254
rect 354022 211018 354204 211254
rect 353604 210934 354204 211018
rect 353604 210698 353786 210934
rect 354022 210698 354204 210934
rect 353604 175254 354204 210698
rect 353604 175018 353786 175254
rect 354022 175018 354204 175254
rect 353604 174934 354204 175018
rect 353604 174698 353786 174934
rect 354022 174698 354204 174934
rect 353604 139254 354204 174698
rect 353604 139018 353786 139254
rect 354022 139018 354204 139254
rect 353604 138934 354204 139018
rect 353604 138698 353786 138934
rect 354022 138698 354204 138934
rect 353604 103254 354204 138698
rect 353604 103018 353786 103254
rect 354022 103018 354204 103254
rect 353604 102934 354204 103018
rect 353604 102698 353786 102934
rect 354022 102698 354204 102934
rect 353604 67254 354204 102698
rect 353604 67018 353786 67254
rect 354022 67018 354204 67254
rect 353604 66934 354204 67018
rect 353604 66698 353786 66934
rect 354022 66698 354204 66934
rect 353604 31254 354204 66698
rect 353604 31018 353786 31254
rect 354022 31018 354204 31254
rect 353604 30934 354204 31018
rect 353604 30698 353786 30934
rect 354022 30698 354204 30934
rect 335604 -6222 335786 -5986
rect 336022 -6222 336204 -5986
rect 335604 -6306 336204 -6222
rect 335604 -6542 335786 -6306
rect 336022 -6542 336204 -6306
rect 335604 -7504 336204 -6542
rect 353604 -6926 354204 30698
rect 360804 704838 361404 705800
rect 360804 704602 360986 704838
rect 361222 704602 361404 704838
rect 360804 704518 361404 704602
rect 360804 704282 360986 704518
rect 361222 704282 361404 704518
rect 360804 686454 361404 704282
rect 360804 686218 360986 686454
rect 361222 686218 361404 686454
rect 360804 686134 361404 686218
rect 360804 685898 360986 686134
rect 361222 685898 361404 686134
rect 360804 650454 361404 685898
rect 360804 650218 360986 650454
rect 361222 650218 361404 650454
rect 360804 650134 361404 650218
rect 360804 649898 360986 650134
rect 361222 649898 361404 650134
rect 360804 614454 361404 649898
rect 360804 614218 360986 614454
rect 361222 614218 361404 614454
rect 360804 614134 361404 614218
rect 360804 613898 360986 614134
rect 361222 613898 361404 614134
rect 360804 578454 361404 613898
rect 360804 578218 360986 578454
rect 361222 578218 361404 578454
rect 360804 578134 361404 578218
rect 360804 577898 360986 578134
rect 361222 577898 361404 578134
rect 360804 542454 361404 577898
rect 360804 542218 360986 542454
rect 361222 542218 361404 542454
rect 360804 542134 361404 542218
rect 360804 541898 360986 542134
rect 361222 541898 361404 542134
rect 360804 506454 361404 541898
rect 360804 506218 360986 506454
rect 361222 506218 361404 506454
rect 360804 506134 361404 506218
rect 360804 505898 360986 506134
rect 361222 505898 361404 506134
rect 360804 470454 361404 505898
rect 360804 470218 360986 470454
rect 361222 470218 361404 470454
rect 360804 470134 361404 470218
rect 360804 469898 360986 470134
rect 361222 469898 361404 470134
rect 360804 434454 361404 469898
rect 360804 434218 360986 434454
rect 361222 434218 361404 434454
rect 360804 434134 361404 434218
rect 360804 433898 360986 434134
rect 361222 433898 361404 434134
rect 360804 398454 361404 433898
rect 360804 398218 360986 398454
rect 361222 398218 361404 398454
rect 360804 398134 361404 398218
rect 360804 397898 360986 398134
rect 361222 397898 361404 398134
rect 360804 362454 361404 397898
rect 360804 362218 360986 362454
rect 361222 362218 361404 362454
rect 360804 362134 361404 362218
rect 360804 361898 360986 362134
rect 361222 361898 361404 362134
rect 360804 326454 361404 361898
rect 360804 326218 360986 326454
rect 361222 326218 361404 326454
rect 360804 326134 361404 326218
rect 360804 325898 360986 326134
rect 361222 325898 361404 326134
rect 360804 290454 361404 325898
rect 360804 290218 360986 290454
rect 361222 290218 361404 290454
rect 360804 290134 361404 290218
rect 360804 289898 360986 290134
rect 361222 289898 361404 290134
rect 360804 254454 361404 289898
rect 360804 254218 360986 254454
rect 361222 254218 361404 254454
rect 360804 254134 361404 254218
rect 360804 253898 360986 254134
rect 361222 253898 361404 254134
rect 360804 218454 361404 253898
rect 360804 218218 360986 218454
rect 361222 218218 361404 218454
rect 360804 218134 361404 218218
rect 360804 217898 360986 218134
rect 361222 217898 361404 218134
rect 360804 182454 361404 217898
rect 360804 182218 360986 182454
rect 361222 182218 361404 182454
rect 360804 182134 361404 182218
rect 360804 181898 360986 182134
rect 361222 181898 361404 182134
rect 360804 146454 361404 181898
rect 360804 146218 360986 146454
rect 361222 146218 361404 146454
rect 360804 146134 361404 146218
rect 360804 145898 360986 146134
rect 361222 145898 361404 146134
rect 360804 110454 361404 145898
rect 360804 110218 360986 110454
rect 361222 110218 361404 110454
rect 360804 110134 361404 110218
rect 360804 109898 360986 110134
rect 361222 109898 361404 110134
rect 360804 74454 361404 109898
rect 360804 74218 360986 74454
rect 361222 74218 361404 74454
rect 360804 74134 361404 74218
rect 360804 73898 360986 74134
rect 361222 73898 361404 74134
rect 360804 38454 361404 73898
rect 360804 38218 360986 38454
rect 361222 38218 361404 38454
rect 360804 38134 361404 38218
rect 360804 37898 360986 38134
rect 361222 37898 361404 38134
rect 360804 2454 361404 37898
rect 360804 2218 360986 2454
rect 361222 2218 361404 2454
rect 360804 2134 361404 2218
rect 360804 1898 360986 2134
rect 361222 1898 361404 2134
rect 360804 -346 361404 1898
rect 360804 -582 360986 -346
rect 361222 -582 361404 -346
rect 360804 -666 361404 -582
rect 360804 -902 360986 -666
rect 361222 -902 361404 -666
rect 360804 -1864 361404 -902
rect 364404 690054 365004 706162
rect 364404 689818 364586 690054
rect 364822 689818 365004 690054
rect 364404 689734 365004 689818
rect 364404 689498 364586 689734
rect 364822 689498 365004 689734
rect 364404 654054 365004 689498
rect 364404 653818 364586 654054
rect 364822 653818 365004 654054
rect 364404 653734 365004 653818
rect 364404 653498 364586 653734
rect 364822 653498 365004 653734
rect 364404 618054 365004 653498
rect 364404 617818 364586 618054
rect 364822 617818 365004 618054
rect 364404 617734 365004 617818
rect 364404 617498 364586 617734
rect 364822 617498 365004 617734
rect 364404 582054 365004 617498
rect 364404 581818 364586 582054
rect 364822 581818 365004 582054
rect 364404 581734 365004 581818
rect 364404 581498 364586 581734
rect 364822 581498 365004 581734
rect 364404 546054 365004 581498
rect 364404 545818 364586 546054
rect 364822 545818 365004 546054
rect 364404 545734 365004 545818
rect 364404 545498 364586 545734
rect 364822 545498 365004 545734
rect 364404 510054 365004 545498
rect 364404 509818 364586 510054
rect 364822 509818 365004 510054
rect 364404 509734 365004 509818
rect 364404 509498 364586 509734
rect 364822 509498 365004 509734
rect 364404 474054 365004 509498
rect 364404 473818 364586 474054
rect 364822 473818 365004 474054
rect 364404 473734 365004 473818
rect 364404 473498 364586 473734
rect 364822 473498 365004 473734
rect 364404 438054 365004 473498
rect 364404 437818 364586 438054
rect 364822 437818 365004 438054
rect 364404 437734 365004 437818
rect 364404 437498 364586 437734
rect 364822 437498 365004 437734
rect 364404 402054 365004 437498
rect 364404 401818 364586 402054
rect 364822 401818 365004 402054
rect 364404 401734 365004 401818
rect 364404 401498 364586 401734
rect 364822 401498 365004 401734
rect 364404 366054 365004 401498
rect 364404 365818 364586 366054
rect 364822 365818 365004 366054
rect 364404 365734 365004 365818
rect 364404 365498 364586 365734
rect 364822 365498 365004 365734
rect 364404 330054 365004 365498
rect 364404 329818 364586 330054
rect 364822 329818 365004 330054
rect 364404 329734 365004 329818
rect 364404 329498 364586 329734
rect 364822 329498 365004 329734
rect 364404 294054 365004 329498
rect 364404 293818 364586 294054
rect 364822 293818 365004 294054
rect 364404 293734 365004 293818
rect 364404 293498 364586 293734
rect 364822 293498 365004 293734
rect 364404 258054 365004 293498
rect 364404 257818 364586 258054
rect 364822 257818 365004 258054
rect 364404 257734 365004 257818
rect 364404 257498 364586 257734
rect 364822 257498 365004 257734
rect 364404 222054 365004 257498
rect 364404 221818 364586 222054
rect 364822 221818 365004 222054
rect 364404 221734 365004 221818
rect 364404 221498 364586 221734
rect 364822 221498 365004 221734
rect 364404 186054 365004 221498
rect 364404 185818 364586 186054
rect 364822 185818 365004 186054
rect 364404 185734 365004 185818
rect 364404 185498 364586 185734
rect 364822 185498 365004 185734
rect 364404 150054 365004 185498
rect 364404 149818 364586 150054
rect 364822 149818 365004 150054
rect 364404 149734 365004 149818
rect 364404 149498 364586 149734
rect 364822 149498 365004 149734
rect 364404 114054 365004 149498
rect 364404 113818 364586 114054
rect 364822 113818 365004 114054
rect 364404 113734 365004 113818
rect 364404 113498 364586 113734
rect 364822 113498 365004 113734
rect 364404 78054 365004 113498
rect 364404 77818 364586 78054
rect 364822 77818 365004 78054
rect 364404 77734 365004 77818
rect 364404 77498 364586 77734
rect 364822 77498 365004 77734
rect 364404 42054 365004 77498
rect 364404 41818 364586 42054
rect 364822 41818 365004 42054
rect 364404 41734 365004 41818
rect 364404 41498 364586 41734
rect 364822 41498 365004 41734
rect 364404 6054 365004 41498
rect 364404 5818 364586 6054
rect 364822 5818 365004 6054
rect 364404 5734 365004 5818
rect 364404 5498 364586 5734
rect 364822 5498 365004 5734
rect 364404 -2226 365004 5498
rect 364404 -2462 364586 -2226
rect 364822 -2462 365004 -2226
rect 364404 -2546 365004 -2462
rect 364404 -2782 364586 -2546
rect 364822 -2782 365004 -2546
rect 364404 -3744 365004 -2782
rect 368004 693654 368604 708042
rect 368004 693418 368186 693654
rect 368422 693418 368604 693654
rect 368004 693334 368604 693418
rect 368004 693098 368186 693334
rect 368422 693098 368604 693334
rect 368004 657654 368604 693098
rect 368004 657418 368186 657654
rect 368422 657418 368604 657654
rect 368004 657334 368604 657418
rect 368004 657098 368186 657334
rect 368422 657098 368604 657334
rect 368004 621654 368604 657098
rect 368004 621418 368186 621654
rect 368422 621418 368604 621654
rect 368004 621334 368604 621418
rect 368004 621098 368186 621334
rect 368422 621098 368604 621334
rect 368004 585654 368604 621098
rect 368004 585418 368186 585654
rect 368422 585418 368604 585654
rect 368004 585334 368604 585418
rect 368004 585098 368186 585334
rect 368422 585098 368604 585334
rect 368004 549654 368604 585098
rect 368004 549418 368186 549654
rect 368422 549418 368604 549654
rect 368004 549334 368604 549418
rect 368004 549098 368186 549334
rect 368422 549098 368604 549334
rect 368004 513654 368604 549098
rect 368004 513418 368186 513654
rect 368422 513418 368604 513654
rect 368004 513334 368604 513418
rect 368004 513098 368186 513334
rect 368422 513098 368604 513334
rect 368004 477654 368604 513098
rect 368004 477418 368186 477654
rect 368422 477418 368604 477654
rect 368004 477334 368604 477418
rect 368004 477098 368186 477334
rect 368422 477098 368604 477334
rect 368004 441654 368604 477098
rect 368004 441418 368186 441654
rect 368422 441418 368604 441654
rect 368004 441334 368604 441418
rect 368004 441098 368186 441334
rect 368422 441098 368604 441334
rect 368004 405654 368604 441098
rect 368004 405418 368186 405654
rect 368422 405418 368604 405654
rect 368004 405334 368604 405418
rect 368004 405098 368186 405334
rect 368422 405098 368604 405334
rect 368004 369654 368604 405098
rect 368004 369418 368186 369654
rect 368422 369418 368604 369654
rect 368004 369334 368604 369418
rect 368004 369098 368186 369334
rect 368422 369098 368604 369334
rect 368004 333654 368604 369098
rect 368004 333418 368186 333654
rect 368422 333418 368604 333654
rect 368004 333334 368604 333418
rect 368004 333098 368186 333334
rect 368422 333098 368604 333334
rect 368004 297654 368604 333098
rect 368004 297418 368186 297654
rect 368422 297418 368604 297654
rect 368004 297334 368604 297418
rect 368004 297098 368186 297334
rect 368422 297098 368604 297334
rect 368004 261654 368604 297098
rect 368004 261418 368186 261654
rect 368422 261418 368604 261654
rect 368004 261334 368604 261418
rect 368004 261098 368186 261334
rect 368422 261098 368604 261334
rect 368004 225654 368604 261098
rect 368004 225418 368186 225654
rect 368422 225418 368604 225654
rect 368004 225334 368604 225418
rect 368004 225098 368186 225334
rect 368422 225098 368604 225334
rect 368004 189654 368604 225098
rect 368004 189418 368186 189654
rect 368422 189418 368604 189654
rect 368004 189334 368604 189418
rect 368004 189098 368186 189334
rect 368422 189098 368604 189334
rect 368004 153654 368604 189098
rect 368004 153418 368186 153654
rect 368422 153418 368604 153654
rect 368004 153334 368604 153418
rect 368004 153098 368186 153334
rect 368422 153098 368604 153334
rect 368004 117654 368604 153098
rect 368004 117418 368186 117654
rect 368422 117418 368604 117654
rect 368004 117334 368604 117418
rect 368004 117098 368186 117334
rect 368422 117098 368604 117334
rect 368004 81654 368604 117098
rect 368004 81418 368186 81654
rect 368422 81418 368604 81654
rect 368004 81334 368604 81418
rect 368004 81098 368186 81334
rect 368422 81098 368604 81334
rect 368004 45654 368604 81098
rect 368004 45418 368186 45654
rect 368422 45418 368604 45654
rect 368004 45334 368604 45418
rect 368004 45098 368186 45334
rect 368422 45098 368604 45334
rect 368004 9654 368604 45098
rect 368004 9418 368186 9654
rect 368422 9418 368604 9654
rect 368004 9334 368604 9418
rect 368004 9098 368186 9334
rect 368422 9098 368604 9334
rect 368004 -4106 368604 9098
rect 368004 -4342 368186 -4106
rect 368422 -4342 368604 -4106
rect 368004 -4426 368604 -4342
rect 368004 -4662 368186 -4426
rect 368422 -4662 368604 -4426
rect 368004 -5624 368604 -4662
rect 371604 697254 372204 709922
rect 389604 711418 390204 711440
rect 389604 711182 389786 711418
rect 390022 711182 390204 711418
rect 389604 711098 390204 711182
rect 389604 710862 389786 711098
rect 390022 710862 390204 711098
rect 386004 709538 386604 709560
rect 386004 709302 386186 709538
rect 386422 709302 386604 709538
rect 386004 709218 386604 709302
rect 386004 708982 386186 709218
rect 386422 708982 386604 709218
rect 382404 707658 383004 707680
rect 382404 707422 382586 707658
rect 382822 707422 383004 707658
rect 382404 707338 383004 707422
rect 382404 707102 382586 707338
rect 382822 707102 383004 707338
rect 371604 697018 371786 697254
rect 372022 697018 372204 697254
rect 371604 696934 372204 697018
rect 371604 696698 371786 696934
rect 372022 696698 372204 696934
rect 371604 661254 372204 696698
rect 371604 661018 371786 661254
rect 372022 661018 372204 661254
rect 371604 660934 372204 661018
rect 371604 660698 371786 660934
rect 372022 660698 372204 660934
rect 371604 625254 372204 660698
rect 371604 625018 371786 625254
rect 372022 625018 372204 625254
rect 371604 624934 372204 625018
rect 371604 624698 371786 624934
rect 372022 624698 372204 624934
rect 371604 589254 372204 624698
rect 371604 589018 371786 589254
rect 372022 589018 372204 589254
rect 371604 588934 372204 589018
rect 371604 588698 371786 588934
rect 372022 588698 372204 588934
rect 371604 553254 372204 588698
rect 371604 553018 371786 553254
rect 372022 553018 372204 553254
rect 371604 552934 372204 553018
rect 371604 552698 371786 552934
rect 372022 552698 372204 552934
rect 371604 517254 372204 552698
rect 371604 517018 371786 517254
rect 372022 517018 372204 517254
rect 371604 516934 372204 517018
rect 371604 516698 371786 516934
rect 372022 516698 372204 516934
rect 371604 481254 372204 516698
rect 371604 481018 371786 481254
rect 372022 481018 372204 481254
rect 371604 480934 372204 481018
rect 371604 480698 371786 480934
rect 372022 480698 372204 480934
rect 371604 445254 372204 480698
rect 371604 445018 371786 445254
rect 372022 445018 372204 445254
rect 371604 444934 372204 445018
rect 371604 444698 371786 444934
rect 372022 444698 372204 444934
rect 371604 409254 372204 444698
rect 371604 409018 371786 409254
rect 372022 409018 372204 409254
rect 371604 408934 372204 409018
rect 371604 408698 371786 408934
rect 372022 408698 372204 408934
rect 371604 373254 372204 408698
rect 371604 373018 371786 373254
rect 372022 373018 372204 373254
rect 371604 372934 372204 373018
rect 371604 372698 371786 372934
rect 372022 372698 372204 372934
rect 371604 337254 372204 372698
rect 371604 337018 371786 337254
rect 372022 337018 372204 337254
rect 371604 336934 372204 337018
rect 371604 336698 371786 336934
rect 372022 336698 372204 336934
rect 371604 301254 372204 336698
rect 371604 301018 371786 301254
rect 372022 301018 372204 301254
rect 371604 300934 372204 301018
rect 371604 300698 371786 300934
rect 372022 300698 372204 300934
rect 371604 265254 372204 300698
rect 371604 265018 371786 265254
rect 372022 265018 372204 265254
rect 371604 264934 372204 265018
rect 371604 264698 371786 264934
rect 372022 264698 372204 264934
rect 371604 229254 372204 264698
rect 371604 229018 371786 229254
rect 372022 229018 372204 229254
rect 371604 228934 372204 229018
rect 371604 228698 371786 228934
rect 372022 228698 372204 228934
rect 371604 193254 372204 228698
rect 371604 193018 371786 193254
rect 372022 193018 372204 193254
rect 371604 192934 372204 193018
rect 371604 192698 371786 192934
rect 372022 192698 372204 192934
rect 371604 157254 372204 192698
rect 371604 157018 371786 157254
rect 372022 157018 372204 157254
rect 371604 156934 372204 157018
rect 371604 156698 371786 156934
rect 372022 156698 372204 156934
rect 371604 121254 372204 156698
rect 371604 121018 371786 121254
rect 372022 121018 372204 121254
rect 371604 120934 372204 121018
rect 371604 120698 371786 120934
rect 372022 120698 372204 120934
rect 371604 85254 372204 120698
rect 371604 85018 371786 85254
rect 372022 85018 372204 85254
rect 371604 84934 372204 85018
rect 371604 84698 371786 84934
rect 372022 84698 372204 84934
rect 371604 49254 372204 84698
rect 371604 49018 371786 49254
rect 372022 49018 372204 49254
rect 371604 48934 372204 49018
rect 371604 48698 371786 48934
rect 372022 48698 372204 48934
rect 371604 13254 372204 48698
rect 371604 13018 371786 13254
rect 372022 13018 372204 13254
rect 371604 12934 372204 13018
rect 371604 12698 371786 12934
rect 372022 12698 372204 12934
rect 353604 -7162 353786 -6926
rect 354022 -7162 354204 -6926
rect 353604 -7246 354204 -7162
rect 353604 -7482 353786 -7246
rect 354022 -7482 354204 -7246
rect 353604 -7504 354204 -7482
rect 371604 -5986 372204 12698
rect 378804 705778 379404 705800
rect 378804 705542 378986 705778
rect 379222 705542 379404 705778
rect 378804 705458 379404 705542
rect 378804 705222 378986 705458
rect 379222 705222 379404 705458
rect 378804 668454 379404 705222
rect 378804 668218 378986 668454
rect 379222 668218 379404 668454
rect 378804 668134 379404 668218
rect 378804 667898 378986 668134
rect 379222 667898 379404 668134
rect 378804 632454 379404 667898
rect 378804 632218 378986 632454
rect 379222 632218 379404 632454
rect 378804 632134 379404 632218
rect 378804 631898 378986 632134
rect 379222 631898 379404 632134
rect 378804 596454 379404 631898
rect 378804 596218 378986 596454
rect 379222 596218 379404 596454
rect 378804 596134 379404 596218
rect 378804 595898 378986 596134
rect 379222 595898 379404 596134
rect 378804 560454 379404 595898
rect 382404 672054 383004 707102
rect 382404 671818 382586 672054
rect 382822 671818 383004 672054
rect 382404 671734 383004 671818
rect 382404 671498 382586 671734
rect 382822 671498 383004 671734
rect 382404 636054 383004 671498
rect 382404 635818 382586 636054
rect 382822 635818 383004 636054
rect 382404 635734 383004 635818
rect 382404 635498 382586 635734
rect 382822 635498 383004 635734
rect 382404 600054 383004 635498
rect 382404 599818 382586 600054
rect 382822 599818 383004 600054
rect 382404 599734 383004 599818
rect 382404 599498 382586 599734
rect 382822 599498 383004 599734
rect 380019 572116 380085 572117
rect 380019 572052 380020 572116
rect 380084 572052 380085 572116
rect 380019 572051 380085 572052
rect 379467 563140 379533 563141
rect 379467 563076 379468 563140
rect 379532 563076 379533 563140
rect 379467 563075 379533 563076
rect 378804 560218 378986 560454
rect 379222 560218 379404 560454
rect 378804 560134 379404 560218
rect 378804 559898 378986 560134
rect 379222 559898 379404 560134
rect 378804 524454 379404 559898
rect 378804 524218 378986 524454
rect 379222 524218 379404 524454
rect 378804 524134 379404 524218
rect 378804 523898 378986 524134
rect 379222 523898 379404 524134
rect 378804 488454 379404 523898
rect 378804 488218 378986 488454
rect 379222 488218 379404 488454
rect 378804 488134 379404 488218
rect 378804 487898 378986 488134
rect 379222 487898 379404 488134
rect 378804 452454 379404 487898
rect 378804 452218 378986 452454
rect 379222 452218 379404 452454
rect 378804 452134 379404 452218
rect 378804 451898 378986 452134
rect 379222 451898 379404 452134
rect 378804 416454 379404 451898
rect 378804 416218 378986 416454
rect 379222 416218 379404 416454
rect 378804 416134 379404 416218
rect 378804 415898 378986 416134
rect 379222 415898 379404 416134
rect 378804 380454 379404 415898
rect 379470 394637 379530 563075
rect 379651 559604 379717 559605
rect 379651 559540 379652 559604
rect 379716 559540 379717 559604
rect 379651 559539 379717 559540
rect 379467 394636 379533 394637
rect 379467 394572 379468 394636
rect 379532 394572 379533 394636
rect 379467 394571 379533 394572
rect 379654 394501 379714 559539
rect 379835 528732 379901 528733
rect 379835 528668 379836 528732
rect 379900 528668 379901 528732
rect 379835 528667 379901 528668
rect 379838 417485 379898 528667
rect 380022 500173 380082 572051
rect 382404 564054 383004 599498
rect 382404 563818 382586 564054
rect 382822 563818 383004 564054
rect 382404 563734 383004 563818
rect 382404 563498 382586 563734
rect 382822 563498 383004 563734
rect 380203 541108 380269 541109
rect 380203 541044 380204 541108
rect 380268 541044 380269 541108
rect 380203 541043 380269 541044
rect 380206 500309 380266 541043
rect 382404 528054 383004 563498
rect 382404 527818 382586 528054
rect 382822 527818 383004 528054
rect 382404 527734 383004 527818
rect 382404 527498 382586 527734
rect 382822 527498 383004 527734
rect 380203 500308 380269 500309
rect 380203 500244 380204 500308
rect 380268 500244 380269 500308
rect 380203 500243 380269 500244
rect 380019 500172 380085 500173
rect 380019 500108 380020 500172
rect 380084 500108 380085 500172
rect 380019 500107 380085 500108
rect 382404 492054 383004 527498
rect 382404 491818 382586 492054
rect 382822 491818 383004 492054
rect 382404 491734 383004 491818
rect 382404 491498 382586 491734
rect 382822 491498 383004 491734
rect 382404 456054 383004 491498
rect 382404 455818 382586 456054
rect 382822 455818 383004 456054
rect 382404 455734 383004 455818
rect 382404 455498 382586 455734
rect 382822 455498 383004 455734
rect 382404 420054 383004 455498
rect 382404 419818 382586 420054
rect 382822 419818 383004 420054
rect 382404 419734 383004 419818
rect 382404 419498 382586 419734
rect 382822 419498 383004 419734
rect 379835 417484 379901 417485
rect 379835 417420 379836 417484
rect 379900 417420 379901 417484
rect 379835 417419 379901 417420
rect 379651 394500 379717 394501
rect 379651 394436 379652 394500
rect 379716 394436 379717 394500
rect 379651 394435 379717 394436
rect 378804 380218 378986 380454
rect 379222 380218 379404 380454
rect 378804 380134 379404 380218
rect 378804 379898 378986 380134
rect 379222 379898 379404 380134
rect 378804 344454 379404 379898
rect 378804 344218 378986 344454
rect 379222 344218 379404 344454
rect 378804 344134 379404 344218
rect 378804 343898 378986 344134
rect 379222 343898 379404 344134
rect 378804 308454 379404 343898
rect 378804 308218 378986 308454
rect 379222 308218 379404 308454
rect 378804 308134 379404 308218
rect 378804 307898 378986 308134
rect 379222 307898 379404 308134
rect 378804 272454 379404 307898
rect 378804 272218 378986 272454
rect 379222 272218 379404 272454
rect 378804 272134 379404 272218
rect 378804 271898 378986 272134
rect 379222 271898 379404 272134
rect 378804 236454 379404 271898
rect 378804 236218 378986 236454
rect 379222 236218 379404 236454
rect 378804 236134 379404 236218
rect 378804 235898 378986 236134
rect 379222 235898 379404 236134
rect 378804 200454 379404 235898
rect 378804 200218 378986 200454
rect 379222 200218 379404 200454
rect 378804 200134 379404 200218
rect 378804 199898 378986 200134
rect 379222 199898 379404 200134
rect 378804 164454 379404 199898
rect 378804 164218 378986 164454
rect 379222 164218 379404 164454
rect 378804 164134 379404 164218
rect 378804 163898 378986 164134
rect 379222 163898 379404 164134
rect 378804 128454 379404 163898
rect 378804 128218 378986 128454
rect 379222 128218 379404 128454
rect 378804 128134 379404 128218
rect 378804 127898 378986 128134
rect 379222 127898 379404 128134
rect 378804 92454 379404 127898
rect 378804 92218 378986 92454
rect 379222 92218 379404 92454
rect 378804 92134 379404 92218
rect 378804 91898 378986 92134
rect 379222 91898 379404 92134
rect 378804 56454 379404 91898
rect 378804 56218 378986 56454
rect 379222 56218 379404 56454
rect 378804 56134 379404 56218
rect 378804 55898 378986 56134
rect 379222 55898 379404 56134
rect 378804 20454 379404 55898
rect 378804 20218 378986 20454
rect 379222 20218 379404 20454
rect 378804 20134 379404 20218
rect 378804 19898 378986 20134
rect 379222 19898 379404 20134
rect 378804 -1286 379404 19898
rect 378804 -1522 378986 -1286
rect 379222 -1522 379404 -1286
rect 378804 -1606 379404 -1522
rect 378804 -1842 378986 -1606
rect 379222 -1842 379404 -1606
rect 378804 -1864 379404 -1842
rect 382404 384054 383004 419498
rect 382404 383818 382586 384054
rect 382822 383818 383004 384054
rect 382404 383734 383004 383818
rect 382404 383498 382586 383734
rect 382822 383498 383004 383734
rect 382404 348054 383004 383498
rect 382404 347818 382586 348054
rect 382822 347818 383004 348054
rect 382404 347734 383004 347818
rect 382404 347498 382586 347734
rect 382822 347498 383004 347734
rect 382404 312054 383004 347498
rect 382404 311818 382586 312054
rect 382822 311818 383004 312054
rect 382404 311734 383004 311818
rect 382404 311498 382586 311734
rect 382822 311498 383004 311734
rect 382404 276054 383004 311498
rect 382404 275818 382586 276054
rect 382822 275818 383004 276054
rect 382404 275734 383004 275818
rect 382404 275498 382586 275734
rect 382822 275498 383004 275734
rect 382404 240054 383004 275498
rect 382404 239818 382586 240054
rect 382822 239818 383004 240054
rect 382404 239734 383004 239818
rect 382404 239498 382586 239734
rect 382822 239498 383004 239734
rect 382404 204054 383004 239498
rect 382404 203818 382586 204054
rect 382822 203818 383004 204054
rect 382404 203734 383004 203818
rect 382404 203498 382586 203734
rect 382822 203498 383004 203734
rect 382404 168054 383004 203498
rect 382404 167818 382586 168054
rect 382822 167818 383004 168054
rect 382404 167734 383004 167818
rect 382404 167498 382586 167734
rect 382822 167498 383004 167734
rect 382404 132054 383004 167498
rect 382404 131818 382586 132054
rect 382822 131818 383004 132054
rect 382404 131734 383004 131818
rect 382404 131498 382586 131734
rect 382822 131498 383004 131734
rect 382404 96054 383004 131498
rect 382404 95818 382586 96054
rect 382822 95818 383004 96054
rect 382404 95734 383004 95818
rect 382404 95498 382586 95734
rect 382822 95498 383004 95734
rect 382404 60054 383004 95498
rect 382404 59818 382586 60054
rect 382822 59818 383004 60054
rect 382404 59734 383004 59818
rect 382404 59498 382586 59734
rect 382822 59498 383004 59734
rect 382404 24054 383004 59498
rect 382404 23818 382586 24054
rect 382822 23818 383004 24054
rect 382404 23734 383004 23818
rect 382404 23498 382586 23734
rect 382822 23498 383004 23734
rect 382404 -3166 383004 23498
rect 382404 -3402 382586 -3166
rect 382822 -3402 383004 -3166
rect 382404 -3486 383004 -3402
rect 382404 -3722 382586 -3486
rect 382822 -3722 383004 -3486
rect 382404 -3744 383004 -3722
rect 386004 675654 386604 708982
rect 386004 675418 386186 675654
rect 386422 675418 386604 675654
rect 386004 675334 386604 675418
rect 386004 675098 386186 675334
rect 386422 675098 386604 675334
rect 386004 639654 386604 675098
rect 386004 639418 386186 639654
rect 386422 639418 386604 639654
rect 386004 639334 386604 639418
rect 386004 639098 386186 639334
rect 386422 639098 386604 639334
rect 386004 603654 386604 639098
rect 386004 603418 386186 603654
rect 386422 603418 386604 603654
rect 386004 603334 386604 603418
rect 386004 603098 386186 603334
rect 386422 603098 386604 603334
rect 386004 567654 386604 603098
rect 386004 567418 386186 567654
rect 386422 567418 386604 567654
rect 386004 567334 386604 567418
rect 386004 567098 386186 567334
rect 386422 567098 386604 567334
rect 386004 531654 386604 567098
rect 386004 531418 386186 531654
rect 386422 531418 386604 531654
rect 386004 531334 386604 531418
rect 386004 531098 386186 531334
rect 386422 531098 386604 531334
rect 386004 495654 386604 531098
rect 386004 495418 386186 495654
rect 386422 495418 386604 495654
rect 386004 495334 386604 495418
rect 386004 495098 386186 495334
rect 386422 495098 386604 495334
rect 386004 459654 386604 495098
rect 386004 459418 386186 459654
rect 386422 459418 386604 459654
rect 386004 459334 386604 459418
rect 386004 459098 386186 459334
rect 386422 459098 386604 459334
rect 386004 423654 386604 459098
rect 386004 423418 386186 423654
rect 386422 423418 386604 423654
rect 386004 423334 386604 423418
rect 386004 423098 386186 423334
rect 386422 423098 386604 423334
rect 386004 387654 386604 423098
rect 386004 387418 386186 387654
rect 386422 387418 386604 387654
rect 386004 387334 386604 387418
rect 386004 387098 386186 387334
rect 386422 387098 386604 387334
rect 386004 351654 386604 387098
rect 386004 351418 386186 351654
rect 386422 351418 386604 351654
rect 386004 351334 386604 351418
rect 386004 351098 386186 351334
rect 386422 351098 386604 351334
rect 386004 315654 386604 351098
rect 386004 315418 386186 315654
rect 386422 315418 386604 315654
rect 386004 315334 386604 315418
rect 386004 315098 386186 315334
rect 386422 315098 386604 315334
rect 386004 279654 386604 315098
rect 386004 279418 386186 279654
rect 386422 279418 386604 279654
rect 386004 279334 386604 279418
rect 386004 279098 386186 279334
rect 386422 279098 386604 279334
rect 386004 243654 386604 279098
rect 386004 243418 386186 243654
rect 386422 243418 386604 243654
rect 386004 243334 386604 243418
rect 386004 243098 386186 243334
rect 386422 243098 386604 243334
rect 386004 207654 386604 243098
rect 386004 207418 386186 207654
rect 386422 207418 386604 207654
rect 386004 207334 386604 207418
rect 386004 207098 386186 207334
rect 386422 207098 386604 207334
rect 386004 171654 386604 207098
rect 386004 171418 386186 171654
rect 386422 171418 386604 171654
rect 386004 171334 386604 171418
rect 386004 171098 386186 171334
rect 386422 171098 386604 171334
rect 386004 135654 386604 171098
rect 386004 135418 386186 135654
rect 386422 135418 386604 135654
rect 386004 135334 386604 135418
rect 386004 135098 386186 135334
rect 386422 135098 386604 135334
rect 386004 99654 386604 135098
rect 386004 99418 386186 99654
rect 386422 99418 386604 99654
rect 386004 99334 386604 99418
rect 386004 99098 386186 99334
rect 386422 99098 386604 99334
rect 386004 63654 386604 99098
rect 386004 63418 386186 63654
rect 386422 63418 386604 63654
rect 386004 63334 386604 63418
rect 386004 63098 386186 63334
rect 386422 63098 386604 63334
rect 386004 27654 386604 63098
rect 386004 27418 386186 27654
rect 386422 27418 386604 27654
rect 386004 27334 386604 27418
rect 386004 27098 386186 27334
rect 386422 27098 386604 27334
rect 386004 -5046 386604 27098
rect 386004 -5282 386186 -5046
rect 386422 -5282 386604 -5046
rect 386004 -5366 386604 -5282
rect 386004 -5602 386186 -5366
rect 386422 -5602 386604 -5366
rect 386004 -5624 386604 -5602
rect 389604 679254 390204 710862
rect 407604 710478 408204 711440
rect 407604 710242 407786 710478
rect 408022 710242 408204 710478
rect 407604 710158 408204 710242
rect 407604 709922 407786 710158
rect 408022 709922 408204 710158
rect 404004 708598 404604 709560
rect 404004 708362 404186 708598
rect 404422 708362 404604 708598
rect 404004 708278 404604 708362
rect 404004 708042 404186 708278
rect 404422 708042 404604 708278
rect 400404 706718 401004 707680
rect 400404 706482 400586 706718
rect 400822 706482 401004 706718
rect 400404 706398 401004 706482
rect 400404 706162 400586 706398
rect 400822 706162 401004 706398
rect 389604 679018 389786 679254
rect 390022 679018 390204 679254
rect 389604 678934 390204 679018
rect 389604 678698 389786 678934
rect 390022 678698 390204 678934
rect 389604 643254 390204 678698
rect 389604 643018 389786 643254
rect 390022 643018 390204 643254
rect 389604 642934 390204 643018
rect 389604 642698 389786 642934
rect 390022 642698 390204 642934
rect 389604 607254 390204 642698
rect 389604 607018 389786 607254
rect 390022 607018 390204 607254
rect 389604 606934 390204 607018
rect 389604 606698 389786 606934
rect 390022 606698 390204 606934
rect 389604 571254 390204 606698
rect 389604 571018 389786 571254
rect 390022 571018 390204 571254
rect 389604 570934 390204 571018
rect 389604 570698 389786 570934
rect 390022 570698 390204 570934
rect 389604 535254 390204 570698
rect 389604 535018 389786 535254
rect 390022 535018 390204 535254
rect 389604 534934 390204 535018
rect 389604 534698 389786 534934
rect 390022 534698 390204 534934
rect 389604 499254 390204 534698
rect 389604 499018 389786 499254
rect 390022 499018 390204 499254
rect 389604 498934 390204 499018
rect 389604 498698 389786 498934
rect 390022 498698 390204 498934
rect 389604 463254 390204 498698
rect 389604 463018 389786 463254
rect 390022 463018 390204 463254
rect 389604 462934 390204 463018
rect 389604 462698 389786 462934
rect 390022 462698 390204 462934
rect 389604 427254 390204 462698
rect 389604 427018 389786 427254
rect 390022 427018 390204 427254
rect 389604 426934 390204 427018
rect 389604 426698 389786 426934
rect 390022 426698 390204 426934
rect 389604 391254 390204 426698
rect 389604 391018 389786 391254
rect 390022 391018 390204 391254
rect 389604 390934 390204 391018
rect 389604 390698 389786 390934
rect 390022 390698 390204 390934
rect 389604 355254 390204 390698
rect 389604 355018 389786 355254
rect 390022 355018 390204 355254
rect 389604 354934 390204 355018
rect 389604 354698 389786 354934
rect 390022 354698 390204 354934
rect 389604 319254 390204 354698
rect 389604 319018 389786 319254
rect 390022 319018 390204 319254
rect 389604 318934 390204 319018
rect 389604 318698 389786 318934
rect 390022 318698 390204 318934
rect 396804 704838 397404 705800
rect 396804 704602 396986 704838
rect 397222 704602 397404 704838
rect 396804 704518 397404 704602
rect 396804 704282 396986 704518
rect 397222 704282 397404 704518
rect 396804 686454 397404 704282
rect 396804 686218 396986 686454
rect 397222 686218 397404 686454
rect 396804 686134 397404 686218
rect 396804 685898 396986 686134
rect 397222 685898 397404 686134
rect 396804 650454 397404 685898
rect 396804 650218 396986 650454
rect 397222 650218 397404 650454
rect 396804 650134 397404 650218
rect 396804 649898 396986 650134
rect 397222 649898 397404 650134
rect 396804 614454 397404 649898
rect 396804 614218 396986 614454
rect 397222 614218 397404 614454
rect 396804 614134 397404 614218
rect 396804 613898 396986 614134
rect 397222 613898 397404 614134
rect 396804 578454 397404 613898
rect 396804 578218 396986 578454
rect 397222 578218 397404 578454
rect 396804 578134 397404 578218
rect 396804 577898 396986 578134
rect 397222 577898 397404 578134
rect 396804 542454 397404 577898
rect 396804 542218 396986 542454
rect 397222 542218 397404 542454
rect 396804 542134 397404 542218
rect 396804 541898 396986 542134
rect 397222 541898 397404 542134
rect 396804 506454 397404 541898
rect 396804 506218 396986 506454
rect 397222 506218 397404 506454
rect 396804 506134 397404 506218
rect 396804 505898 396986 506134
rect 397222 505898 397404 506134
rect 396804 470454 397404 505898
rect 396804 470218 396986 470454
rect 397222 470218 397404 470454
rect 396804 470134 397404 470218
rect 396804 469898 396986 470134
rect 397222 469898 397404 470134
rect 396804 434454 397404 469898
rect 396804 434218 396986 434454
rect 397222 434218 397404 434454
rect 396804 434134 397404 434218
rect 396804 433898 396986 434134
rect 397222 433898 397404 434134
rect 396804 398454 397404 433898
rect 396804 398218 396986 398454
rect 397222 398218 397404 398454
rect 396804 398134 397404 398218
rect 396804 397898 396986 398134
rect 397222 397898 397404 398134
rect 396804 362454 397404 397898
rect 396804 362218 396986 362454
rect 397222 362218 397404 362454
rect 396804 362134 397404 362218
rect 396804 361898 396986 362134
rect 397222 361898 397404 362134
rect 396804 326454 397404 361898
rect 396804 326218 396986 326454
rect 397222 326218 397404 326454
rect 396804 326134 397404 326218
rect 396804 325898 396986 326134
rect 397222 325898 397404 326134
rect 389604 283254 390204 318698
rect 391059 318748 391125 318749
rect 391059 318684 391060 318748
rect 391124 318684 391125 318748
rect 391059 318683 391125 318684
rect 391062 309229 391122 318683
rect 391059 309228 391125 309229
rect 391059 309164 391060 309228
rect 391124 309164 391125 309228
rect 391059 309163 391125 309164
rect 391059 299436 391125 299437
rect 391059 299372 391060 299436
rect 391124 299372 391125 299436
rect 391059 299371 391125 299372
rect 391062 289917 391122 299371
rect 396804 290454 397404 325898
rect 396804 290218 396986 290454
rect 397222 290218 397404 290454
rect 396804 290134 397404 290218
rect 391059 289916 391125 289917
rect 391059 289852 391060 289916
rect 391124 289852 391125 289916
rect 391059 289851 391125 289852
rect 396804 289898 396986 290134
rect 397222 289898 397404 290134
rect 389604 283018 389786 283254
rect 390022 283018 390204 283254
rect 389604 282934 390204 283018
rect 389604 282698 389786 282934
rect 390022 282698 390204 282934
rect 389604 247254 390204 282698
rect 391059 280124 391125 280125
rect 391059 280060 391060 280124
rect 391124 280060 391125 280124
rect 391059 280059 391125 280060
rect 391062 270605 391122 280059
rect 391059 270604 391125 270605
rect 391059 270540 391060 270604
rect 391124 270540 391125 270604
rect 391059 270539 391125 270540
rect 389604 247018 389786 247254
rect 390022 247018 390204 247254
rect 389604 246934 390204 247018
rect 389604 246698 389786 246934
rect 390022 246698 390204 246934
rect 389604 211254 390204 246698
rect 389604 211018 389786 211254
rect 390022 211018 390204 211254
rect 389604 210934 390204 211018
rect 389604 210698 389786 210934
rect 390022 210698 390204 210934
rect 389604 175254 390204 210698
rect 389604 175018 389786 175254
rect 390022 175018 390204 175254
rect 389604 174934 390204 175018
rect 389604 174698 389786 174934
rect 390022 174698 390204 174934
rect 389604 139254 390204 174698
rect 389604 139018 389786 139254
rect 390022 139018 390204 139254
rect 389604 138934 390204 139018
rect 389604 138698 389786 138934
rect 390022 138698 390204 138934
rect 389604 103254 390204 138698
rect 389604 103018 389786 103254
rect 390022 103018 390204 103254
rect 389604 102934 390204 103018
rect 389604 102698 389786 102934
rect 390022 102698 390204 102934
rect 389604 67254 390204 102698
rect 389604 67018 389786 67254
rect 390022 67018 390204 67254
rect 389604 66934 390204 67018
rect 389604 66698 389786 66934
rect 390022 66698 390204 66934
rect 389604 31254 390204 66698
rect 389604 31018 389786 31254
rect 390022 31018 390204 31254
rect 389604 30934 390204 31018
rect 389604 30698 389786 30934
rect 390022 30698 390204 30934
rect 371604 -6222 371786 -5986
rect 372022 -6222 372204 -5986
rect 371604 -6306 372204 -6222
rect 371604 -6542 371786 -6306
rect 372022 -6542 372204 -6306
rect 371604 -7504 372204 -6542
rect 389604 -6926 390204 30698
rect 396804 254454 397404 289898
rect 396804 254218 396986 254454
rect 397222 254218 397404 254454
rect 396804 254134 397404 254218
rect 396804 253898 396986 254134
rect 397222 253898 397404 254134
rect 396804 218454 397404 253898
rect 396804 218218 396986 218454
rect 397222 218218 397404 218454
rect 396804 218134 397404 218218
rect 396804 217898 396986 218134
rect 397222 217898 397404 218134
rect 396804 182454 397404 217898
rect 396804 182218 396986 182454
rect 397222 182218 397404 182454
rect 396804 182134 397404 182218
rect 396804 181898 396986 182134
rect 397222 181898 397404 182134
rect 396804 146454 397404 181898
rect 396804 146218 396986 146454
rect 397222 146218 397404 146454
rect 396804 146134 397404 146218
rect 396804 145898 396986 146134
rect 397222 145898 397404 146134
rect 396804 110454 397404 145898
rect 396804 110218 396986 110454
rect 397222 110218 397404 110454
rect 396804 110134 397404 110218
rect 396804 109898 396986 110134
rect 397222 109898 397404 110134
rect 396804 74454 397404 109898
rect 396804 74218 396986 74454
rect 397222 74218 397404 74454
rect 396804 74134 397404 74218
rect 396804 73898 396986 74134
rect 397222 73898 397404 74134
rect 396804 38454 397404 73898
rect 396804 38218 396986 38454
rect 397222 38218 397404 38454
rect 396804 38134 397404 38218
rect 396804 37898 396986 38134
rect 397222 37898 397404 38134
rect 396804 2454 397404 37898
rect 396804 2218 396986 2454
rect 397222 2218 397404 2454
rect 396804 2134 397404 2218
rect 396804 1898 396986 2134
rect 397222 1898 397404 2134
rect 396804 -346 397404 1898
rect 396804 -582 396986 -346
rect 397222 -582 397404 -346
rect 396804 -666 397404 -582
rect 396804 -902 396986 -666
rect 397222 -902 397404 -666
rect 396804 -1864 397404 -902
rect 400404 690054 401004 706162
rect 400404 689818 400586 690054
rect 400822 689818 401004 690054
rect 400404 689734 401004 689818
rect 400404 689498 400586 689734
rect 400822 689498 401004 689734
rect 400404 654054 401004 689498
rect 400404 653818 400586 654054
rect 400822 653818 401004 654054
rect 400404 653734 401004 653818
rect 400404 653498 400586 653734
rect 400822 653498 401004 653734
rect 400404 618054 401004 653498
rect 400404 617818 400586 618054
rect 400822 617818 401004 618054
rect 400404 617734 401004 617818
rect 400404 617498 400586 617734
rect 400822 617498 401004 617734
rect 400404 582054 401004 617498
rect 400404 581818 400586 582054
rect 400822 581818 401004 582054
rect 400404 581734 401004 581818
rect 400404 581498 400586 581734
rect 400822 581498 401004 581734
rect 400404 546054 401004 581498
rect 400404 545818 400586 546054
rect 400822 545818 401004 546054
rect 400404 545734 401004 545818
rect 400404 545498 400586 545734
rect 400822 545498 401004 545734
rect 400404 510054 401004 545498
rect 400404 509818 400586 510054
rect 400822 509818 401004 510054
rect 400404 509734 401004 509818
rect 400404 509498 400586 509734
rect 400822 509498 401004 509734
rect 400404 474054 401004 509498
rect 400404 473818 400586 474054
rect 400822 473818 401004 474054
rect 400404 473734 401004 473818
rect 400404 473498 400586 473734
rect 400822 473498 401004 473734
rect 400404 438054 401004 473498
rect 400404 437818 400586 438054
rect 400822 437818 401004 438054
rect 400404 437734 401004 437818
rect 400404 437498 400586 437734
rect 400822 437498 401004 437734
rect 400404 402054 401004 437498
rect 400404 401818 400586 402054
rect 400822 401818 401004 402054
rect 400404 401734 401004 401818
rect 400404 401498 400586 401734
rect 400822 401498 401004 401734
rect 400404 366054 401004 401498
rect 400404 365818 400586 366054
rect 400822 365818 401004 366054
rect 400404 365734 401004 365818
rect 400404 365498 400586 365734
rect 400822 365498 401004 365734
rect 400404 330054 401004 365498
rect 400404 329818 400586 330054
rect 400822 329818 401004 330054
rect 400404 329734 401004 329818
rect 400404 329498 400586 329734
rect 400822 329498 401004 329734
rect 400404 294054 401004 329498
rect 400404 293818 400586 294054
rect 400822 293818 401004 294054
rect 400404 293734 401004 293818
rect 400404 293498 400586 293734
rect 400822 293498 401004 293734
rect 400404 258054 401004 293498
rect 400404 257818 400586 258054
rect 400822 257818 401004 258054
rect 400404 257734 401004 257818
rect 400404 257498 400586 257734
rect 400822 257498 401004 257734
rect 400404 222054 401004 257498
rect 400404 221818 400586 222054
rect 400822 221818 401004 222054
rect 400404 221734 401004 221818
rect 400404 221498 400586 221734
rect 400822 221498 401004 221734
rect 400404 186054 401004 221498
rect 400404 185818 400586 186054
rect 400822 185818 401004 186054
rect 400404 185734 401004 185818
rect 400404 185498 400586 185734
rect 400822 185498 401004 185734
rect 400404 150054 401004 185498
rect 400404 149818 400586 150054
rect 400822 149818 401004 150054
rect 400404 149734 401004 149818
rect 400404 149498 400586 149734
rect 400822 149498 401004 149734
rect 400404 114054 401004 149498
rect 400404 113818 400586 114054
rect 400822 113818 401004 114054
rect 400404 113734 401004 113818
rect 400404 113498 400586 113734
rect 400822 113498 401004 113734
rect 400404 78054 401004 113498
rect 400404 77818 400586 78054
rect 400822 77818 401004 78054
rect 400404 77734 401004 77818
rect 400404 77498 400586 77734
rect 400822 77498 401004 77734
rect 400404 42054 401004 77498
rect 400404 41818 400586 42054
rect 400822 41818 401004 42054
rect 400404 41734 401004 41818
rect 400404 41498 400586 41734
rect 400822 41498 401004 41734
rect 400404 6054 401004 41498
rect 400404 5818 400586 6054
rect 400822 5818 401004 6054
rect 400404 5734 401004 5818
rect 400404 5498 400586 5734
rect 400822 5498 401004 5734
rect 400404 -2226 401004 5498
rect 400404 -2462 400586 -2226
rect 400822 -2462 401004 -2226
rect 400404 -2546 401004 -2462
rect 400404 -2782 400586 -2546
rect 400822 -2782 401004 -2546
rect 400404 -3744 401004 -2782
rect 404004 693654 404604 708042
rect 404004 693418 404186 693654
rect 404422 693418 404604 693654
rect 404004 693334 404604 693418
rect 404004 693098 404186 693334
rect 404422 693098 404604 693334
rect 404004 657654 404604 693098
rect 404004 657418 404186 657654
rect 404422 657418 404604 657654
rect 404004 657334 404604 657418
rect 404004 657098 404186 657334
rect 404422 657098 404604 657334
rect 404004 621654 404604 657098
rect 404004 621418 404186 621654
rect 404422 621418 404604 621654
rect 404004 621334 404604 621418
rect 404004 621098 404186 621334
rect 404422 621098 404604 621334
rect 404004 585654 404604 621098
rect 404004 585418 404186 585654
rect 404422 585418 404604 585654
rect 404004 585334 404604 585418
rect 404004 585098 404186 585334
rect 404422 585098 404604 585334
rect 404004 549654 404604 585098
rect 404004 549418 404186 549654
rect 404422 549418 404604 549654
rect 404004 549334 404604 549418
rect 404004 549098 404186 549334
rect 404422 549098 404604 549334
rect 404004 513654 404604 549098
rect 404004 513418 404186 513654
rect 404422 513418 404604 513654
rect 404004 513334 404604 513418
rect 404004 513098 404186 513334
rect 404422 513098 404604 513334
rect 404004 477654 404604 513098
rect 404004 477418 404186 477654
rect 404422 477418 404604 477654
rect 404004 477334 404604 477418
rect 404004 477098 404186 477334
rect 404422 477098 404604 477334
rect 404004 441654 404604 477098
rect 404004 441418 404186 441654
rect 404422 441418 404604 441654
rect 404004 441334 404604 441418
rect 404004 441098 404186 441334
rect 404422 441098 404604 441334
rect 404004 405654 404604 441098
rect 404004 405418 404186 405654
rect 404422 405418 404604 405654
rect 404004 405334 404604 405418
rect 404004 405098 404186 405334
rect 404422 405098 404604 405334
rect 404004 369654 404604 405098
rect 404004 369418 404186 369654
rect 404422 369418 404604 369654
rect 404004 369334 404604 369418
rect 404004 369098 404186 369334
rect 404422 369098 404604 369334
rect 404004 333654 404604 369098
rect 404004 333418 404186 333654
rect 404422 333418 404604 333654
rect 404004 333334 404604 333418
rect 404004 333098 404186 333334
rect 404422 333098 404604 333334
rect 404004 297654 404604 333098
rect 404004 297418 404186 297654
rect 404422 297418 404604 297654
rect 404004 297334 404604 297418
rect 404004 297098 404186 297334
rect 404422 297098 404604 297334
rect 404004 261654 404604 297098
rect 404004 261418 404186 261654
rect 404422 261418 404604 261654
rect 404004 261334 404604 261418
rect 404004 261098 404186 261334
rect 404422 261098 404604 261334
rect 404004 225654 404604 261098
rect 404004 225418 404186 225654
rect 404422 225418 404604 225654
rect 404004 225334 404604 225418
rect 404004 225098 404186 225334
rect 404422 225098 404604 225334
rect 404004 189654 404604 225098
rect 404004 189418 404186 189654
rect 404422 189418 404604 189654
rect 404004 189334 404604 189418
rect 404004 189098 404186 189334
rect 404422 189098 404604 189334
rect 404004 153654 404604 189098
rect 404004 153418 404186 153654
rect 404422 153418 404604 153654
rect 404004 153334 404604 153418
rect 404004 153098 404186 153334
rect 404422 153098 404604 153334
rect 404004 117654 404604 153098
rect 404004 117418 404186 117654
rect 404422 117418 404604 117654
rect 404004 117334 404604 117418
rect 404004 117098 404186 117334
rect 404422 117098 404604 117334
rect 404004 81654 404604 117098
rect 404004 81418 404186 81654
rect 404422 81418 404604 81654
rect 404004 81334 404604 81418
rect 404004 81098 404186 81334
rect 404422 81098 404604 81334
rect 404004 45654 404604 81098
rect 404004 45418 404186 45654
rect 404422 45418 404604 45654
rect 404004 45334 404604 45418
rect 404004 45098 404186 45334
rect 404422 45098 404604 45334
rect 404004 9654 404604 45098
rect 404004 9418 404186 9654
rect 404422 9418 404604 9654
rect 404004 9334 404604 9418
rect 404004 9098 404186 9334
rect 404422 9098 404604 9334
rect 404004 -4106 404604 9098
rect 404004 -4342 404186 -4106
rect 404422 -4342 404604 -4106
rect 404004 -4426 404604 -4342
rect 404004 -4662 404186 -4426
rect 404422 -4662 404604 -4426
rect 404004 -5624 404604 -4662
rect 407604 697254 408204 709922
rect 425604 711418 426204 711440
rect 425604 711182 425786 711418
rect 426022 711182 426204 711418
rect 425604 711098 426204 711182
rect 425604 710862 425786 711098
rect 426022 710862 426204 711098
rect 422004 709538 422604 709560
rect 422004 709302 422186 709538
rect 422422 709302 422604 709538
rect 422004 709218 422604 709302
rect 422004 708982 422186 709218
rect 422422 708982 422604 709218
rect 418404 707658 419004 707680
rect 418404 707422 418586 707658
rect 418822 707422 419004 707658
rect 418404 707338 419004 707422
rect 418404 707102 418586 707338
rect 418822 707102 419004 707338
rect 407604 697018 407786 697254
rect 408022 697018 408204 697254
rect 407604 696934 408204 697018
rect 407604 696698 407786 696934
rect 408022 696698 408204 696934
rect 407604 661254 408204 696698
rect 407604 661018 407786 661254
rect 408022 661018 408204 661254
rect 407604 660934 408204 661018
rect 407604 660698 407786 660934
rect 408022 660698 408204 660934
rect 407604 625254 408204 660698
rect 407604 625018 407786 625254
rect 408022 625018 408204 625254
rect 407604 624934 408204 625018
rect 407604 624698 407786 624934
rect 408022 624698 408204 624934
rect 407604 589254 408204 624698
rect 407604 589018 407786 589254
rect 408022 589018 408204 589254
rect 407604 588934 408204 589018
rect 407604 588698 407786 588934
rect 408022 588698 408204 588934
rect 407604 553254 408204 588698
rect 407604 553018 407786 553254
rect 408022 553018 408204 553254
rect 407604 552934 408204 553018
rect 407604 552698 407786 552934
rect 408022 552698 408204 552934
rect 407604 517254 408204 552698
rect 407604 517018 407786 517254
rect 408022 517018 408204 517254
rect 407604 516934 408204 517018
rect 407604 516698 407786 516934
rect 408022 516698 408204 516934
rect 407604 481254 408204 516698
rect 407604 481018 407786 481254
rect 408022 481018 408204 481254
rect 407604 480934 408204 481018
rect 407604 480698 407786 480934
rect 408022 480698 408204 480934
rect 407604 445254 408204 480698
rect 407604 445018 407786 445254
rect 408022 445018 408204 445254
rect 407604 444934 408204 445018
rect 407604 444698 407786 444934
rect 408022 444698 408204 444934
rect 407604 409254 408204 444698
rect 407604 409018 407786 409254
rect 408022 409018 408204 409254
rect 407604 408934 408204 409018
rect 407604 408698 407786 408934
rect 408022 408698 408204 408934
rect 407604 373254 408204 408698
rect 407604 373018 407786 373254
rect 408022 373018 408204 373254
rect 407604 372934 408204 373018
rect 407604 372698 407786 372934
rect 408022 372698 408204 372934
rect 407604 337254 408204 372698
rect 407604 337018 407786 337254
rect 408022 337018 408204 337254
rect 407604 336934 408204 337018
rect 407604 336698 407786 336934
rect 408022 336698 408204 336934
rect 407604 301254 408204 336698
rect 407604 301018 407786 301254
rect 408022 301018 408204 301254
rect 407604 300934 408204 301018
rect 407604 300698 407786 300934
rect 408022 300698 408204 300934
rect 407604 265254 408204 300698
rect 407604 265018 407786 265254
rect 408022 265018 408204 265254
rect 407604 264934 408204 265018
rect 407604 264698 407786 264934
rect 408022 264698 408204 264934
rect 407604 229254 408204 264698
rect 407604 229018 407786 229254
rect 408022 229018 408204 229254
rect 407604 228934 408204 229018
rect 407604 228698 407786 228934
rect 408022 228698 408204 228934
rect 407604 193254 408204 228698
rect 407604 193018 407786 193254
rect 408022 193018 408204 193254
rect 407604 192934 408204 193018
rect 407604 192698 407786 192934
rect 408022 192698 408204 192934
rect 407604 157254 408204 192698
rect 407604 157018 407786 157254
rect 408022 157018 408204 157254
rect 407604 156934 408204 157018
rect 407604 156698 407786 156934
rect 408022 156698 408204 156934
rect 407604 121254 408204 156698
rect 407604 121018 407786 121254
rect 408022 121018 408204 121254
rect 407604 120934 408204 121018
rect 407604 120698 407786 120934
rect 408022 120698 408204 120934
rect 407604 85254 408204 120698
rect 407604 85018 407786 85254
rect 408022 85018 408204 85254
rect 407604 84934 408204 85018
rect 407604 84698 407786 84934
rect 408022 84698 408204 84934
rect 407604 49254 408204 84698
rect 407604 49018 407786 49254
rect 408022 49018 408204 49254
rect 407604 48934 408204 49018
rect 407604 48698 407786 48934
rect 408022 48698 408204 48934
rect 407604 13254 408204 48698
rect 407604 13018 407786 13254
rect 408022 13018 408204 13254
rect 407604 12934 408204 13018
rect 407604 12698 407786 12934
rect 408022 12698 408204 12934
rect 389604 -7162 389786 -6926
rect 390022 -7162 390204 -6926
rect 389604 -7246 390204 -7162
rect 389604 -7482 389786 -7246
rect 390022 -7482 390204 -7246
rect 389604 -7504 390204 -7482
rect 407604 -5986 408204 12698
rect 414804 705778 415404 705800
rect 414804 705542 414986 705778
rect 415222 705542 415404 705778
rect 414804 705458 415404 705542
rect 414804 705222 414986 705458
rect 415222 705222 415404 705458
rect 414804 668454 415404 705222
rect 414804 668218 414986 668454
rect 415222 668218 415404 668454
rect 414804 668134 415404 668218
rect 414804 667898 414986 668134
rect 415222 667898 415404 668134
rect 414804 632454 415404 667898
rect 414804 632218 414986 632454
rect 415222 632218 415404 632454
rect 414804 632134 415404 632218
rect 414804 631898 414986 632134
rect 415222 631898 415404 632134
rect 414804 596454 415404 631898
rect 414804 596218 414986 596454
rect 415222 596218 415404 596454
rect 414804 596134 415404 596218
rect 414804 595898 414986 596134
rect 415222 595898 415404 596134
rect 414804 560454 415404 595898
rect 414804 560218 414986 560454
rect 415222 560218 415404 560454
rect 414804 560134 415404 560218
rect 414804 559898 414986 560134
rect 415222 559898 415404 560134
rect 414804 524454 415404 559898
rect 414804 524218 414986 524454
rect 415222 524218 415404 524454
rect 414804 524134 415404 524218
rect 414804 523898 414986 524134
rect 415222 523898 415404 524134
rect 414804 488454 415404 523898
rect 414804 488218 414986 488454
rect 415222 488218 415404 488454
rect 414804 488134 415404 488218
rect 414804 487898 414986 488134
rect 415222 487898 415404 488134
rect 414804 452454 415404 487898
rect 414804 452218 414986 452454
rect 415222 452218 415404 452454
rect 414804 452134 415404 452218
rect 414804 451898 414986 452134
rect 415222 451898 415404 452134
rect 414804 416454 415404 451898
rect 414804 416218 414986 416454
rect 415222 416218 415404 416454
rect 414804 416134 415404 416218
rect 414804 415898 414986 416134
rect 415222 415898 415404 416134
rect 414804 380454 415404 415898
rect 414804 380218 414986 380454
rect 415222 380218 415404 380454
rect 414804 380134 415404 380218
rect 414804 379898 414986 380134
rect 415222 379898 415404 380134
rect 414804 344454 415404 379898
rect 414804 344218 414986 344454
rect 415222 344218 415404 344454
rect 414804 344134 415404 344218
rect 414804 343898 414986 344134
rect 415222 343898 415404 344134
rect 414804 308454 415404 343898
rect 414804 308218 414986 308454
rect 415222 308218 415404 308454
rect 414804 308134 415404 308218
rect 414804 307898 414986 308134
rect 415222 307898 415404 308134
rect 414804 272454 415404 307898
rect 414804 272218 414986 272454
rect 415222 272218 415404 272454
rect 414804 272134 415404 272218
rect 414804 271898 414986 272134
rect 415222 271898 415404 272134
rect 414804 236454 415404 271898
rect 414804 236218 414986 236454
rect 415222 236218 415404 236454
rect 414804 236134 415404 236218
rect 414804 235898 414986 236134
rect 415222 235898 415404 236134
rect 414804 200454 415404 235898
rect 414804 200218 414986 200454
rect 415222 200218 415404 200454
rect 414804 200134 415404 200218
rect 414804 199898 414986 200134
rect 415222 199898 415404 200134
rect 414804 164454 415404 199898
rect 414804 164218 414986 164454
rect 415222 164218 415404 164454
rect 414804 164134 415404 164218
rect 414804 163898 414986 164134
rect 415222 163898 415404 164134
rect 414804 128454 415404 163898
rect 414804 128218 414986 128454
rect 415222 128218 415404 128454
rect 414804 128134 415404 128218
rect 414804 127898 414986 128134
rect 415222 127898 415404 128134
rect 414804 92454 415404 127898
rect 414804 92218 414986 92454
rect 415222 92218 415404 92454
rect 414804 92134 415404 92218
rect 414804 91898 414986 92134
rect 415222 91898 415404 92134
rect 414804 56454 415404 91898
rect 414804 56218 414986 56454
rect 415222 56218 415404 56454
rect 414804 56134 415404 56218
rect 414804 55898 414986 56134
rect 415222 55898 415404 56134
rect 414804 20454 415404 55898
rect 414804 20218 414986 20454
rect 415222 20218 415404 20454
rect 414804 20134 415404 20218
rect 414804 19898 414986 20134
rect 415222 19898 415404 20134
rect 414804 -1286 415404 19898
rect 414804 -1522 414986 -1286
rect 415222 -1522 415404 -1286
rect 414804 -1606 415404 -1522
rect 414804 -1842 414986 -1606
rect 415222 -1842 415404 -1606
rect 414804 -1864 415404 -1842
rect 418404 672054 419004 707102
rect 418404 671818 418586 672054
rect 418822 671818 419004 672054
rect 418404 671734 419004 671818
rect 418404 671498 418586 671734
rect 418822 671498 419004 671734
rect 418404 636054 419004 671498
rect 418404 635818 418586 636054
rect 418822 635818 419004 636054
rect 418404 635734 419004 635818
rect 418404 635498 418586 635734
rect 418822 635498 419004 635734
rect 418404 600054 419004 635498
rect 418404 599818 418586 600054
rect 418822 599818 419004 600054
rect 418404 599734 419004 599818
rect 418404 599498 418586 599734
rect 418822 599498 419004 599734
rect 418404 564054 419004 599498
rect 418404 563818 418586 564054
rect 418822 563818 419004 564054
rect 418404 563734 419004 563818
rect 418404 563498 418586 563734
rect 418822 563498 419004 563734
rect 418404 528054 419004 563498
rect 418404 527818 418586 528054
rect 418822 527818 419004 528054
rect 418404 527734 419004 527818
rect 418404 527498 418586 527734
rect 418822 527498 419004 527734
rect 418404 492054 419004 527498
rect 418404 491818 418586 492054
rect 418822 491818 419004 492054
rect 418404 491734 419004 491818
rect 418404 491498 418586 491734
rect 418822 491498 419004 491734
rect 418404 456054 419004 491498
rect 418404 455818 418586 456054
rect 418822 455818 419004 456054
rect 418404 455734 419004 455818
rect 418404 455498 418586 455734
rect 418822 455498 419004 455734
rect 418404 420054 419004 455498
rect 418404 419818 418586 420054
rect 418822 419818 419004 420054
rect 418404 419734 419004 419818
rect 418404 419498 418586 419734
rect 418822 419498 419004 419734
rect 418404 384054 419004 419498
rect 418404 383818 418586 384054
rect 418822 383818 419004 384054
rect 418404 383734 419004 383818
rect 418404 383498 418586 383734
rect 418822 383498 419004 383734
rect 418404 348054 419004 383498
rect 418404 347818 418586 348054
rect 418822 347818 419004 348054
rect 418404 347734 419004 347818
rect 418404 347498 418586 347734
rect 418822 347498 419004 347734
rect 418404 312054 419004 347498
rect 418404 311818 418586 312054
rect 418822 311818 419004 312054
rect 418404 311734 419004 311818
rect 418404 311498 418586 311734
rect 418822 311498 419004 311734
rect 418404 276054 419004 311498
rect 418404 275818 418586 276054
rect 418822 275818 419004 276054
rect 418404 275734 419004 275818
rect 418404 275498 418586 275734
rect 418822 275498 419004 275734
rect 418404 240054 419004 275498
rect 418404 239818 418586 240054
rect 418822 239818 419004 240054
rect 418404 239734 419004 239818
rect 418404 239498 418586 239734
rect 418822 239498 419004 239734
rect 418404 204054 419004 239498
rect 418404 203818 418586 204054
rect 418822 203818 419004 204054
rect 418404 203734 419004 203818
rect 418404 203498 418586 203734
rect 418822 203498 419004 203734
rect 418404 168054 419004 203498
rect 418404 167818 418586 168054
rect 418822 167818 419004 168054
rect 418404 167734 419004 167818
rect 418404 167498 418586 167734
rect 418822 167498 419004 167734
rect 418404 132054 419004 167498
rect 418404 131818 418586 132054
rect 418822 131818 419004 132054
rect 418404 131734 419004 131818
rect 418404 131498 418586 131734
rect 418822 131498 419004 131734
rect 418404 96054 419004 131498
rect 418404 95818 418586 96054
rect 418822 95818 419004 96054
rect 418404 95734 419004 95818
rect 418404 95498 418586 95734
rect 418822 95498 419004 95734
rect 418404 60054 419004 95498
rect 422004 675654 422604 708982
rect 422004 675418 422186 675654
rect 422422 675418 422604 675654
rect 422004 675334 422604 675418
rect 422004 675098 422186 675334
rect 422422 675098 422604 675334
rect 422004 639654 422604 675098
rect 422004 639418 422186 639654
rect 422422 639418 422604 639654
rect 422004 639334 422604 639418
rect 422004 639098 422186 639334
rect 422422 639098 422604 639334
rect 422004 603654 422604 639098
rect 422004 603418 422186 603654
rect 422422 603418 422604 603654
rect 422004 603334 422604 603418
rect 422004 603098 422186 603334
rect 422422 603098 422604 603334
rect 422004 567654 422604 603098
rect 422004 567418 422186 567654
rect 422422 567418 422604 567654
rect 422004 567334 422604 567418
rect 422004 567098 422186 567334
rect 422422 567098 422604 567334
rect 422004 531654 422604 567098
rect 422004 531418 422186 531654
rect 422422 531418 422604 531654
rect 422004 531334 422604 531418
rect 422004 531098 422186 531334
rect 422422 531098 422604 531334
rect 422004 495654 422604 531098
rect 422004 495418 422186 495654
rect 422422 495418 422604 495654
rect 422004 495334 422604 495418
rect 422004 495098 422186 495334
rect 422422 495098 422604 495334
rect 422004 459654 422604 495098
rect 422004 459418 422186 459654
rect 422422 459418 422604 459654
rect 422004 459334 422604 459418
rect 422004 459098 422186 459334
rect 422422 459098 422604 459334
rect 422004 423654 422604 459098
rect 422004 423418 422186 423654
rect 422422 423418 422604 423654
rect 422004 423334 422604 423418
rect 422004 423098 422186 423334
rect 422422 423098 422604 423334
rect 422004 387654 422604 423098
rect 422004 387418 422186 387654
rect 422422 387418 422604 387654
rect 422004 387334 422604 387418
rect 422004 387098 422186 387334
rect 422422 387098 422604 387334
rect 422004 351654 422604 387098
rect 422004 351418 422186 351654
rect 422422 351418 422604 351654
rect 422004 351334 422604 351418
rect 422004 351098 422186 351334
rect 422422 351098 422604 351334
rect 422004 315654 422604 351098
rect 422004 315418 422186 315654
rect 422422 315418 422604 315654
rect 422004 315334 422604 315418
rect 422004 315098 422186 315334
rect 422422 315098 422604 315334
rect 422004 279654 422604 315098
rect 422004 279418 422186 279654
rect 422422 279418 422604 279654
rect 422004 279334 422604 279418
rect 422004 279098 422186 279334
rect 422422 279098 422604 279334
rect 422004 243654 422604 279098
rect 422004 243418 422186 243654
rect 422422 243418 422604 243654
rect 422004 243334 422604 243418
rect 422004 243098 422186 243334
rect 422422 243098 422604 243334
rect 422004 207654 422604 243098
rect 422004 207418 422186 207654
rect 422422 207418 422604 207654
rect 422004 207334 422604 207418
rect 422004 207098 422186 207334
rect 422422 207098 422604 207334
rect 422004 171654 422604 207098
rect 422004 171418 422186 171654
rect 422422 171418 422604 171654
rect 422004 171334 422604 171418
rect 422004 171098 422186 171334
rect 422422 171098 422604 171334
rect 422004 135654 422604 171098
rect 422004 135418 422186 135654
rect 422422 135418 422604 135654
rect 422004 135334 422604 135418
rect 422004 135098 422186 135334
rect 422422 135098 422604 135334
rect 422004 99654 422604 135098
rect 422004 99418 422186 99654
rect 422422 99418 422604 99654
rect 422004 99334 422604 99418
rect 422004 99098 422186 99334
rect 422422 99098 422604 99334
rect 422004 63654 422604 99098
rect 422004 63418 422186 63654
rect 422422 63418 422604 63654
rect 422004 63334 422604 63418
rect 422004 63098 422186 63334
rect 422422 63098 422604 63334
rect 420683 61436 420749 61437
rect 420683 61372 420684 61436
rect 420748 61372 420749 61436
rect 420683 61371 420749 61372
rect 418404 59818 418586 60054
rect 418822 59818 419004 60054
rect 418404 59734 419004 59818
rect 418404 59498 418586 59734
rect 418822 59498 419004 59734
rect 418404 24054 419004 59498
rect 420686 48381 420746 61371
rect 420683 48380 420749 48381
rect 420683 48316 420684 48380
rect 420748 48316 420749 48380
rect 420683 48315 420749 48316
rect 420683 42124 420749 42125
rect 420683 42060 420684 42124
rect 420748 42060 420749 42124
rect 420683 42059 420749 42060
rect 420686 29069 420746 42059
rect 420683 29068 420749 29069
rect 420683 29004 420684 29068
rect 420748 29004 420749 29068
rect 420683 29003 420749 29004
rect 418404 23818 418586 24054
rect 418822 23818 419004 24054
rect 418404 23734 419004 23818
rect 418404 23498 418586 23734
rect 418822 23498 419004 23734
rect 418404 -3166 419004 23498
rect 418404 -3402 418586 -3166
rect 418822 -3402 419004 -3166
rect 418404 -3486 419004 -3402
rect 418404 -3722 418586 -3486
rect 418822 -3722 419004 -3486
rect 418404 -3744 419004 -3722
rect 422004 27654 422604 63098
rect 422004 27418 422186 27654
rect 422422 27418 422604 27654
rect 422004 27334 422604 27418
rect 422004 27098 422186 27334
rect 422422 27098 422604 27334
rect 422004 -5046 422604 27098
rect 422004 -5282 422186 -5046
rect 422422 -5282 422604 -5046
rect 422004 -5366 422604 -5282
rect 422004 -5602 422186 -5366
rect 422422 -5602 422604 -5366
rect 422004 -5624 422604 -5602
rect 425604 679254 426204 710862
rect 443604 710478 444204 711440
rect 443604 710242 443786 710478
rect 444022 710242 444204 710478
rect 443604 710158 444204 710242
rect 443604 709922 443786 710158
rect 444022 709922 444204 710158
rect 440004 708598 440604 709560
rect 440004 708362 440186 708598
rect 440422 708362 440604 708598
rect 440004 708278 440604 708362
rect 440004 708042 440186 708278
rect 440422 708042 440604 708278
rect 436404 706718 437004 707680
rect 436404 706482 436586 706718
rect 436822 706482 437004 706718
rect 436404 706398 437004 706482
rect 436404 706162 436586 706398
rect 436822 706162 437004 706398
rect 425604 679018 425786 679254
rect 426022 679018 426204 679254
rect 425604 678934 426204 679018
rect 425604 678698 425786 678934
rect 426022 678698 426204 678934
rect 425604 643254 426204 678698
rect 425604 643018 425786 643254
rect 426022 643018 426204 643254
rect 425604 642934 426204 643018
rect 425604 642698 425786 642934
rect 426022 642698 426204 642934
rect 425604 607254 426204 642698
rect 425604 607018 425786 607254
rect 426022 607018 426204 607254
rect 425604 606934 426204 607018
rect 425604 606698 425786 606934
rect 426022 606698 426204 606934
rect 425604 571254 426204 606698
rect 425604 571018 425786 571254
rect 426022 571018 426204 571254
rect 425604 570934 426204 571018
rect 425604 570698 425786 570934
rect 426022 570698 426204 570934
rect 425604 535254 426204 570698
rect 425604 535018 425786 535254
rect 426022 535018 426204 535254
rect 425604 534934 426204 535018
rect 425604 534698 425786 534934
rect 426022 534698 426204 534934
rect 425604 499254 426204 534698
rect 425604 499018 425786 499254
rect 426022 499018 426204 499254
rect 425604 498934 426204 499018
rect 425604 498698 425786 498934
rect 426022 498698 426204 498934
rect 425604 463254 426204 498698
rect 425604 463018 425786 463254
rect 426022 463018 426204 463254
rect 425604 462934 426204 463018
rect 425604 462698 425786 462934
rect 426022 462698 426204 462934
rect 425604 427254 426204 462698
rect 425604 427018 425786 427254
rect 426022 427018 426204 427254
rect 425604 426934 426204 427018
rect 425604 426698 425786 426934
rect 426022 426698 426204 426934
rect 425604 391254 426204 426698
rect 425604 391018 425786 391254
rect 426022 391018 426204 391254
rect 425604 390934 426204 391018
rect 425604 390698 425786 390934
rect 426022 390698 426204 390934
rect 425604 355254 426204 390698
rect 425604 355018 425786 355254
rect 426022 355018 426204 355254
rect 425604 354934 426204 355018
rect 425604 354698 425786 354934
rect 426022 354698 426204 354934
rect 425604 319254 426204 354698
rect 425604 319018 425786 319254
rect 426022 319018 426204 319254
rect 425604 318934 426204 319018
rect 425604 318698 425786 318934
rect 426022 318698 426204 318934
rect 425604 283254 426204 318698
rect 425604 283018 425786 283254
rect 426022 283018 426204 283254
rect 425604 282934 426204 283018
rect 425604 282698 425786 282934
rect 426022 282698 426204 282934
rect 425604 247254 426204 282698
rect 425604 247018 425786 247254
rect 426022 247018 426204 247254
rect 425604 246934 426204 247018
rect 425604 246698 425786 246934
rect 426022 246698 426204 246934
rect 425604 211254 426204 246698
rect 425604 211018 425786 211254
rect 426022 211018 426204 211254
rect 425604 210934 426204 211018
rect 425604 210698 425786 210934
rect 426022 210698 426204 210934
rect 425604 175254 426204 210698
rect 425604 175018 425786 175254
rect 426022 175018 426204 175254
rect 425604 174934 426204 175018
rect 425604 174698 425786 174934
rect 426022 174698 426204 174934
rect 425604 139254 426204 174698
rect 425604 139018 425786 139254
rect 426022 139018 426204 139254
rect 425604 138934 426204 139018
rect 425604 138698 425786 138934
rect 426022 138698 426204 138934
rect 425604 103254 426204 138698
rect 425604 103018 425786 103254
rect 426022 103018 426204 103254
rect 425604 102934 426204 103018
rect 425604 102698 425786 102934
rect 426022 102698 426204 102934
rect 425604 67254 426204 102698
rect 425604 67018 425786 67254
rect 426022 67018 426204 67254
rect 425604 66934 426204 67018
rect 425604 66698 425786 66934
rect 426022 66698 426204 66934
rect 425604 31254 426204 66698
rect 425604 31018 425786 31254
rect 426022 31018 426204 31254
rect 425604 30934 426204 31018
rect 425604 30698 425786 30934
rect 426022 30698 426204 30934
rect 407604 -6222 407786 -5986
rect 408022 -6222 408204 -5986
rect 407604 -6306 408204 -6222
rect 407604 -6542 407786 -6306
rect 408022 -6542 408204 -6306
rect 407604 -7504 408204 -6542
rect 425604 -6926 426204 30698
rect 432804 704838 433404 705800
rect 432804 704602 432986 704838
rect 433222 704602 433404 704838
rect 432804 704518 433404 704602
rect 432804 704282 432986 704518
rect 433222 704282 433404 704518
rect 432804 686454 433404 704282
rect 432804 686218 432986 686454
rect 433222 686218 433404 686454
rect 432804 686134 433404 686218
rect 432804 685898 432986 686134
rect 433222 685898 433404 686134
rect 432804 650454 433404 685898
rect 432804 650218 432986 650454
rect 433222 650218 433404 650454
rect 432804 650134 433404 650218
rect 432804 649898 432986 650134
rect 433222 649898 433404 650134
rect 432804 614454 433404 649898
rect 432804 614218 432986 614454
rect 433222 614218 433404 614454
rect 432804 614134 433404 614218
rect 432804 613898 432986 614134
rect 433222 613898 433404 614134
rect 432804 578454 433404 613898
rect 432804 578218 432986 578454
rect 433222 578218 433404 578454
rect 432804 578134 433404 578218
rect 432804 577898 432986 578134
rect 433222 577898 433404 578134
rect 432804 542454 433404 577898
rect 432804 542218 432986 542454
rect 433222 542218 433404 542454
rect 432804 542134 433404 542218
rect 432804 541898 432986 542134
rect 433222 541898 433404 542134
rect 432804 506454 433404 541898
rect 432804 506218 432986 506454
rect 433222 506218 433404 506454
rect 432804 506134 433404 506218
rect 432804 505898 432986 506134
rect 433222 505898 433404 506134
rect 432804 470454 433404 505898
rect 432804 470218 432986 470454
rect 433222 470218 433404 470454
rect 432804 470134 433404 470218
rect 432804 469898 432986 470134
rect 433222 469898 433404 470134
rect 432804 434454 433404 469898
rect 432804 434218 432986 434454
rect 433222 434218 433404 434454
rect 432804 434134 433404 434218
rect 432804 433898 432986 434134
rect 433222 433898 433404 434134
rect 432804 398454 433404 433898
rect 432804 398218 432986 398454
rect 433222 398218 433404 398454
rect 432804 398134 433404 398218
rect 432804 397898 432986 398134
rect 433222 397898 433404 398134
rect 432804 362454 433404 397898
rect 432804 362218 432986 362454
rect 433222 362218 433404 362454
rect 432804 362134 433404 362218
rect 432804 361898 432986 362134
rect 433222 361898 433404 362134
rect 432804 326454 433404 361898
rect 432804 326218 432986 326454
rect 433222 326218 433404 326454
rect 432804 326134 433404 326218
rect 432804 325898 432986 326134
rect 433222 325898 433404 326134
rect 432804 290454 433404 325898
rect 432804 290218 432986 290454
rect 433222 290218 433404 290454
rect 432804 290134 433404 290218
rect 432804 289898 432986 290134
rect 433222 289898 433404 290134
rect 432804 254454 433404 289898
rect 432804 254218 432986 254454
rect 433222 254218 433404 254454
rect 432804 254134 433404 254218
rect 432804 253898 432986 254134
rect 433222 253898 433404 254134
rect 432804 218454 433404 253898
rect 432804 218218 432986 218454
rect 433222 218218 433404 218454
rect 432804 218134 433404 218218
rect 432804 217898 432986 218134
rect 433222 217898 433404 218134
rect 432804 182454 433404 217898
rect 432804 182218 432986 182454
rect 433222 182218 433404 182454
rect 432804 182134 433404 182218
rect 432804 181898 432986 182134
rect 433222 181898 433404 182134
rect 432804 146454 433404 181898
rect 432804 146218 432986 146454
rect 433222 146218 433404 146454
rect 432804 146134 433404 146218
rect 432804 145898 432986 146134
rect 433222 145898 433404 146134
rect 432804 110454 433404 145898
rect 432804 110218 432986 110454
rect 433222 110218 433404 110454
rect 432804 110134 433404 110218
rect 432804 109898 432986 110134
rect 433222 109898 433404 110134
rect 432804 74454 433404 109898
rect 432804 74218 432986 74454
rect 433222 74218 433404 74454
rect 432804 74134 433404 74218
rect 432804 73898 432986 74134
rect 433222 73898 433404 74134
rect 432804 38454 433404 73898
rect 432804 38218 432986 38454
rect 433222 38218 433404 38454
rect 432804 38134 433404 38218
rect 432804 37898 432986 38134
rect 433222 37898 433404 38134
rect 432804 2454 433404 37898
rect 432804 2218 432986 2454
rect 433222 2218 433404 2454
rect 432804 2134 433404 2218
rect 432804 1898 432986 2134
rect 433222 1898 433404 2134
rect 432804 -346 433404 1898
rect 432804 -582 432986 -346
rect 433222 -582 433404 -346
rect 432804 -666 433404 -582
rect 432804 -902 432986 -666
rect 433222 -902 433404 -666
rect 432804 -1864 433404 -902
rect 436404 690054 437004 706162
rect 436404 689818 436586 690054
rect 436822 689818 437004 690054
rect 436404 689734 437004 689818
rect 436404 689498 436586 689734
rect 436822 689498 437004 689734
rect 436404 654054 437004 689498
rect 436404 653818 436586 654054
rect 436822 653818 437004 654054
rect 436404 653734 437004 653818
rect 436404 653498 436586 653734
rect 436822 653498 437004 653734
rect 436404 618054 437004 653498
rect 436404 617818 436586 618054
rect 436822 617818 437004 618054
rect 436404 617734 437004 617818
rect 436404 617498 436586 617734
rect 436822 617498 437004 617734
rect 436404 582054 437004 617498
rect 436404 581818 436586 582054
rect 436822 581818 437004 582054
rect 436404 581734 437004 581818
rect 436404 581498 436586 581734
rect 436822 581498 437004 581734
rect 436404 546054 437004 581498
rect 436404 545818 436586 546054
rect 436822 545818 437004 546054
rect 436404 545734 437004 545818
rect 436404 545498 436586 545734
rect 436822 545498 437004 545734
rect 436404 510054 437004 545498
rect 436404 509818 436586 510054
rect 436822 509818 437004 510054
rect 436404 509734 437004 509818
rect 436404 509498 436586 509734
rect 436822 509498 437004 509734
rect 436404 474054 437004 509498
rect 436404 473818 436586 474054
rect 436822 473818 437004 474054
rect 436404 473734 437004 473818
rect 436404 473498 436586 473734
rect 436822 473498 437004 473734
rect 436404 438054 437004 473498
rect 436404 437818 436586 438054
rect 436822 437818 437004 438054
rect 436404 437734 437004 437818
rect 436404 437498 436586 437734
rect 436822 437498 437004 437734
rect 436404 402054 437004 437498
rect 436404 401818 436586 402054
rect 436822 401818 437004 402054
rect 436404 401734 437004 401818
rect 436404 401498 436586 401734
rect 436822 401498 437004 401734
rect 436404 366054 437004 401498
rect 436404 365818 436586 366054
rect 436822 365818 437004 366054
rect 436404 365734 437004 365818
rect 436404 365498 436586 365734
rect 436822 365498 437004 365734
rect 436404 330054 437004 365498
rect 436404 329818 436586 330054
rect 436822 329818 437004 330054
rect 436404 329734 437004 329818
rect 436404 329498 436586 329734
rect 436822 329498 437004 329734
rect 436404 294054 437004 329498
rect 436404 293818 436586 294054
rect 436822 293818 437004 294054
rect 436404 293734 437004 293818
rect 436404 293498 436586 293734
rect 436822 293498 437004 293734
rect 436404 258054 437004 293498
rect 436404 257818 436586 258054
rect 436822 257818 437004 258054
rect 436404 257734 437004 257818
rect 436404 257498 436586 257734
rect 436822 257498 437004 257734
rect 436404 222054 437004 257498
rect 436404 221818 436586 222054
rect 436822 221818 437004 222054
rect 436404 221734 437004 221818
rect 436404 221498 436586 221734
rect 436822 221498 437004 221734
rect 436404 186054 437004 221498
rect 436404 185818 436586 186054
rect 436822 185818 437004 186054
rect 436404 185734 437004 185818
rect 436404 185498 436586 185734
rect 436822 185498 437004 185734
rect 436404 150054 437004 185498
rect 436404 149818 436586 150054
rect 436822 149818 437004 150054
rect 436404 149734 437004 149818
rect 436404 149498 436586 149734
rect 436822 149498 437004 149734
rect 436404 114054 437004 149498
rect 436404 113818 436586 114054
rect 436822 113818 437004 114054
rect 436404 113734 437004 113818
rect 436404 113498 436586 113734
rect 436822 113498 437004 113734
rect 436404 78054 437004 113498
rect 436404 77818 436586 78054
rect 436822 77818 437004 78054
rect 436404 77734 437004 77818
rect 436404 77498 436586 77734
rect 436822 77498 437004 77734
rect 436404 42054 437004 77498
rect 436404 41818 436586 42054
rect 436822 41818 437004 42054
rect 436404 41734 437004 41818
rect 436404 41498 436586 41734
rect 436822 41498 437004 41734
rect 436404 6054 437004 41498
rect 436404 5818 436586 6054
rect 436822 5818 437004 6054
rect 436404 5734 437004 5818
rect 436404 5498 436586 5734
rect 436822 5498 437004 5734
rect 436404 -2226 437004 5498
rect 436404 -2462 436586 -2226
rect 436822 -2462 437004 -2226
rect 436404 -2546 437004 -2462
rect 436404 -2782 436586 -2546
rect 436822 -2782 437004 -2546
rect 436404 -3744 437004 -2782
rect 440004 693654 440604 708042
rect 440004 693418 440186 693654
rect 440422 693418 440604 693654
rect 440004 693334 440604 693418
rect 440004 693098 440186 693334
rect 440422 693098 440604 693334
rect 440004 657654 440604 693098
rect 440004 657418 440186 657654
rect 440422 657418 440604 657654
rect 440004 657334 440604 657418
rect 440004 657098 440186 657334
rect 440422 657098 440604 657334
rect 440004 621654 440604 657098
rect 440004 621418 440186 621654
rect 440422 621418 440604 621654
rect 440004 621334 440604 621418
rect 440004 621098 440186 621334
rect 440422 621098 440604 621334
rect 440004 585654 440604 621098
rect 440004 585418 440186 585654
rect 440422 585418 440604 585654
rect 440004 585334 440604 585418
rect 440004 585098 440186 585334
rect 440422 585098 440604 585334
rect 440004 549654 440604 585098
rect 440004 549418 440186 549654
rect 440422 549418 440604 549654
rect 440004 549334 440604 549418
rect 440004 549098 440186 549334
rect 440422 549098 440604 549334
rect 440004 513654 440604 549098
rect 440004 513418 440186 513654
rect 440422 513418 440604 513654
rect 440004 513334 440604 513418
rect 440004 513098 440186 513334
rect 440422 513098 440604 513334
rect 440004 477654 440604 513098
rect 440004 477418 440186 477654
rect 440422 477418 440604 477654
rect 440004 477334 440604 477418
rect 440004 477098 440186 477334
rect 440422 477098 440604 477334
rect 440004 441654 440604 477098
rect 440004 441418 440186 441654
rect 440422 441418 440604 441654
rect 440004 441334 440604 441418
rect 440004 441098 440186 441334
rect 440422 441098 440604 441334
rect 440004 405654 440604 441098
rect 440004 405418 440186 405654
rect 440422 405418 440604 405654
rect 440004 405334 440604 405418
rect 440004 405098 440186 405334
rect 440422 405098 440604 405334
rect 440004 369654 440604 405098
rect 440004 369418 440186 369654
rect 440422 369418 440604 369654
rect 440004 369334 440604 369418
rect 440004 369098 440186 369334
rect 440422 369098 440604 369334
rect 440004 333654 440604 369098
rect 440004 333418 440186 333654
rect 440422 333418 440604 333654
rect 440004 333334 440604 333418
rect 440004 333098 440186 333334
rect 440422 333098 440604 333334
rect 440004 297654 440604 333098
rect 440004 297418 440186 297654
rect 440422 297418 440604 297654
rect 440004 297334 440604 297418
rect 440004 297098 440186 297334
rect 440422 297098 440604 297334
rect 440004 261654 440604 297098
rect 440004 261418 440186 261654
rect 440422 261418 440604 261654
rect 440004 261334 440604 261418
rect 440004 261098 440186 261334
rect 440422 261098 440604 261334
rect 440004 225654 440604 261098
rect 440004 225418 440186 225654
rect 440422 225418 440604 225654
rect 440004 225334 440604 225418
rect 440004 225098 440186 225334
rect 440422 225098 440604 225334
rect 440004 189654 440604 225098
rect 440004 189418 440186 189654
rect 440422 189418 440604 189654
rect 440004 189334 440604 189418
rect 440004 189098 440186 189334
rect 440422 189098 440604 189334
rect 440004 153654 440604 189098
rect 440004 153418 440186 153654
rect 440422 153418 440604 153654
rect 440004 153334 440604 153418
rect 440004 153098 440186 153334
rect 440422 153098 440604 153334
rect 440004 117654 440604 153098
rect 440004 117418 440186 117654
rect 440422 117418 440604 117654
rect 440004 117334 440604 117418
rect 440004 117098 440186 117334
rect 440422 117098 440604 117334
rect 440004 81654 440604 117098
rect 440004 81418 440186 81654
rect 440422 81418 440604 81654
rect 440004 81334 440604 81418
rect 440004 81098 440186 81334
rect 440422 81098 440604 81334
rect 440004 45654 440604 81098
rect 440004 45418 440186 45654
rect 440422 45418 440604 45654
rect 440004 45334 440604 45418
rect 440004 45098 440186 45334
rect 440422 45098 440604 45334
rect 440004 9654 440604 45098
rect 440004 9418 440186 9654
rect 440422 9418 440604 9654
rect 440004 9334 440604 9418
rect 440004 9098 440186 9334
rect 440422 9098 440604 9334
rect 440004 -4106 440604 9098
rect 440004 -4342 440186 -4106
rect 440422 -4342 440604 -4106
rect 440004 -4426 440604 -4342
rect 440004 -4662 440186 -4426
rect 440422 -4662 440604 -4426
rect 440004 -5624 440604 -4662
rect 443604 697254 444204 709922
rect 461604 711418 462204 711440
rect 461604 711182 461786 711418
rect 462022 711182 462204 711418
rect 461604 711098 462204 711182
rect 461604 710862 461786 711098
rect 462022 710862 462204 711098
rect 458004 709538 458604 709560
rect 458004 709302 458186 709538
rect 458422 709302 458604 709538
rect 458004 709218 458604 709302
rect 458004 708982 458186 709218
rect 458422 708982 458604 709218
rect 454404 707658 455004 707680
rect 454404 707422 454586 707658
rect 454822 707422 455004 707658
rect 454404 707338 455004 707422
rect 454404 707102 454586 707338
rect 454822 707102 455004 707338
rect 443604 697018 443786 697254
rect 444022 697018 444204 697254
rect 443604 696934 444204 697018
rect 443604 696698 443786 696934
rect 444022 696698 444204 696934
rect 443604 661254 444204 696698
rect 443604 661018 443786 661254
rect 444022 661018 444204 661254
rect 443604 660934 444204 661018
rect 443604 660698 443786 660934
rect 444022 660698 444204 660934
rect 443604 625254 444204 660698
rect 443604 625018 443786 625254
rect 444022 625018 444204 625254
rect 443604 624934 444204 625018
rect 443604 624698 443786 624934
rect 444022 624698 444204 624934
rect 443604 589254 444204 624698
rect 443604 589018 443786 589254
rect 444022 589018 444204 589254
rect 443604 588934 444204 589018
rect 443604 588698 443786 588934
rect 444022 588698 444204 588934
rect 443604 553254 444204 588698
rect 443604 553018 443786 553254
rect 444022 553018 444204 553254
rect 443604 552934 444204 553018
rect 443604 552698 443786 552934
rect 444022 552698 444204 552934
rect 443604 517254 444204 552698
rect 443604 517018 443786 517254
rect 444022 517018 444204 517254
rect 443604 516934 444204 517018
rect 443604 516698 443786 516934
rect 444022 516698 444204 516934
rect 443604 481254 444204 516698
rect 443604 481018 443786 481254
rect 444022 481018 444204 481254
rect 443604 480934 444204 481018
rect 443604 480698 443786 480934
rect 444022 480698 444204 480934
rect 443604 445254 444204 480698
rect 443604 445018 443786 445254
rect 444022 445018 444204 445254
rect 443604 444934 444204 445018
rect 443604 444698 443786 444934
rect 444022 444698 444204 444934
rect 443604 409254 444204 444698
rect 443604 409018 443786 409254
rect 444022 409018 444204 409254
rect 443604 408934 444204 409018
rect 443604 408698 443786 408934
rect 444022 408698 444204 408934
rect 443604 373254 444204 408698
rect 443604 373018 443786 373254
rect 444022 373018 444204 373254
rect 443604 372934 444204 373018
rect 443604 372698 443786 372934
rect 444022 372698 444204 372934
rect 443604 337254 444204 372698
rect 443604 337018 443786 337254
rect 444022 337018 444204 337254
rect 443604 336934 444204 337018
rect 443604 336698 443786 336934
rect 444022 336698 444204 336934
rect 443604 301254 444204 336698
rect 443604 301018 443786 301254
rect 444022 301018 444204 301254
rect 443604 300934 444204 301018
rect 443604 300698 443786 300934
rect 444022 300698 444204 300934
rect 443604 265254 444204 300698
rect 443604 265018 443786 265254
rect 444022 265018 444204 265254
rect 443604 264934 444204 265018
rect 443604 264698 443786 264934
rect 444022 264698 444204 264934
rect 443604 229254 444204 264698
rect 443604 229018 443786 229254
rect 444022 229018 444204 229254
rect 443604 228934 444204 229018
rect 443604 228698 443786 228934
rect 444022 228698 444204 228934
rect 443604 193254 444204 228698
rect 443604 193018 443786 193254
rect 444022 193018 444204 193254
rect 443604 192934 444204 193018
rect 443604 192698 443786 192934
rect 444022 192698 444204 192934
rect 443604 157254 444204 192698
rect 443604 157018 443786 157254
rect 444022 157018 444204 157254
rect 443604 156934 444204 157018
rect 443604 156698 443786 156934
rect 444022 156698 444204 156934
rect 443604 121254 444204 156698
rect 443604 121018 443786 121254
rect 444022 121018 444204 121254
rect 443604 120934 444204 121018
rect 443604 120698 443786 120934
rect 444022 120698 444204 120934
rect 443604 85254 444204 120698
rect 443604 85018 443786 85254
rect 444022 85018 444204 85254
rect 443604 84934 444204 85018
rect 443604 84698 443786 84934
rect 444022 84698 444204 84934
rect 443604 49254 444204 84698
rect 443604 49018 443786 49254
rect 444022 49018 444204 49254
rect 443604 48934 444204 49018
rect 443604 48698 443786 48934
rect 444022 48698 444204 48934
rect 443604 13254 444204 48698
rect 443604 13018 443786 13254
rect 444022 13018 444204 13254
rect 443604 12934 444204 13018
rect 443604 12698 443786 12934
rect 444022 12698 444204 12934
rect 425604 -7162 425786 -6926
rect 426022 -7162 426204 -6926
rect 425604 -7246 426204 -7162
rect 425604 -7482 425786 -7246
rect 426022 -7482 426204 -7246
rect 425604 -7504 426204 -7482
rect 443604 -5986 444204 12698
rect 450804 705778 451404 705800
rect 450804 705542 450986 705778
rect 451222 705542 451404 705778
rect 450804 705458 451404 705542
rect 450804 705222 450986 705458
rect 451222 705222 451404 705458
rect 450804 668454 451404 705222
rect 450804 668218 450986 668454
rect 451222 668218 451404 668454
rect 450804 668134 451404 668218
rect 450804 667898 450986 668134
rect 451222 667898 451404 668134
rect 450804 632454 451404 667898
rect 450804 632218 450986 632454
rect 451222 632218 451404 632454
rect 450804 632134 451404 632218
rect 450804 631898 450986 632134
rect 451222 631898 451404 632134
rect 450804 596454 451404 631898
rect 450804 596218 450986 596454
rect 451222 596218 451404 596454
rect 450804 596134 451404 596218
rect 450804 595898 450986 596134
rect 451222 595898 451404 596134
rect 450804 560454 451404 595898
rect 450804 560218 450986 560454
rect 451222 560218 451404 560454
rect 450804 560134 451404 560218
rect 450804 559898 450986 560134
rect 451222 559898 451404 560134
rect 450804 524454 451404 559898
rect 450804 524218 450986 524454
rect 451222 524218 451404 524454
rect 450804 524134 451404 524218
rect 450804 523898 450986 524134
rect 451222 523898 451404 524134
rect 450804 488454 451404 523898
rect 450804 488218 450986 488454
rect 451222 488218 451404 488454
rect 450804 488134 451404 488218
rect 450804 487898 450986 488134
rect 451222 487898 451404 488134
rect 450804 452454 451404 487898
rect 450804 452218 450986 452454
rect 451222 452218 451404 452454
rect 450804 452134 451404 452218
rect 450804 451898 450986 452134
rect 451222 451898 451404 452134
rect 450804 416454 451404 451898
rect 450804 416218 450986 416454
rect 451222 416218 451404 416454
rect 450804 416134 451404 416218
rect 450804 415898 450986 416134
rect 451222 415898 451404 416134
rect 450804 380454 451404 415898
rect 450804 380218 450986 380454
rect 451222 380218 451404 380454
rect 450804 380134 451404 380218
rect 450804 379898 450986 380134
rect 451222 379898 451404 380134
rect 450804 344454 451404 379898
rect 450804 344218 450986 344454
rect 451222 344218 451404 344454
rect 450804 344134 451404 344218
rect 450804 343898 450986 344134
rect 451222 343898 451404 344134
rect 450804 308454 451404 343898
rect 450804 308218 450986 308454
rect 451222 308218 451404 308454
rect 450804 308134 451404 308218
rect 450804 307898 450986 308134
rect 451222 307898 451404 308134
rect 450804 272454 451404 307898
rect 450804 272218 450986 272454
rect 451222 272218 451404 272454
rect 450804 272134 451404 272218
rect 450804 271898 450986 272134
rect 451222 271898 451404 272134
rect 450804 236454 451404 271898
rect 450804 236218 450986 236454
rect 451222 236218 451404 236454
rect 450804 236134 451404 236218
rect 450804 235898 450986 236134
rect 451222 235898 451404 236134
rect 450804 200454 451404 235898
rect 450804 200218 450986 200454
rect 451222 200218 451404 200454
rect 450804 200134 451404 200218
rect 450804 199898 450986 200134
rect 451222 199898 451404 200134
rect 450804 164454 451404 199898
rect 450804 164218 450986 164454
rect 451222 164218 451404 164454
rect 450804 164134 451404 164218
rect 450804 163898 450986 164134
rect 451222 163898 451404 164134
rect 450804 128454 451404 163898
rect 450804 128218 450986 128454
rect 451222 128218 451404 128454
rect 450804 128134 451404 128218
rect 450804 127898 450986 128134
rect 451222 127898 451404 128134
rect 450804 92454 451404 127898
rect 450804 92218 450986 92454
rect 451222 92218 451404 92454
rect 450804 92134 451404 92218
rect 450804 91898 450986 92134
rect 451222 91898 451404 92134
rect 450804 56454 451404 91898
rect 450804 56218 450986 56454
rect 451222 56218 451404 56454
rect 450804 56134 451404 56218
rect 450804 55898 450986 56134
rect 451222 55898 451404 56134
rect 450804 20454 451404 55898
rect 450804 20218 450986 20454
rect 451222 20218 451404 20454
rect 450804 20134 451404 20218
rect 450804 19898 450986 20134
rect 451222 19898 451404 20134
rect 450804 -1286 451404 19898
rect 450804 -1522 450986 -1286
rect 451222 -1522 451404 -1286
rect 450804 -1606 451404 -1522
rect 450804 -1842 450986 -1606
rect 451222 -1842 451404 -1606
rect 450804 -1864 451404 -1842
rect 454404 672054 455004 707102
rect 454404 671818 454586 672054
rect 454822 671818 455004 672054
rect 454404 671734 455004 671818
rect 454404 671498 454586 671734
rect 454822 671498 455004 671734
rect 454404 636054 455004 671498
rect 454404 635818 454586 636054
rect 454822 635818 455004 636054
rect 454404 635734 455004 635818
rect 454404 635498 454586 635734
rect 454822 635498 455004 635734
rect 454404 600054 455004 635498
rect 454404 599818 454586 600054
rect 454822 599818 455004 600054
rect 454404 599734 455004 599818
rect 454404 599498 454586 599734
rect 454822 599498 455004 599734
rect 454404 564054 455004 599498
rect 454404 563818 454586 564054
rect 454822 563818 455004 564054
rect 454404 563734 455004 563818
rect 454404 563498 454586 563734
rect 454822 563498 455004 563734
rect 454404 528054 455004 563498
rect 454404 527818 454586 528054
rect 454822 527818 455004 528054
rect 454404 527734 455004 527818
rect 454404 527498 454586 527734
rect 454822 527498 455004 527734
rect 454404 492054 455004 527498
rect 454404 491818 454586 492054
rect 454822 491818 455004 492054
rect 454404 491734 455004 491818
rect 454404 491498 454586 491734
rect 454822 491498 455004 491734
rect 454404 456054 455004 491498
rect 454404 455818 454586 456054
rect 454822 455818 455004 456054
rect 454404 455734 455004 455818
rect 454404 455498 454586 455734
rect 454822 455498 455004 455734
rect 454404 420054 455004 455498
rect 454404 419818 454586 420054
rect 454822 419818 455004 420054
rect 454404 419734 455004 419818
rect 454404 419498 454586 419734
rect 454822 419498 455004 419734
rect 454404 384054 455004 419498
rect 454404 383818 454586 384054
rect 454822 383818 455004 384054
rect 454404 383734 455004 383818
rect 454404 383498 454586 383734
rect 454822 383498 455004 383734
rect 454404 348054 455004 383498
rect 454404 347818 454586 348054
rect 454822 347818 455004 348054
rect 454404 347734 455004 347818
rect 454404 347498 454586 347734
rect 454822 347498 455004 347734
rect 454404 312054 455004 347498
rect 454404 311818 454586 312054
rect 454822 311818 455004 312054
rect 454404 311734 455004 311818
rect 454404 311498 454586 311734
rect 454822 311498 455004 311734
rect 454404 276054 455004 311498
rect 454404 275818 454586 276054
rect 454822 275818 455004 276054
rect 454404 275734 455004 275818
rect 454404 275498 454586 275734
rect 454822 275498 455004 275734
rect 454404 240054 455004 275498
rect 454404 239818 454586 240054
rect 454822 239818 455004 240054
rect 454404 239734 455004 239818
rect 454404 239498 454586 239734
rect 454822 239498 455004 239734
rect 454404 204054 455004 239498
rect 454404 203818 454586 204054
rect 454822 203818 455004 204054
rect 454404 203734 455004 203818
rect 454404 203498 454586 203734
rect 454822 203498 455004 203734
rect 454404 168054 455004 203498
rect 454404 167818 454586 168054
rect 454822 167818 455004 168054
rect 454404 167734 455004 167818
rect 454404 167498 454586 167734
rect 454822 167498 455004 167734
rect 454404 132054 455004 167498
rect 454404 131818 454586 132054
rect 454822 131818 455004 132054
rect 454404 131734 455004 131818
rect 454404 131498 454586 131734
rect 454822 131498 455004 131734
rect 454404 96054 455004 131498
rect 454404 95818 454586 96054
rect 454822 95818 455004 96054
rect 454404 95734 455004 95818
rect 454404 95498 454586 95734
rect 454822 95498 455004 95734
rect 454404 60054 455004 95498
rect 454404 59818 454586 60054
rect 454822 59818 455004 60054
rect 454404 59734 455004 59818
rect 454404 59498 454586 59734
rect 454822 59498 455004 59734
rect 454404 24054 455004 59498
rect 454404 23818 454586 24054
rect 454822 23818 455004 24054
rect 454404 23734 455004 23818
rect 454404 23498 454586 23734
rect 454822 23498 455004 23734
rect 454404 -3166 455004 23498
rect 454404 -3402 454586 -3166
rect 454822 -3402 455004 -3166
rect 454404 -3486 455004 -3402
rect 454404 -3722 454586 -3486
rect 454822 -3722 455004 -3486
rect 454404 -3744 455004 -3722
rect 458004 675654 458604 708982
rect 458004 675418 458186 675654
rect 458422 675418 458604 675654
rect 458004 675334 458604 675418
rect 458004 675098 458186 675334
rect 458422 675098 458604 675334
rect 458004 639654 458604 675098
rect 458004 639418 458186 639654
rect 458422 639418 458604 639654
rect 458004 639334 458604 639418
rect 458004 639098 458186 639334
rect 458422 639098 458604 639334
rect 458004 603654 458604 639098
rect 458004 603418 458186 603654
rect 458422 603418 458604 603654
rect 458004 603334 458604 603418
rect 458004 603098 458186 603334
rect 458422 603098 458604 603334
rect 458004 567654 458604 603098
rect 458004 567418 458186 567654
rect 458422 567418 458604 567654
rect 458004 567334 458604 567418
rect 458004 567098 458186 567334
rect 458422 567098 458604 567334
rect 458004 531654 458604 567098
rect 458004 531418 458186 531654
rect 458422 531418 458604 531654
rect 458004 531334 458604 531418
rect 458004 531098 458186 531334
rect 458422 531098 458604 531334
rect 458004 495654 458604 531098
rect 458004 495418 458186 495654
rect 458422 495418 458604 495654
rect 458004 495334 458604 495418
rect 458004 495098 458186 495334
rect 458422 495098 458604 495334
rect 458004 459654 458604 495098
rect 458004 459418 458186 459654
rect 458422 459418 458604 459654
rect 458004 459334 458604 459418
rect 458004 459098 458186 459334
rect 458422 459098 458604 459334
rect 458004 423654 458604 459098
rect 458004 423418 458186 423654
rect 458422 423418 458604 423654
rect 458004 423334 458604 423418
rect 458004 423098 458186 423334
rect 458422 423098 458604 423334
rect 458004 387654 458604 423098
rect 458004 387418 458186 387654
rect 458422 387418 458604 387654
rect 458004 387334 458604 387418
rect 458004 387098 458186 387334
rect 458422 387098 458604 387334
rect 458004 351654 458604 387098
rect 458004 351418 458186 351654
rect 458422 351418 458604 351654
rect 458004 351334 458604 351418
rect 458004 351098 458186 351334
rect 458422 351098 458604 351334
rect 458004 315654 458604 351098
rect 458004 315418 458186 315654
rect 458422 315418 458604 315654
rect 458004 315334 458604 315418
rect 458004 315098 458186 315334
rect 458422 315098 458604 315334
rect 458004 279654 458604 315098
rect 458004 279418 458186 279654
rect 458422 279418 458604 279654
rect 458004 279334 458604 279418
rect 458004 279098 458186 279334
rect 458422 279098 458604 279334
rect 458004 243654 458604 279098
rect 458004 243418 458186 243654
rect 458422 243418 458604 243654
rect 458004 243334 458604 243418
rect 458004 243098 458186 243334
rect 458422 243098 458604 243334
rect 458004 207654 458604 243098
rect 458004 207418 458186 207654
rect 458422 207418 458604 207654
rect 458004 207334 458604 207418
rect 458004 207098 458186 207334
rect 458422 207098 458604 207334
rect 458004 171654 458604 207098
rect 458004 171418 458186 171654
rect 458422 171418 458604 171654
rect 458004 171334 458604 171418
rect 458004 171098 458186 171334
rect 458422 171098 458604 171334
rect 458004 135654 458604 171098
rect 458004 135418 458186 135654
rect 458422 135418 458604 135654
rect 458004 135334 458604 135418
rect 458004 135098 458186 135334
rect 458422 135098 458604 135334
rect 458004 99654 458604 135098
rect 458004 99418 458186 99654
rect 458422 99418 458604 99654
rect 458004 99334 458604 99418
rect 458004 99098 458186 99334
rect 458422 99098 458604 99334
rect 458004 63654 458604 99098
rect 458004 63418 458186 63654
rect 458422 63418 458604 63654
rect 458004 63334 458604 63418
rect 458004 63098 458186 63334
rect 458422 63098 458604 63334
rect 458004 27654 458604 63098
rect 458004 27418 458186 27654
rect 458422 27418 458604 27654
rect 458004 27334 458604 27418
rect 458004 27098 458186 27334
rect 458422 27098 458604 27334
rect 458004 -5046 458604 27098
rect 458004 -5282 458186 -5046
rect 458422 -5282 458604 -5046
rect 458004 -5366 458604 -5282
rect 458004 -5602 458186 -5366
rect 458422 -5602 458604 -5366
rect 458004 -5624 458604 -5602
rect 461604 679254 462204 710862
rect 479604 710478 480204 711440
rect 479604 710242 479786 710478
rect 480022 710242 480204 710478
rect 479604 710158 480204 710242
rect 479604 709922 479786 710158
rect 480022 709922 480204 710158
rect 476004 708598 476604 709560
rect 476004 708362 476186 708598
rect 476422 708362 476604 708598
rect 476004 708278 476604 708362
rect 476004 708042 476186 708278
rect 476422 708042 476604 708278
rect 472404 706718 473004 707680
rect 472404 706482 472586 706718
rect 472822 706482 473004 706718
rect 472404 706398 473004 706482
rect 472404 706162 472586 706398
rect 472822 706162 473004 706398
rect 461604 679018 461786 679254
rect 462022 679018 462204 679254
rect 461604 678934 462204 679018
rect 461604 678698 461786 678934
rect 462022 678698 462204 678934
rect 461604 643254 462204 678698
rect 461604 643018 461786 643254
rect 462022 643018 462204 643254
rect 461604 642934 462204 643018
rect 461604 642698 461786 642934
rect 462022 642698 462204 642934
rect 461604 607254 462204 642698
rect 461604 607018 461786 607254
rect 462022 607018 462204 607254
rect 461604 606934 462204 607018
rect 461604 606698 461786 606934
rect 462022 606698 462204 606934
rect 461604 571254 462204 606698
rect 461604 571018 461786 571254
rect 462022 571018 462204 571254
rect 461604 570934 462204 571018
rect 461604 570698 461786 570934
rect 462022 570698 462204 570934
rect 461604 535254 462204 570698
rect 461604 535018 461786 535254
rect 462022 535018 462204 535254
rect 461604 534934 462204 535018
rect 461604 534698 461786 534934
rect 462022 534698 462204 534934
rect 461604 499254 462204 534698
rect 461604 499018 461786 499254
rect 462022 499018 462204 499254
rect 461604 498934 462204 499018
rect 461604 498698 461786 498934
rect 462022 498698 462204 498934
rect 461604 463254 462204 498698
rect 461604 463018 461786 463254
rect 462022 463018 462204 463254
rect 461604 462934 462204 463018
rect 461604 462698 461786 462934
rect 462022 462698 462204 462934
rect 461604 427254 462204 462698
rect 461604 427018 461786 427254
rect 462022 427018 462204 427254
rect 461604 426934 462204 427018
rect 461604 426698 461786 426934
rect 462022 426698 462204 426934
rect 461604 391254 462204 426698
rect 461604 391018 461786 391254
rect 462022 391018 462204 391254
rect 461604 390934 462204 391018
rect 461604 390698 461786 390934
rect 462022 390698 462204 390934
rect 461604 355254 462204 390698
rect 461604 355018 461786 355254
rect 462022 355018 462204 355254
rect 461604 354934 462204 355018
rect 461604 354698 461786 354934
rect 462022 354698 462204 354934
rect 461604 319254 462204 354698
rect 461604 319018 461786 319254
rect 462022 319018 462204 319254
rect 461604 318934 462204 319018
rect 461604 318698 461786 318934
rect 462022 318698 462204 318934
rect 461604 283254 462204 318698
rect 461604 283018 461786 283254
rect 462022 283018 462204 283254
rect 461604 282934 462204 283018
rect 461604 282698 461786 282934
rect 462022 282698 462204 282934
rect 461604 247254 462204 282698
rect 461604 247018 461786 247254
rect 462022 247018 462204 247254
rect 461604 246934 462204 247018
rect 461604 246698 461786 246934
rect 462022 246698 462204 246934
rect 461604 211254 462204 246698
rect 461604 211018 461786 211254
rect 462022 211018 462204 211254
rect 461604 210934 462204 211018
rect 461604 210698 461786 210934
rect 462022 210698 462204 210934
rect 461604 175254 462204 210698
rect 461604 175018 461786 175254
rect 462022 175018 462204 175254
rect 461604 174934 462204 175018
rect 461604 174698 461786 174934
rect 462022 174698 462204 174934
rect 461604 139254 462204 174698
rect 461604 139018 461786 139254
rect 462022 139018 462204 139254
rect 461604 138934 462204 139018
rect 461604 138698 461786 138934
rect 462022 138698 462204 138934
rect 461604 103254 462204 138698
rect 461604 103018 461786 103254
rect 462022 103018 462204 103254
rect 461604 102934 462204 103018
rect 461604 102698 461786 102934
rect 462022 102698 462204 102934
rect 461604 67254 462204 102698
rect 461604 67018 461786 67254
rect 462022 67018 462204 67254
rect 461604 66934 462204 67018
rect 461604 66698 461786 66934
rect 462022 66698 462204 66934
rect 461604 31254 462204 66698
rect 461604 31018 461786 31254
rect 462022 31018 462204 31254
rect 461604 30934 462204 31018
rect 461604 30698 461786 30934
rect 462022 30698 462204 30934
rect 443604 -6222 443786 -5986
rect 444022 -6222 444204 -5986
rect 443604 -6306 444204 -6222
rect 443604 -6542 443786 -6306
rect 444022 -6542 444204 -6306
rect 443604 -7504 444204 -6542
rect 461604 -6926 462204 30698
rect 468804 704838 469404 705800
rect 468804 704602 468986 704838
rect 469222 704602 469404 704838
rect 468804 704518 469404 704602
rect 468804 704282 468986 704518
rect 469222 704282 469404 704518
rect 468804 686454 469404 704282
rect 468804 686218 468986 686454
rect 469222 686218 469404 686454
rect 468804 686134 469404 686218
rect 468804 685898 468986 686134
rect 469222 685898 469404 686134
rect 468804 650454 469404 685898
rect 468804 650218 468986 650454
rect 469222 650218 469404 650454
rect 468804 650134 469404 650218
rect 468804 649898 468986 650134
rect 469222 649898 469404 650134
rect 468804 614454 469404 649898
rect 468804 614218 468986 614454
rect 469222 614218 469404 614454
rect 468804 614134 469404 614218
rect 468804 613898 468986 614134
rect 469222 613898 469404 614134
rect 468804 578454 469404 613898
rect 468804 578218 468986 578454
rect 469222 578218 469404 578454
rect 468804 578134 469404 578218
rect 468804 577898 468986 578134
rect 469222 577898 469404 578134
rect 468804 542454 469404 577898
rect 468804 542218 468986 542454
rect 469222 542218 469404 542454
rect 468804 542134 469404 542218
rect 468804 541898 468986 542134
rect 469222 541898 469404 542134
rect 468804 506454 469404 541898
rect 468804 506218 468986 506454
rect 469222 506218 469404 506454
rect 468804 506134 469404 506218
rect 468804 505898 468986 506134
rect 469222 505898 469404 506134
rect 468804 470454 469404 505898
rect 468804 470218 468986 470454
rect 469222 470218 469404 470454
rect 468804 470134 469404 470218
rect 468804 469898 468986 470134
rect 469222 469898 469404 470134
rect 468804 434454 469404 469898
rect 468804 434218 468986 434454
rect 469222 434218 469404 434454
rect 468804 434134 469404 434218
rect 468804 433898 468986 434134
rect 469222 433898 469404 434134
rect 468804 398454 469404 433898
rect 468804 398218 468986 398454
rect 469222 398218 469404 398454
rect 468804 398134 469404 398218
rect 468804 397898 468986 398134
rect 469222 397898 469404 398134
rect 468804 362454 469404 397898
rect 468804 362218 468986 362454
rect 469222 362218 469404 362454
rect 468804 362134 469404 362218
rect 468804 361898 468986 362134
rect 469222 361898 469404 362134
rect 468804 326454 469404 361898
rect 468804 326218 468986 326454
rect 469222 326218 469404 326454
rect 468804 326134 469404 326218
rect 468804 325898 468986 326134
rect 469222 325898 469404 326134
rect 468804 290454 469404 325898
rect 468804 290218 468986 290454
rect 469222 290218 469404 290454
rect 468804 290134 469404 290218
rect 468804 289898 468986 290134
rect 469222 289898 469404 290134
rect 468804 254454 469404 289898
rect 468804 254218 468986 254454
rect 469222 254218 469404 254454
rect 468804 254134 469404 254218
rect 468804 253898 468986 254134
rect 469222 253898 469404 254134
rect 468804 218454 469404 253898
rect 468804 218218 468986 218454
rect 469222 218218 469404 218454
rect 468804 218134 469404 218218
rect 468804 217898 468986 218134
rect 469222 217898 469404 218134
rect 468804 182454 469404 217898
rect 468804 182218 468986 182454
rect 469222 182218 469404 182454
rect 468804 182134 469404 182218
rect 468804 181898 468986 182134
rect 469222 181898 469404 182134
rect 468804 146454 469404 181898
rect 468804 146218 468986 146454
rect 469222 146218 469404 146454
rect 468804 146134 469404 146218
rect 468804 145898 468986 146134
rect 469222 145898 469404 146134
rect 468804 110454 469404 145898
rect 468804 110218 468986 110454
rect 469222 110218 469404 110454
rect 468804 110134 469404 110218
rect 468804 109898 468986 110134
rect 469222 109898 469404 110134
rect 468804 74454 469404 109898
rect 468804 74218 468986 74454
rect 469222 74218 469404 74454
rect 468804 74134 469404 74218
rect 468804 73898 468986 74134
rect 469222 73898 469404 74134
rect 468804 38454 469404 73898
rect 468804 38218 468986 38454
rect 469222 38218 469404 38454
rect 468804 38134 469404 38218
rect 468804 37898 468986 38134
rect 469222 37898 469404 38134
rect 468804 2454 469404 37898
rect 468804 2218 468986 2454
rect 469222 2218 469404 2454
rect 468804 2134 469404 2218
rect 468804 1898 468986 2134
rect 469222 1898 469404 2134
rect 468804 -346 469404 1898
rect 468804 -582 468986 -346
rect 469222 -582 469404 -346
rect 468804 -666 469404 -582
rect 468804 -902 468986 -666
rect 469222 -902 469404 -666
rect 468804 -1864 469404 -902
rect 472404 690054 473004 706162
rect 472404 689818 472586 690054
rect 472822 689818 473004 690054
rect 472404 689734 473004 689818
rect 472404 689498 472586 689734
rect 472822 689498 473004 689734
rect 472404 654054 473004 689498
rect 472404 653818 472586 654054
rect 472822 653818 473004 654054
rect 472404 653734 473004 653818
rect 472404 653498 472586 653734
rect 472822 653498 473004 653734
rect 472404 618054 473004 653498
rect 472404 617818 472586 618054
rect 472822 617818 473004 618054
rect 472404 617734 473004 617818
rect 472404 617498 472586 617734
rect 472822 617498 473004 617734
rect 472404 582054 473004 617498
rect 472404 581818 472586 582054
rect 472822 581818 473004 582054
rect 472404 581734 473004 581818
rect 472404 581498 472586 581734
rect 472822 581498 473004 581734
rect 472404 546054 473004 581498
rect 472404 545818 472586 546054
rect 472822 545818 473004 546054
rect 472404 545734 473004 545818
rect 472404 545498 472586 545734
rect 472822 545498 473004 545734
rect 472404 510054 473004 545498
rect 472404 509818 472586 510054
rect 472822 509818 473004 510054
rect 472404 509734 473004 509818
rect 472404 509498 472586 509734
rect 472822 509498 473004 509734
rect 472404 474054 473004 509498
rect 472404 473818 472586 474054
rect 472822 473818 473004 474054
rect 472404 473734 473004 473818
rect 472404 473498 472586 473734
rect 472822 473498 473004 473734
rect 472404 438054 473004 473498
rect 472404 437818 472586 438054
rect 472822 437818 473004 438054
rect 472404 437734 473004 437818
rect 472404 437498 472586 437734
rect 472822 437498 473004 437734
rect 472404 402054 473004 437498
rect 472404 401818 472586 402054
rect 472822 401818 473004 402054
rect 472404 401734 473004 401818
rect 472404 401498 472586 401734
rect 472822 401498 473004 401734
rect 472404 366054 473004 401498
rect 472404 365818 472586 366054
rect 472822 365818 473004 366054
rect 472404 365734 473004 365818
rect 472404 365498 472586 365734
rect 472822 365498 473004 365734
rect 472404 330054 473004 365498
rect 472404 329818 472586 330054
rect 472822 329818 473004 330054
rect 472404 329734 473004 329818
rect 472404 329498 472586 329734
rect 472822 329498 473004 329734
rect 472404 294054 473004 329498
rect 472404 293818 472586 294054
rect 472822 293818 473004 294054
rect 472404 293734 473004 293818
rect 472404 293498 472586 293734
rect 472822 293498 473004 293734
rect 472404 258054 473004 293498
rect 472404 257818 472586 258054
rect 472822 257818 473004 258054
rect 472404 257734 473004 257818
rect 472404 257498 472586 257734
rect 472822 257498 473004 257734
rect 472404 222054 473004 257498
rect 472404 221818 472586 222054
rect 472822 221818 473004 222054
rect 472404 221734 473004 221818
rect 472404 221498 472586 221734
rect 472822 221498 473004 221734
rect 472404 186054 473004 221498
rect 472404 185818 472586 186054
rect 472822 185818 473004 186054
rect 472404 185734 473004 185818
rect 472404 185498 472586 185734
rect 472822 185498 473004 185734
rect 472404 150054 473004 185498
rect 472404 149818 472586 150054
rect 472822 149818 473004 150054
rect 472404 149734 473004 149818
rect 472404 149498 472586 149734
rect 472822 149498 473004 149734
rect 472404 114054 473004 149498
rect 472404 113818 472586 114054
rect 472822 113818 473004 114054
rect 472404 113734 473004 113818
rect 472404 113498 472586 113734
rect 472822 113498 473004 113734
rect 472404 78054 473004 113498
rect 472404 77818 472586 78054
rect 472822 77818 473004 78054
rect 472404 77734 473004 77818
rect 472404 77498 472586 77734
rect 472822 77498 473004 77734
rect 472404 42054 473004 77498
rect 472404 41818 472586 42054
rect 472822 41818 473004 42054
rect 472404 41734 473004 41818
rect 472404 41498 472586 41734
rect 472822 41498 473004 41734
rect 472404 6054 473004 41498
rect 472404 5818 472586 6054
rect 472822 5818 473004 6054
rect 472404 5734 473004 5818
rect 472404 5498 472586 5734
rect 472822 5498 473004 5734
rect 472404 -2226 473004 5498
rect 472404 -2462 472586 -2226
rect 472822 -2462 473004 -2226
rect 472404 -2546 473004 -2462
rect 472404 -2782 472586 -2546
rect 472822 -2782 473004 -2546
rect 472404 -3744 473004 -2782
rect 476004 693654 476604 708042
rect 476004 693418 476186 693654
rect 476422 693418 476604 693654
rect 476004 693334 476604 693418
rect 476004 693098 476186 693334
rect 476422 693098 476604 693334
rect 476004 657654 476604 693098
rect 476004 657418 476186 657654
rect 476422 657418 476604 657654
rect 476004 657334 476604 657418
rect 476004 657098 476186 657334
rect 476422 657098 476604 657334
rect 476004 621654 476604 657098
rect 476004 621418 476186 621654
rect 476422 621418 476604 621654
rect 476004 621334 476604 621418
rect 476004 621098 476186 621334
rect 476422 621098 476604 621334
rect 476004 585654 476604 621098
rect 476004 585418 476186 585654
rect 476422 585418 476604 585654
rect 476004 585334 476604 585418
rect 476004 585098 476186 585334
rect 476422 585098 476604 585334
rect 476004 549654 476604 585098
rect 476004 549418 476186 549654
rect 476422 549418 476604 549654
rect 476004 549334 476604 549418
rect 476004 549098 476186 549334
rect 476422 549098 476604 549334
rect 476004 513654 476604 549098
rect 476004 513418 476186 513654
rect 476422 513418 476604 513654
rect 476004 513334 476604 513418
rect 476004 513098 476186 513334
rect 476422 513098 476604 513334
rect 476004 477654 476604 513098
rect 476004 477418 476186 477654
rect 476422 477418 476604 477654
rect 476004 477334 476604 477418
rect 476004 477098 476186 477334
rect 476422 477098 476604 477334
rect 476004 441654 476604 477098
rect 476004 441418 476186 441654
rect 476422 441418 476604 441654
rect 476004 441334 476604 441418
rect 476004 441098 476186 441334
rect 476422 441098 476604 441334
rect 476004 405654 476604 441098
rect 476004 405418 476186 405654
rect 476422 405418 476604 405654
rect 476004 405334 476604 405418
rect 476004 405098 476186 405334
rect 476422 405098 476604 405334
rect 476004 369654 476604 405098
rect 476004 369418 476186 369654
rect 476422 369418 476604 369654
rect 476004 369334 476604 369418
rect 476004 369098 476186 369334
rect 476422 369098 476604 369334
rect 476004 333654 476604 369098
rect 476004 333418 476186 333654
rect 476422 333418 476604 333654
rect 476004 333334 476604 333418
rect 476004 333098 476186 333334
rect 476422 333098 476604 333334
rect 476004 297654 476604 333098
rect 476004 297418 476186 297654
rect 476422 297418 476604 297654
rect 476004 297334 476604 297418
rect 476004 297098 476186 297334
rect 476422 297098 476604 297334
rect 476004 261654 476604 297098
rect 476004 261418 476186 261654
rect 476422 261418 476604 261654
rect 476004 261334 476604 261418
rect 476004 261098 476186 261334
rect 476422 261098 476604 261334
rect 476004 225654 476604 261098
rect 476004 225418 476186 225654
rect 476422 225418 476604 225654
rect 476004 225334 476604 225418
rect 476004 225098 476186 225334
rect 476422 225098 476604 225334
rect 476004 189654 476604 225098
rect 476004 189418 476186 189654
rect 476422 189418 476604 189654
rect 476004 189334 476604 189418
rect 476004 189098 476186 189334
rect 476422 189098 476604 189334
rect 476004 153654 476604 189098
rect 476004 153418 476186 153654
rect 476422 153418 476604 153654
rect 476004 153334 476604 153418
rect 476004 153098 476186 153334
rect 476422 153098 476604 153334
rect 476004 117654 476604 153098
rect 476004 117418 476186 117654
rect 476422 117418 476604 117654
rect 476004 117334 476604 117418
rect 476004 117098 476186 117334
rect 476422 117098 476604 117334
rect 476004 81654 476604 117098
rect 476004 81418 476186 81654
rect 476422 81418 476604 81654
rect 476004 81334 476604 81418
rect 476004 81098 476186 81334
rect 476422 81098 476604 81334
rect 476004 45654 476604 81098
rect 476004 45418 476186 45654
rect 476422 45418 476604 45654
rect 476004 45334 476604 45418
rect 476004 45098 476186 45334
rect 476422 45098 476604 45334
rect 476004 9654 476604 45098
rect 476004 9418 476186 9654
rect 476422 9418 476604 9654
rect 476004 9334 476604 9418
rect 476004 9098 476186 9334
rect 476422 9098 476604 9334
rect 476004 -4106 476604 9098
rect 476004 -4342 476186 -4106
rect 476422 -4342 476604 -4106
rect 476004 -4426 476604 -4342
rect 476004 -4662 476186 -4426
rect 476422 -4662 476604 -4426
rect 476004 -5624 476604 -4662
rect 479604 697254 480204 709922
rect 497604 711418 498204 711440
rect 497604 711182 497786 711418
rect 498022 711182 498204 711418
rect 497604 711098 498204 711182
rect 497604 710862 497786 711098
rect 498022 710862 498204 711098
rect 494004 709538 494604 709560
rect 494004 709302 494186 709538
rect 494422 709302 494604 709538
rect 494004 709218 494604 709302
rect 494004 708982 494186 709218
rect 494422 708982 494604 709218
rect 490404 707658 491004 707680
rect 490404 707422 490586 707658
rect 490822 707422 491004 707658
rect 490404 707338 491004 707422
rect 490404 707102 490586 707338
rect 490822 707102 491004 707338
rect 479604 697018 479786 697254
rect 480022 697018 480204 697254
rect 479604 696934 480204 697018
rect 479604 696698 479786 696934
rect 480022 696698 480204 696934
rect 479604 661254 480204 696698
rect 479604 661018 479786 661254
rect 480022 661018 480204 661254
rect 479604 660934 480204 661018
rect 479604 660698 479786 660934
rect 480022 660698 480204 660934
rect 479604 625254 480204 660698
rect 479604 625018 479786 625254
rect 480022 625018 480204 625254
rect 479604 624934 480204 625018
rect 479604 624698 479786 624934
rect 480022 624698 480204 624934
rect 479604 589254 480204 624698
rect 479604 589018 479786 589254
rect 480022 589018 480204 589254
rect 479604 588934 480204 589018
rect 479604 588698 479786 588934
rect 480022 588698 480204 588934
rect 479604 553254 480204 588698
rect 479604 553018 479786 553254
rect 480022 553018 480204 553254
rect 479604 552934 480204 553018
rect 479604 552698 479786 552934
rect 480022 552698 480204 552934
rect 479604 517254 480204 552698
rect 479604 517018 479786 517254
rect 480022 517018 480204 517254
rect 479604 516934 480204 517018
rect 479604 516698 479786 516934
rect 480022 516698 480204 516934
rect 479604 481254 480204 516698
rect 479604 481018 479786 481254
rect 480022 481018 480204 481254
rect 479604 480934 480204 481018
rect 479604 480698 479786 480934
rect 480022 480698 480204 480934
rect 479604 445254 480204 480698
rect 479604 445018 479786 445254
rect 480022 445018 480204 445254
rect 479604 444934 480204 445018
rect 479604 444698 479786 444934
rect 480022 444698 480204 444934
rect 479604 409254 480204 444698
rect 479604 409018 479786 409254
rect 480022 409018 480204 409254
rect 479604 408934 480204 409018
rect 479604 408698 479786 408934
rect 480022 408698 480204 408934
rect 479604 373254 480204 408698
rect 479604 373018 479786 373254
rect 480022 373018 480204 373254
rect 479604 372934 480204 373018
rect 479604 372698 479786 372934
rect 480022 372698 480204 372934
rect 479604 337254 480204 372698
rect 479604 337018 479786 337254
rect 480022 337018 480204 337254
rect 479604 336934 480204 337018
rect 479604 336698 479786 336934
rect 480022 336698 480204 336934
rect 479604 301254 480204 336698
rect 479604 301018 479786 301254
rect 480022 301018 480204 301254
rect 479604 300934 480204 301018
rect 479604 300698 479786 300934
rect 480022 300698 480204 300934
rect 479604 265254 480204 300698
rect 479604 265018 479786 265254
rect 480022 265018 480204 265254
rect 479604 264934 480204 265018
rect 479604 264698 479786 264934
rect 480022 264698 480204 264934
rect 479604 229254 480204 264698
rect 479604 229018 479786 229254
rect 480022 229018 480204 229254
rect 479604 228934 480204 229018
rect 479604 228698 479786 228934
rect 480022 228698 480204 228934
rect 479604 193254 480204 228698
rect 479604 193018 479786 193254
rect 480022 193018 480204 193254
rect 479604 192934 480204 193018
rect 479604 192698 479786 192934
rect 480022 192698 480204 192934
rect 479604 157254 480204 192698
rect 479604 157018 479786 157254
rect 480022 157018 480204 157254
rect 479604 156934 480204 157018
rect 479604 156698 479786 156934
rect 480022 156698 480204 156934
rect 479604 121254 480204 156698
rect 479604 121018 479786 121254
rect 480022 121018 480204 121254
rect 479604 120934 480204 121018
rect 479604 120698 479786 120934
rect 480022 120698 480204 120934
rect 479604 85254 480204 120698
rect 479604 85018 479786 85254
rect 480022 85018 480204 85254
rect 479604 84934 480204 85018
rect 479604 84698 479786 84934
rect 480022 84698 480204 84934
rect 479604 49254 480204 84698
rect 479604 49018 479786 49254
rect 480022 49018 480204 49254
rect 479604 48934 480204 49018
rect 479604 48698 479786 48934
rect 480022 48698 480204 48934
rect 479604 13254 480204 48698
rect 479604 13018 479786 13254
rect 480022 13018 480204 13254
rect 479604 12934 480204 13018
rect 479604 12698 479786 12934
rect 480022 12698 480204 12934
rect 461604 -7162 461786 -6926
rect 462022 -7162 462204 -6926
rect 461604 -7246 462204 -7162
rect 461604 -7482 461786 -7246
rect 462022 -7482 462204 -7246
rect 461604 -7504 462204 -7482
rect 479604 -5986 480204 12698
rect 486804 705778 487404 705800
rect 486804 705542 486986 705778
rect 487222 705542 487404 705778
rect 486804 705458 487404 705542
rect 486804 705222 486986 705458
rect 487222 705222 487404 705458
rect 486804 668454 487404 705222
rect 486804 668218 486986 668454
rect 487222 668218 487404 668454
rect 486804 668134 487404 668218
rect 486804 667898 486986 668134
rect 487222 667898 487404 668134
rect 486804 632454 487404 667898
rect 486804 632218 486986 632454
rect 487222 632218 487404 632454
rect 486804 632134 487404 632218
rect 486804 631898 486986 632134
rect 487222 631898 487404 632134
rect 486804 596454 487404 631898
rect 486804 596218 486986 596454
rect 487222 596218 487404 596454
rect 486804 596134 487404 596218
rect 486804 595898 486986 596134
rect 487222 595898 487404 596134
rect 486804 560454 487404 595898
rect 486804 560218 486986 560454
rect 487222 560218 487404 560454
rect 486804 560134 487404 560218
rect 486804 559898 486986 560134
rect 487222 559898 487404 560134
rect 486804 524454 487404 559898
rect 486804 524218 486986 524454
rect 487222 524218 487404 524454
rect 486804 524134 487404 524218
rect 486804 523898 486986 524134
rect 487222 523898 487404 524134
rect 486804 488454 487404 523898
rect 486804 488218 486986 488454
rect 487222 488218 487404 488454
rect 486804 488134 487404 488218
rect 486804 487898 486986 488134
rect 487222 487898 487404 488134
rect 486804 452454 487404 487898
rect 486804 452218 486986 452454
rect 487222 452218 487404 452454
rect 486804 452134 487404 452218
rect 486804 451898 486986 452134
rect 487222 451898 487404 452134
rect 486804 416454 487404 451898
rect 486804 416218 486986 416454
rect 487222 416218 487404 416454
rect 486804 416134 487404 416218
rect 486804 415898 486986 416134
rect 487222 415898 487404 416134
rect 486804 380454 487404 415898
rect 486804 380218 486986 380454
rect 487222 380218 487404 380454
rect 486804 380134 487404 380218
rect 486804 379898 486986 380134
rect 487222 379898 487404 380134
rect 486804 344454 487404 379898
rect 486804 344218 486986 344454
rect 487222 344218 487404 344454
rect 486804 344134 487404 344218
rect 486804 343898 486986 344134
rect 487222 343898 487404 344134
rect 486804 308454 487404 343898
rect 486804 308218 486986 308454
rect 487222 308218 487404 308454
rect 486804 308134 487404 308218
rect 486804 307898 486986 308134
rect 487222 307898 487404 308134
rect 486804 272454 487404 307898
rect 486804 272218 486986 272454
rect 487222 272218 487404 272454
rect 486804 272134 487404 272218
rect 486804 271898 486986 272134
rect 487222 271898 487404 272134
rect 486804 236454 487404 271898
rect 486804 236218 486986 236454
rect 487222 236218 487404 236454
rect 486804 236134 487404 236218
rect 486804 235898 486986 236134
rect 487222 235898 487404 236134
rect 486804 200454 487404 235898
rect 486804 200218 486986 200454
rect 487222 200218 487404 200454
rect 486804 200134 487404 200218
rect 486804 199898 486986 200134
rect 487222 199898 487404 200134
rect 486804 164454 487404 199898
rect 486804 164218 486986 164454
rect 487222 164218 487404 164454
rect 486804 164134 487404 164218
rect 486804 163898 486986 164134
rect 487222 163898 487404 164134
rect 486804 128454 487404 163898
rect 486804 128218 486986 128454
rect 487222 128218 487404 128454
rect 486804 128134 487404 128218
rect 486804 127898 486986 128134
rect 487222 127898 487404 128134
rect 486804 92454 487404 127898
rect 486804 92218 486986 92454
rect 487222 92218 487404 92454
rect 486804 92134 487404 92218
rect 486804 91898 486986 92134
rect 487222 91898 487404 92134
rect 486804 56454 487404 91898
rect 486804 56218 486986 56454
rect 487222 56218 487404 56454
rect 486804 56134 487404 56218
rect 486804 55898 486986 56134
rect 487222 55898 487404 56134
rect 486804 20454 487404 55898
rect 486804 20218 486986 20454
rect 487222 20218 487404 20454
rect 486804 20134 487404 20218
rect 486804 19898 486986 20134
rect 487222 19898 487404 20134
rect 486804 -1286 487404 19898
rect 486804 -1522 486986 -1286
rect 487222 -1522 487404 -1286
rect 486804 -1606 487404 -1522
rect 486804 -1842 486986 -1606
rect 487222 -1842 487404 -1606
rect 486804 -1864 487404 -1842
rect 490404 672054 491004 707102
rect 490404 671818 490586 672054
rect 490822 671818 491004 672054
rect 490404 671734 491004 671818
rect 490404 671498 490586 671734
rect 490822 671498 491004 671734
rect 490404 636054 491004 671498
rect 490404 635818 490586 636054
rect 490822 635818 491004 636054
rect 490404 635734 491004 635818
rect 490404 635498 490586 635734
rect 490822 635498 491004 635734
rect 490404 600054 491004 635498
rect 490404 599818 490586 600054
rect 490822 599818 491004 600054
rect 490404 599734 491004 599818
rect 490404 599498 490586 599734
rect 490822 599498 491004 599734
rect 490404 564054 491004 599498
rect 490404 563818 490586 564054
rect 490822 563818 491004 564054
rect 490404 563734 491004 563818
rect 490404 563498 490586 563734
rect 490822 563498 491004 563734
rect 490404 528054 491004 563498
rect 490404 527818 490586 528054
rect 490822 527818 491004 528054
rect 490404 527734 491004 527818
rect 490404 527498 490586 527734
rect 490822 527498 491004 527734
rect 490404 492054 491004 527498
rect 490404 491818 490586 492054
rect 490822 491818 491004 492054
rect 490404 491734 491004 491818
rect 490404 491498 490586 491734
rect 490822 491498 491004 491734
rect 490404 456054 491004 491498
rect 490404 455818 490586 456054
rect 490822 455818 491004 456054
rect 490404 455734 491004 455818
rect 490404 455498 490586 455734
rect 490822 455498 491004 455734
rect 490404 420054 491004 455498
rect 490404 419818 490586 420054
rect 490822 419818 491004 420054
rect 490404 419734 491004 419818
rect 490404 419498 490586 419734
rect 490822 419498 491004 419734
rect 490404 384054 491004 419498
rect 490404 383818 490586 384054
rect 490822 383818 491004 384054
rect 490404 383734 491004 383818
rect 490404 383498 490586 383734
rect 490822 383498 491004 383734
rect 490404 348054 491004 383498
rect 490404 347818 490586 348054
rect 490822 347818 491004 348054
rect 490404 347734 491004 347818
rect 490404 347498 490586 347734
rect 490822 347498 491004 347734
rect 490404 312054 491004 347498
rect 490404 311818 490586 312054
rect 490822 311818 491004 312054
rect 490404 311734 491004 311818
rect 490404 311498 490586 311734
rect 490822 311498 491004 311734
rect 490404 276054 491004 311498
rect 490404 275818 490586 276054
rect 490822 275818 491004 276054
rect 490404 275734 491004 275818
rect 490404 275498 490586 275734
rect 490822 275498 491004 275734
rect 490404 240054 491004 275498
rect 490404 239818 490586 240054
rect 490822 239818 491004 240054
rect 490404 239734 491004 239818
rect 490404 239498 490586 239734
rect 490822 239498 491004 239734
rect 490404 204054 491004 239498
rect 490404 203818 490586 204054
rect 490822 203818 491004 204054
rect 490404 203734 491004 203818
rect 490404 203498 490586 203734
rect 490822 203498 491004 203734
rect 490404 168054 491004 203498
rect 490404 167818 490586 168054
rect 490822 167818 491004 168054
rect 490404 167734 491004 167818
rect 490404 167498 490586 167734
rect 490822 167498 491004 167734
rect 490404 132054 491004 167498
rect 490404 131818 490586 132054
rect 490822 131818 491004 132054
rect 490404 131734 491004 131818
rect 490404 131498 490586 131734
rect 490822 131498 491004 131734
rect 490404 96054 491004 131498
rect 490404 95818 490586 96054
rect 490822 95818 491004 96054
rect 490404 95734 491004 95818
rect 490404 95498 490586 95734
rect 490822 95498 491004 95734
rect 490404 60054 491004 95498
rect 490404 59818 490586 60054
rect 490822 59818 491004 60054
rect 490404 59734 491004 59818
rect 490404 59498 490586 59734
rect 490822 59498 491004 59734
rect 490404 24054 491004 59498
rect 490404 23818 490586 24054
rect 490822 23818 491004 24054
rect 490404 23734 491004 23818
rect 490404 23498 490586 23734
rect 490822 23498 491004 23734
rect 490404 -3166 491004 23498
rect 490404 -3402 490586 -3166
rect 490822 -3402 491004 -3166
rect 490404 -3486 491004 -3402
rect 490404 -3722 490586 -3486
rect 490822 -3722 491004 -3486
rect 490404 -3744 491004 -3722
rect 494004 675654 494604 708982
rect 494004 675418 494186 675654
rect 494422 675418 494604 675654
rect 494004 675334 494604 675418
rect 494004 675098 494186 675334
rect 494422 675098 494604 675334
rect 494004 639654 494604 675098
rect 494004 639418 494186 639654
rect 494422 639418 494604 639654
rect 494004 639334 494604 639418
rect 494004 639098 494186 639334
rect 494422 639098 494604 639334
rect 494004 603654 494604 639098
rect 494004 603418 494186 603654
rect 494422 603418 494604 603654
rect 494004 603334 494604 603418
rect 494004 603098 494186 603334
rect 494422 603098 494604 603334
rect 494004 567654 494604 603098
rect 494004 567418 494186 567654
rect 494422 567418 494604 567654
rect 494004 567334 494604 567418
rect 494004 567098 494186 567334
rect 494422 567098 494604 567334
rect 494004 531654 494604 567098
rect 494004 531418 494186 531654
rect 494422 531418 494604 531654
rect 494004 531334 494604 531418
rect 494004 531098 494186 531334
rect 494422 531098 494604 531334
rect 494004 495654 494604 531098
rect 494004 495418 494186 495654
rect 494422 495418 494604 495654
rect 494004 495334 494604 495418
rect 494004 495098 494186 495334
rect 494422 495098 494604 495334
rect 494004 459654 494604 495098
rect 494004 459418 494186 459654
rect 494422 459418 494604 459654
rect 494004 459334 494604 459418
rect 494004 459098 494186 459334
rect 494422 459098 494604 459334
rect 494004 423654 494604 459098
rect 494004 423418 494186 423654
rect 494422 423418 494604 423654
rect 494004 423334 494604 423418
rect 494004 423098 494186 423334
rect 494422 423098 494604 423334
rect 494004 387654 494604 423098
rect 494004 387418 494186 387654
rect 494422 387418 494604 387654
rect 494004 387334 494604 387418
rect 494004 387098 494186 387334
rect 494422 387098 494604 387334
rect 494004 351654 494604 387098
rect 494004 351418 494186 351654
rect 494422 351418 494604 351654
rect 494004 351334 494604 351418
rect 494004 351098 494186 351334
rect 494422 351098 494604 351334
rect 494004 315654 494604 351098
rect 494004 315418 494186 315654
rect 494422 315418 494604 315654
rect 494004 315334 494604 315418
rect 494004 315098 494186 315334
rect 494422 315098 494604 315334
rect 494004 279654 494604 315098
rect 494004 279418 494186 279654
rect 494422 279418 494604 279654
rect 494004 279334 494604 279418
rect 494004 279098 494186 279334
rect 494422 279098 494604 279334
rect 494004 243654 494604 279098
rect 494004 243418 494186 243654
rect 494422 243418 494604 243654
rect 494004 243334 494604 243418
rect 494004 243098 494186 243334
rect 494422 243098 494604 243334
rect 494004 207654 494604 243098
rect 494004 207418 494186 207654
rect 494422 207418 494604 207654
rect 494004 207334 494604 207418
rect 494004 207098 494186 207334
rect 494422 207098 494604 207334
rect 494004 171654 494604 207098
rect 494004 171418 494186 171654
rect 494422 171418 494604 171654
rect 494004 171334 494604 171418
rect 494004 171098 494186 171334
rect 494422 171098 494604 171334
rect 494004 135654 494604 171098
rect 494004 135418 494186 135654
rect 494422 135418 494604 135654
rect 494004 135334 494604 135418
rect 494004 135098 494186 135334
rect 494422 135098 494604 135334
rect 494004 99654 494604 135098
rect 494004 99418 494186 99654
rect 494422 99418 494604 99654
rect 494004 99334 494604 99418
rect 494004 99098 494186 99334
rect 494422 99098 494604 99334
rect 494004 63654 494604 99098
rect 494004 63418 494186 63654
rect 494422 63418 494604 63654
rect 494004 63334 494604 63418
rect 494004 63098 494186 63334
rect 494422 63098 494604 63334
rect 494004 27654 494604 63098
rect 494004 27418 494186 27654
rect 494422 27418 494604 27654
rect 494004 27334 494604 27418
rect 494004 27098 494186 27334
rect 494422 27098 494604 27334
rect 494004 -5046 494604 27098
rect 494004 -5282 494186 -5046
rect 494422 -5282 494604 -5046
rect 494004 -5366 494604 -5282
rect 494004 -5602 494186 -5366
rect 494422 -5602 494604 -5366
rect 494004 -5624 494604 -5602
rect 497604 679254 498204 710862
rect 515604 710478 516204 711440
rect 515604 710242 515786 710478
rect 516022 710242 516204 710478
rect 515604 710158 516204 710242
rect 515604 709922 515786 710158
rect 516022 709922 516204 710158
rect 512004 708598 512604 709560
rect 512004 708362 512186 708598
rect 512422 708362 512604 708598
rect 512004 708278 512604 708362
rect 512004 708042 512186 708278
rect 512422 708042 512604 708278
rect 508404 706718 509004 707680
rect 508404 706482 508586 706718
rect 508822 706482 509004 706718
rect 508404 706398 509004 706482
rect 508404 706162 508586 706398
rect 508822 706162 509004 706398
rect 497604 679018 497786 679254
rect 498022 679018 498204 679254
rect 497604 678934 498204 679018
rect 497604 678698 497786 678934
rect 498022 678698 498204 678934
rect 497604 643254 498204 678698
rect 497604 643018 497786 643254
rect 498022 643018 498204 643254
rect 497604 642934 498204 643018
rect 497604 642698 497786 642934
rect 498022 642698 498204 642934
rect 497604 607254 498204 642698
rect 497604 607018 497786 607254
rect 498022 607018 498204 607254
rect 497604 606934 498204 607018
rect 497604 606698 497786 606934
rect 498022 606698 498204 606934
rect 497604 571254 498204 606698
rect 497604 571018 497786 571254
rect 498022 571018 498204 571254
rect 497604 570934 498204 571018
rect 497604 570698 497786 570934
rect 498022 570698 498204 570934
rect 497604 535254 498204 570698
rect 497604 535018 497786 535254
rect 498022 535018 498204 535254
rect 497604 534934 498204 535018
rect 497604 534698 497786 534934
rect 498022 534698 498204 534934
rect 497604 499254 498204 534698
rect 497604 499018 497786 499254
rect 498022 499018 498204 499254
rect 497604 498934 498204 499018
rect 497604 498698 497786 498934
rect 498022 498698 498204 498934
rect 497604 463254 498204 498698
rect 497604 463018 497786 463254
rect 498022 463018 498204 463254
rect 497604 462934 498204 463018
rect 497604 462698 497786 462934
rect 498022 462698 498204 462934
rect 497604 427254 498204 462698
rect 497604 427018 497786 427254
rect 498022 427018 498204 427254
rect 497604 426934 498204 427018
rect 497604 426698 497786 426934
rect 498022 426698 498204 426934
rect 497604 391254 498204 426698
rect 497604 391018 497786 391254
rect 498022 391018 498204 391254
rect 497604 390934 498204 391018
rect 497604 390698 497786 390934
rect 498022 390698 498204 390934
rect 497604 355254 498204 390698
rect 497604 355018 497786 355254
rect 498022 355018 498204 355254
rect 497604 354934 498204 355018
rect 497604 354698 497786 354934
rect 498022 354698 498204 354934
rect 497604 319254 498204 354698
rect 497604 319018 497786 319254
rect 498022 319018 498204 319254
rect 497604 318934 498204 319018
rect 497604 318698 497786 318934
rect 498022 318698 498204 318934
rect 497604 283254 498204 318698
rect 497604 283018 497786 283254
rect 498022 283018 498204 283254
rect 497604 282934 498204 283018
rect 497604 282698 497786 282934
rect 498022 282698 498204 282934
rect 497604 247254 498204 282698
rect 497604 247018 497786 247254
rect 498022 247018 498204 247254
rect 497604 246934 498204 247018
rect 497604 246698 497786 246934
rect 498022 246698 498204 246934
rect 497604 211254 498204 246698
rect 497604 211018 497786 211254
rect 498022 211018 498204 211254
rect 497604 210934 498204 211018
rect 497604 210698 497786 210934
rect 498022 210698 498204 210934
rect 497604 175254 498204 210698
rect 497604 175018 497786 175254
rect 498022 175018 498204 175254
rect 497604 174934 498204 175018
rect 497604 174698 497786 174934
rect 498022 174698 498204 174934
rect 497604 139254 498204 174698
rect 497604 139018 497786 139254
rect 498022 139018 498204 139254
rect 497604 138934 498204 139018
rect 497604 138698 497786 138934
rect 498022 138698 498204 138934
rect 497604 103254 498204 138698
rect 497604 103018 497786 103254
rect 498022 103018 498204 103254
rect 497604 102934 498204 103018
rect 497604 102698 497786 102934
rect 498022 102698 498204 102934
rect 497604 67254 498204 102698
rect 497604 67018 497786 67254
rect 498022 67018 498204 67254
rect 497604 66934 498204 67018
rect 497604 66698 497786 66934
rect 498022 66698 498204 66934
rect 497604 31254 498204 66698
rect 497604 31018 497786 31254
rect 498022 31018 498204 31254
rect 497604 30934 498204 31018
rect 497604 30698 497786 30934
rect 498022 30698 498204 30934
rect 479604 -6222 479786 -5986
rect 480022 -6222 480204 -5986
rect 479604 -6306 480204 -6222
rect 479604 -6542 479786 -6306
rect 480022 -6542 480204 -6306
rect 479604 -7504 480204 -6542
rect 497604 -6926 498204 30698
rect 504804 704838 505404 705800
rect 504804 704602 504986 704838
rect 505222 704602 505404 704838
rect 504804 704518 505404 704602
rect 504804 704282 504986 704518
rect 505222 704282 505404 704518
rect 504804 686454 505404 704282
rect 504804 686218 504986 686454
rect 505222 686218 505404 686454
rect 504804 686134 505404 686218
rect 504804 685898 504986 686134
rect 505222 685898 505404 686134
rect 504804 650454 505404 685898
rect 504804 650218 504986 650454
rect 505222 650218 505404 650454
rect 504804 650134 505404 650218
rect 504804 649898 504986 650134
rect 505222 649898 505404 650134
rect 504804 614454 505404 649898
rect 504804 614218 504986 614454
rect 505222 614218 505404 614454
rect 504804 614134 505404 614218
rect 504804 613898 504986 614134
rect 505222 613898 505404 614134
rect 504804 578454 505404 613898
rect 504804 578218 504986 578454
rect 505222 578218 505404 578454
rect 504804 578134 505404 578218
rect 504804 577898 504986 578134
rect 505222 577898 505404 578134
rect 504804 542454 505404 577898
rect 504804 542218 504986 542454
rect 505222 542218 505404 542454
rect 504804 542134 505404 542218
rect 504804 541898 504986 542134
rect 505222 541898 505404 542134
rect 504804 506454 505404 541898
rect 504804 506218 504986 506454
rect 505222 506218 505404 506454
rect 504804 506134 505404 506218
rect 504804 505898 504986 506134
rect 505222 505898 505404 506134
rect 504804 470454 505404 505898
rect 504804 470218 504986 470454
rect 505222 470218 505404 470454
rect 504804 470134 505404 470218
rect 504804 469898 504986 470134
rect 505222 469898 505404 470134
rect 504804 434454 505404 469898
rect 504804 434218 504986 434454
rect 505222 434218 505404 434454
rect 504804 434134 505404 434218
rect 504804 433898 504986 434134
rect 505222 433898 505404 434134
rect 504804 398454 505404 433898
rect 504804 398218 504986 398454
rect 505222 398218 505404 398454
rect 504804 398134 505404 398218
rect 504804 397898 504986 398134
rect 505222 397898 505404 398134
rect 504804 362454 505404 397898
rect 504804 362218 504986 362454
rect 505222 362218 505404 362454
rect 504804 362134 505404 362218
rect 504804 361898 504986 362134
rect 505222 361898 505404 362134
rect 504804 326454 505404 361898
rect 504804 326218 504986 326454
rect 505222 326218 505404 326454
rect 504804 326134 505404 326218
rect 504804 325898 504986 326134
rect 505222 325898 505404 326134
rect 504804 290454 505404 325898
rect 504804 290218 504986 290454
rect 505222 290218 505404 290454
rect 504804 290134 505404 290218
rect 504804 289898 504986 290134
rect 505222 289898 505404 290134
rect 504804 254454 505404 289898
rect 504804 254218 504986 254454
rect 505222 254218 505404 254454
rect 504804 254134 505404 254218
rect 504804 253898 504986 254134
rect 505222 253898 505404 254134
rect 504804 218454 505404 253898
rect 504804 218218 504986 218454
rect 505222 218218 505404 218454
rect 504804 218134 505404 218218
rect 504804 217898 504986 218134
rect 505222 217898 505404 218134
rect 504804 182454 505404 217898
rect 504804 182218 504986 182454
rect 505222 182218 505404 182454
rect 504804 182134 505404 182218
rect 504804 181898 504986 182134
rect 505222 181898 505404 182134
rect 504804 146454 505404 181898
rect 504804 146218 504986 146454
rect 505222 146218 505404 146454
rect 504804 146134 505404 146218
rect 504804 145898 504986 146134
rect 505222 145898 505404 146134
rect 504804 110454 505404 145898
rect 504804 110218 504986 110454
rect 505222 110218 505404 110454
rect 504804 110134 505404 110218
rect 504804 109898 504986 110134
rect 505222 109898 505404 110134
rect 504804 74454 505404 109898
rect 504804 74218 504986 74454
rect 505222 74218 505404 74454
rect 504804 74134 505404 74218
rect 504804 73898 504986 74134
rect 505222 73898 505404 74134
rect 504804 38454 505404 73898
rect 504804 38218 504986 38454
rect 505222 38218 505404 38454
rect 504804 38134 505404 38218
rect 504804 37898 504986 38134
rect 505222 37898 505404 38134
rect 504804 2454 505404 37898
rect 504804 2218 504986 2454
rect 505222 2218 505404 2454
rect 504804 2134 505404 2218
rect 504804 1898 504986 2134
rect 505222 1898 505404 2134
rect 504804 -346 505404 1898
rect 504804 -582 504986 -346
rect 505222 -582 505404 -346
rect 504804 -666 505404 -582
rect 504804 -902 504986 -666
rect 505222 -902 505404 -666
rect 504804 -1864 505404 -902
rect 508404 690054 509004 706162
rect 508404 689818 508586 690054
rect 508822 689818 509004 690054
rect 508404 689734 509004 689818
rect 508404 689498 508586 689734
rect 508822 689498 509004 689734
rect 508404 654054 509004 689498
rect 508404 653818 508586 654054
rect 508822 653818 509004 654054
rect 508404 653734 509004 653818
rect 508404 653498 508586 653734
rect 508822 653498 509004 653734
rect 508404 618054 509004 653498
rect 508404 617818 508586 618054
rect 508822 617818 509004 618054
rect 508404 617734 509004 617818
rect 508404 617498 508586 617734
rect 508822 617498 509004 617734
rect 508404 582054 509004 617498
rect 508404 581818 508586 582054
rect 508822 581818 509004 582054
rect 508404 581734 509004 581818
rect 508404 581498 508586 581734
rect 508822 581498 509004 581734
rect 508404 546054 509004 581498
rect 508404 545818 508586 546054
rect 508822 545818 509004 546054
rect 508404 545734 509004 545818
rect 508404 545498 508586 545734
rect 508822 545498 509004 545734
rect 508404 510054 509004 545498
rect 508404 509818 508586 510054
rect 508822 509818 509004 510054
rect 508404 509734 509004 509818
rect 508404 509498 508586 509734
rect 508822 509498 509004 509734
rect 508404 474054 509004 509498
rect 508404 473818 508586 474054
rect 508822 473818 509004 474054
rect 508404 473734 509004 473818
rect 508404 473498 508586 473734
rect 508822 473498 509004 473734
rect 508404 438054 509004 473498
rect 508404 437818 508586 438054
rect 508822 437818 509004 438054
rect 508404 437734 509004 437818
rect 508404 437498 508586 437734
rect 508822 437498 509004 437734
rect 508404 402054 509004 437498
rect 508404 401818 508586 402054
rect 508822 401818 509004 402054
rect 508404 401734 509004 401818
rect 508404 401498 508586 401734
rect 508822 401498 509004 401734
rect 508404 366054 509004 401498
rect 508404 365818 508586 366054
rect 508822 365818 509004 366054
rect 508404 365734 509004 365818
rect 508404 365498 508586 365734
rect 508822 365498 509004 365734
rect 508404 330054 509004 365498
rect 508404 329818 508586 330054
rect 508822 329818 509004 330054
rect 508404 329734 509004 329818
rect 508404 329498 508586 329734
rect 508822 329498 509004 329734
rect 508404 294054 509004 329498
rect 508404 293818 508586 294054
rect 508822 293818 509004 294054
rect 508404 293734 509004 293818
rect 508404 293498 508586 293734
rect 508822 293498 509004 293734
rect 508404 258054 509004 293498
rect 508404 257818 508586 258054
rect 508822 257818 509004 258054
rect 508404 257734 509004 257818
rect 508404 257498 508586 257734
rect 508822 257498 509004 257734
rect 508404 222054 509004 257498
rect 508404 221818 508586 222054
rect 508822 221818 509004 222054
rect 508404 221734 509004 221818
rect 508404 221498 508586 221734
rect 508822 221498 509004 221734
rect 508404 186054 509004 221498
rect 508404 185818 508586 186054
rect 508822 185818 509004 186054
rect 508404 185734 509004 185818
rect 508404 185498 508586 185734
rect 508822 185498 509004 185734
rect 508404 150054 509004 185498
rect 508404 149818 508586 150054
rect 508822 149818 509004 150054
rect 508404 149734 509004 149818
rect 508404 149498 508586 149734
rect 508822 149498 509004 149734
rect 508404 114054 509004 149498
rect 508404 113818 508586 114054
rect 508822 113818 509004 114054
rect 508404 113734 509004 113818
rect 508404 113498 508586 113734
rect 508822 113498 509004 113734
rect 508404 78054 509004 113498
rect 508404 77818 508586 78054
rect 508822 77818 509004 78054
rect 508404 77734 509004 77818
rect 508404 77498 508586 77734
rect 508822 77498 509004 77734
rect 508404 42054 509004 77498
rect 508404 41818 508586 42054
rect 508822 41818 509004 42054
rect 508404 41734 509004 41818
rect 508404 41498 508586 41734
rect 508822 41498 509004 41734
rect 508404 6054 509004 41498
rect 508404 5818 508586 6054
rect 508822 5818 509004 6054
rect 508404 5734 509004 5818
rect 508404 5498 508586 5734
rect 508822 5498 509004 5734
rect 508404 -2226 509004 5498
rect 508404 -2462 508586 -2226
rect 508822 -2462 509004 -2226
rect 508404 -2546 509004 -2462
rect 508404 -2782 508586 -2546
rect 508822 -2782 509004 -2546
rect 508404 -3744 509004 -2782
rect 512004 693654 512604 708042
rect 512004 693418 512186 693654
rect 512422 693418 512604 693654
rect 512004 693334 512604 693418
rect 512004 693098 512186 693334
rect 512422 693098 512604 693334
rect 512004 657654 512604 693098
rect 512004 657418 512186 657654
rect 512422 657418 512604 657654
rect 512004 657334 512604 657418
rect 512004 657098 512186 657334
rect 512422 657098 512604 657334
rect 512004 621654 512604 657098
rect 512004 621418 512186 621654
rect 512422 621418 512604 621654
rect 512004 621334 512604 621418
rect 512004 621098 512186 621334
rect 512422 621098 512604 621334
rect 512004 585654 512604 621098
rect 512004 585418 512186 585654
rect 512422 585418 512604 585654
rect 512004 585334 512604 585418
rect 512004 585098 512186 585334
rect 512422 585098 512604 585334
rect 512004 549654 512604 585098
rect 512004 549418 512186 549654
rect 512422 549418 512604 549654
rect 512004 549334 512604 549418
rect 512004 549098 512186 549334
rect 512422 549098 512604 549334
rect 512004 513654 512604 549098
rect 512004 513418 512186 513654
rect 512422 513418 512604 513654
rect 512004 513334 512604 513418
rect 512004 513098 512186 513334
rect 512422 513098 512604 513334
rect 512004 477654 512604 513098
rect 512004 477418 512186 477654
rect 512422 477418 512604 477654
rect 512004 477334 512604 477418
rect 512004 477098 512186 477334
rect 512422 477098 512604 477334
rect 512004 441654 512604 477098
rect 512004 441418 512186 441654
rect 512422 441418 512604 441654
rect 512004 441334 512604 441418
rect 512004 441098 512186 441334
rect 512422 441098 512604 441334
rect 512004 405654 512604 441098
rect 512004 405418 512186 405654
rect 512422 405418 512604 405654
rect 512004 405334 512604 405418
rect 512004 405098 512186 405334
rect 512422 405098 512604 405334
rect 512004 369654 512604 405098
rect 512004 369418 512186 369654
rect 512422 369418 512604 369654
rect 512004 369334 512604 369418
rect 512004 369098 512186 369334
rect 512422 369098 512604 369334
rect 512004 333654 512604 369098
rect 512004 333418 512186 333654
rect 512422 333418 512604 333654
rect 512004 333334 512604 333418
rect 512004 333098 512186 333334
rect 512422 333098 512604 333334
rect 512004 297654 512604 333098
rect 512004 297418 512186 297654
rect 512422 297418 512604 297654
rect 512004 297334 512604 297418
rect 512004 297098 512186 297334
rect 512422 297098 512604 297334
rect 512004 261654 512604 297098
rect 512004 261418 512186 261654
rect 512422 261418 512604 261654
rect 512004 261334 512604 261418
rect 512004 261098 512186 261334
rect 512422 261098 512604 261334
rect 512004 225654 512604 261098
rect 512004 225418 512186 225654
rect 512422 225418 512604 225654
rect 512004 225334 512604 225418
rect 512004 225098 512186 225334
rect 512422 225098 512604 225334
rect 512004 189654 512604 225098
rect 512004 189418 512186 189654
rect 512422 189418 512604 189654
rect 512004 189334 512604 189418
rect 512004 189098 512186 189334
rect 512422 189098 512604 189334
rect 512004 153654 512604 189098
rect 512004 153418 512186 153654
rect 512422 153418 512604 153654
rect 512004 153334 512604 153418
rect 512004 153098 512186 153334
rect 512422 153098 512604 153334
rect 512004 117654 512604 153098
rect 512004 117418 512186 117654
rect 512422 117418 512604 117654
rect 512004 117334 512604 117418
rect 512004 117098 512186 117334
rect 512422 117098 512604 117334
rect 512004 81654 512604 117098
rect 512004 81418 512186 81654
rect 512422 81418 512604 81654
rect 512004 81334 512604 81418
rect 512004 81098 512186 81334
rect 512422 81098 512604 81334
rect 512004 45654 512604 81098
rect 512004 45418 512186 45654
rect 512422 45418 512604 45654
rect 512004 45334 512604 45418
rect 512004 45098 512186 45334
rect 512422 45098 512604 45334
rect 512004 9654 512604 45098
rect 512004 9418 512186 9654
rect 512422 9418 512604 9654
rect 512004 9334 512604 9418
rect 512004 9098 512186 9334
rect 512422 9098 512604 9334
rect 512004 -4106 512604 9098
rect 512004 -4342 512186 -4106
rect 512422 -4342 512604 -4106
rect 512004 -4426 512604 -4342
rect 512004 -4662 512186 -4426
rect 512422 -4662 512604 -4426
rect 512004 -5624 512604 -4662
rect 515604 697254 516204 709922
rect 533604 711418 534204 711440
rect 533604 711182 533786 711418
rect 534022 711182 534204 711418
rect 533604 711098 534204 711182
rect 533604 710862 533786 711098
rect 534022 710862 534204 711098
rect 530004 709538 530604 709560
rect 530004 709302 530186 709538
rect 530422 709302 530604 709538
rect 530004 709218 530604 709302
rect 530004 708982 530186 709218
rect 530422 708982 530604 709218
rect 526404 707658 527004 707680
rect 526404 707422 526586 707658
rect 526822 707422 527004 707658
rect 526404 707338 527004 707422
rect 526404 707102 526586 707338
rect 526822 707102 527004 707338
rect 515604 697018 515786 697254
rect 516022 697018 516204 697254
rect 515604 696934 516204 697018
rect 515604 696698 515786 696934
rect 516022 696698 516204 696934
rect 515604 661254 516204 696698
rect 515604 661018 515786 661254
rect 516022 661018 516204 661254
rect 515604 660934 516204 661018
rect 515604 660698 515786 660934
rect 516022 660698 516204 660934
rect 515604 625254 516204 660698
rect 515604 625018 515786 625254
rect 516022 625018 516204 625254
rect 515604 624934 516204 625018
rect 515604 624698 515786 624934
rect 516022 624698 516204 624934
rect 515604 589254 516204 624698
rect 515604 589018 515786 589254
rect 516022 589018 516204 589254
rect 515604 588934 516204 589018
rect 515604 588698 515786 588934
rect 516022 588698 516204 588934
rect 515604 553254 516204 588698
rect 515604 553018 515786 553254
rect 516022 553018 516204 553254
rect 515604 552934 516204 553018
rect 515604 552698 515786 552934
rect 516022 552698 516204 552934
rect 515604 517254 516204 552698
rect 515604 517018 515786 517254
rect 516022 517018 516204 517254
rect 515604 516934 516204 517018
rect 515604 516698 515786 516934
rect 516022 516698 516204 516934
rect 515604 481254 516204 516698
rect 515604 481018 515786 481254
rect 516022 481018 516204 481254
rect 515604 480934 516204 481018
rect 515604 480698 515786 480934
rect 516022 480698 516204 480934
rect 515604 445254 516204 480698
rect 515604 445018 515786 445254
rect 516022 445018 516204 445254
rect 515604 444934 516204 445018
rect 515604 444698 515786 444934
rect 516022 444698 516204 444934
rect 515604 409254 516204 444698
rect 515604 409018 515786 409254
rect 516022 409018 516204 409254
rect 515604 408934 516204 409018
rect 515604 408698 515786 408934
rect 516022 408698 516204 408934
rect 515604 373254 516204 408698
rect 515604 373018 515786 373254
rect 516022 373018 516204 373254
rect 515604 372934 516204 373018
rect 515604 372698 515786 372934
rect 516022 372698 516204 372934
rect 515604 337254 516204 372698
rect 515604 337018 515786 337254
rect 516022 337018 516204 337254
rect 515604 336934 516204 337018
rect 515604 336698 515786 336934
rect 516022 336698 516204 336934
rect 515604 301254 516204 336698
rect 515604 301018 515786 301254
rect 516022 301018 516204 301254
rect 515604 300934 516204 301018
rect 515604 300698 515786 300934
rect 516022 300698 516204 300934
rect 515604 265254 516204 300698
rect 515604 265018 515786 265254
rect 516022 265018 516204 265254
rect 515604 264934 516204 265018
rect 515604 264698 515786 264934
rect 516022 264698 516204 264934
rect 515604 229254 516204 264698
rect 515604 229018 515786 229254
rect 516022 229018 516204 229254
rect 515604 228934 516204 229018
rect 515604 228698 515786 228934
rect 516022 228698 516204 228934
rect 515604 193254 516204 228698
rect 515604 193018 515786 193254
rect 516022 193018 516204 193254
rect 515604 192934 516204 193018
rect 515604 192698 515786 192934
rect 516022 192698 516204 192934
rect 515604 157254 516204 192698
rect 515604 157018 515786 157254
rect 516022 157018 516204 157254
rect 515604 156934 516204 157018
rect 515604 156698 515786 156934
rect 516022 156698 516204 156934
rect 515604 121254 516204 156698
rect 515604 121018 515786 121254
rect 516022 121018 516204 121254
rect 515604 120934 516204 121018
rect 515604 120698 515786 120934
rect 516022 120698 516204 120934
rect 515604 85254 516204 120698
rect 515604 85018 515786 85254
rect 516022 85018 516204 85254
rect 515604 84934 516204 85018
rect 515604 84698 515786 84934
rect 516022 84698 516204 84934
rect 515604 49254 516204 84698
rect 515604 49018 515786 49254
rect 516022 49018 516204 49254
rect 515604 48934 516204 49018
rect 515604 48698 515786 48934
rect 516022 48698 516204 48934
rect 515604 13254 516204 48698
rect 515604 13018 515786 13254
rect 516022 13018 516204 13254
rect 515604 12934 516204 13018
rect 515604 12698 515786 12934
rect 516022 12698 516204 12934
rect 497604 -7162 497786 -6926
rect 498022 -7162 498204 -6926
rect 497604 -7246 498204 -7162
rect 497604 -7482 497786 -7246
rect 498022 -7482 498204 -7246
rect 497604 -7504 498204 -7482
rect 515604 -5986 516204 12698
rect 522804 705778 523404 705800
rect 522804 705542 522986 705778
rect 523222 705542 523404 705778
rect 522804 705458 523404 705542
rect 522804 705222 522986 705458
rect 523222 705222 523404 705458
rect 522804 668454 523404 705222
rect 522804 668218 522986 668454
rect 523222 668218 523404 668454
rect 522804 668134 523404 668218
rect 522804 667898 522986 668134
rect 523222 667898 523404 668134
rect 522804 632454 523404 667898
rect 522804 632218 522986 632454
rect 523222 632218 523404 632454
rect 522804 632134 523404 632218
rect 522804 631898 522986 632134
rect 523222 631898 523404 632134
rect 522804 596454 523404 631898
rect 522804 596218 522986 596454
rect 523222 596218 523404 596454
rect 522804 596134 523404 596218
rect 522804 595898 522986 596134
rect 523222 595898 523404 596134
rect 522804 560454 523404 595898
rect 522804 560218 522986 560454
rect 523222 560218 523404 560454
rect 522804 560134 523404 560218
rect 522804 559898 522986 560134
rect 523222 559898 523404 560134
rect 522804 524454 523404 559898
rect 522804 524218 522986 524454
rect 523222 524218 523404 524454
rect 522804 524134 523404 524218
rect 522804 523898 522986 524134
rect 523222 523898 523404 524134
rect 522804 488454 523404 523898
rect 522804 488218 522986 488454
rect 523222 488218 523404 488454
rect 522804 488134 523404 488218
rect 522804 487898 522986 488134
rect 523222 487898 523404 488134
rect 522804 452454 523404 487898
rect 522804 452218 522986 452454
rect 523222 452218 523404 452454
rect 522804 452134 523404 452218
rect 522804 451898 522986 452134
rect 523222 451898 523404 452134
rect 522804 416454 523404 451898
rect 522804 416218 522986 416454
rect 523222 416218 523404 416454
rect 522804 416134 523404 416218
rect 522804 415898 522986 416134
rect 523222 415898 523404 416134
rect 522804 380454 523404 415898
rect 522804 380218 522986 380454
rect 523222 380218 523404 380454
rect 522804 380134 523404 380218
rect 522804 379898 522986 380134
rect 523222 379898 523404 380134
rect 522804 344454 523404 379898
rect 522804 344218 522986 344454
rect 523222 344218 523404 344454
rect 522804 344134 523404 344218
rect 522804 343898 522986 344134
rect 523222 343898 523404 344134
rect 522804 308454 523404 343898
rect 522804 308218 522986 308454
rect 523222 308218 523404 308454
rect 522804 308134 523404 308218
rect 522804 307898 522986 308134
rect 523222 307898 523404 308134
rect 522804 272454 523404 307898
rect 522804 272218 522986 272454
rect 523222 272218 523404 272454
rect 522804 272134 523404 272218
rect 522804 271898 522986 272134
rect 523222 271898 523404 272134
rect 522804 236454 523404 271898
rect 522804 236218 522986 236454
rect 523222 236218 523404 236454
rect 522804 236134 523404 236218
rect 522804 235898 522986 236134
rect 523222 235898 523404 236134
rect 522804 200454 523404 235898
rect 522804 200218 522986 200454
rect 523222 200218 523404 200454
rect 522804 200134 523404 200218
rect 522804 199898 522986 200134
rect 523222 199898 523404 200134
rect 522804 164454 523404 199898
rect 522804 164218 522986 164454
rect 523222 164218 523404 164454
rect 522804 164134 523404 164218
rect 522804 163898 522986 164134
rect 523222 163898 523404 164134
rect 522804 128454 523404 163898
rect 522804 128218 522986 128454
rect 523222 128218 523404 128454
rect 522804 128134 523404 128218
rect 522804 127898 522986 128134
rect 523222 127898 523404 128134
rect 522804 92454 523404 127898
rect 522804 92218 522986 92454
rect 523222 92218 523404 92454
rect 522804 92134 523404 92218
rect 522804 91898 522986 92134
rect 523222 91898 523404 92134
rect 522804 56454 523404 91898
rect 522804 56218 522986 56454
rect 523222 56218 523404 56454
rect 522804 56134 523404 56218
rect 522804 55898 522986 56134
rect 523222 55898 523404 56134
rect 522804 20454 523404 55898
rect 522804 20218 522986 20454
rect 523222 20218 523404 20454
rect 522804 20134 523404 20218
rect 522804 19898 522986 20134
rect 523222 19898 523404 20134
rect 522804 -1286 523404 19898
rect 522804 -1522 522986 -1286
rect 523222 -1522 523404 -1286
rect 522804 -1606 523404 -1522
rect 522804 -1842 522986 -1606
rect 523222 -1842 523404 -1606
rect 522804 -1864 523404 -1842
rect 526404 672054 527004 707102
rect 526404 671818 526586 672054
rect 526822 671818 527004 672054
rect 526404 671734 527004 671818
rect 526404 671498 526586 671734
rect 526822 671498 527004 671734
rect 526404 636054 527004 671498
rect 526404 635818 526586 636054
rect 526822 635818 527004 636054
rect 526404 635734 527004 635818
rect 526404 635498 526586 635734
rect 526822 635498 527004 635734
rect 526404 600054 527004 635498
rect 526404 599818 526586 600054
rect 526822 599818 527004 600054
rect 526404 599734 527004 599818
rect 526404 599498 526586 599734
rect 526822 599498 527004 599734
rect 526404 564054 527004 599498
rect 526404 563818 526586 564054
rect 526822 563818 527004 564054
rect 526404 563734 527004 563818
rect 526404 563498 526586 563734
rect 526822 563498 527004 563734
rect 526404 528054 527004 563498
rect 526404 527818 526586 528054
rect 526822 527818 527004 528054
rect 526404 527734 527004 527818
rect 526404 527498 526586 527734
rect 526822 527498 527004 527734
rect 526404 492054 527004 527498
rect 526404 491818 526586 492054
rect 526822 491818 527004 492054
rect 526404 491734 527004 491818
rect 526404 491498 526586 491734
rect 526822 491498 527004 491734
rect 526404 456054 527004 491498
rect 526404 455818 526586 456054
rect 526822 455818 527004 456054
rect 526404 455734 527004 455818
rect 526404 455498 526586 455734
rect 526822 455498 527004 455734
rect 526404 420054 527004 455498
rect 526404 419818 526586 420054
rect 526822 419818 527004 420054
rect 526404 419734 527004 419818
rect 526404 419498 526586 419734
rect 526822 419498 527004 419734
rect 526404 384054 527004 419498
rect 526404 383818 526586 384054
rect 526822 383818 527004 384054
rect 526404 383734 527004 383818
rect 526404 383498 526586 383734
rect 526822 383498 527004 383734
rect 526404 348054 527004 383498
rect 526404 347818 526586 348054
rect 526822 347818 527004 348054
rect 526404 347734 527004 347818
rect 526404 347498 526586 347734
rect 526822 347498 527004 347734
rect 526404 312054 527004 347498
rect 526404 311818 526586 312054
rect 526822 311818 527004 312054
rect 526404 311734 527004 311818
rect 526404 311498 526586 311734
rect 526822 311498 527004 311734
rect 526404 276054 527004 311498
rect 526404 275818 526586 276054
rect 526822 275818 527004 276054
rect 526404 275734 527004 275818
rect 526404 275498 526586 275734
rect 526822 275498 527004 275734
rect 526404 240054 527004 275498
rect 526404 239818 526586 240054
rect 526822 239818 527004 240054
rect 526404 239734 527004 239818
rect 526404 239498 526586 239734
rect 526822 239498 527004 239734
rect 526404 204054 527004 239498
rect 526404 203818 526586 204054
rect 526822 203818 527004 204054
rect 526404 203734 527004 203818
rect 526404 203498 526586 203734
rect 526822 203498 527004 203734
rect 526404 168054 527004 203498
rect 526404 167818 526586 168054
rect 526822 167818 527004 168054
rect 526404 167734 527004 167818
rect 526404 167498 526586 167734
rect 526822 167498 527004 167734
rect 526404 132054 527004 167498
rect 526404 131818 526586 132054
rect 526822 131818 527004 132054
rect 526404 131734 527004 131818
rect 526404 131498 526586 131734
rect 526822 131498 527004 131734
rect 526404 96054 527004 131498
rect 526404 95818 526586 96054
rect 526822 95818 527004 96054
rect 526404 95734 527004 95818
rect 526404 95498 526586 95734
rect 526822 95498 527004 95734
rect 526404 60054 527004 95498
rect 526404 59818 526586 60054
rect 526822 59818 527004 60054
rect 526404 59734 527004 59818
rect 526404 59498 526586 59734
rect 526822 59498 527004 59734
rect 526404 24054 527004 59498
rect 526404 23818 526586 24054
rect 526822 23818 527004 24054
rect 526404 23734 527004 23818
rect 526404 23498 526586 23734
rect 526822 23498 527004 23734
rect 526404 -3166 527004 23498
rect 526404 -3402 526586 -3166
rect 526822 -3402 527004 -3166
rect 526404 -3486 527004 -3402
rect 526404 -3722 526586 -3486
rect 526822 -3722 527004 -3486
rect 526404 -3744 527004 -3722
rect 530004 675654 530604 708982
rect 530004 675418 530186 675654
rect 530422 675418 530604 675654
rect 530004 675334 530604 675418
rect 530004 675098 530186 675334
rect 530422 675098 530604 675334
rect 530004 639654 530604 675098
rect 530004 639418 530186 639654
rect 530422 639418 530604 639654
rect 530004 639334 530604 639418
rect 530004 639098 530186 639334
rect 530422 639098 530604 639334
rect 530004 603654 530604 639098
rect 530004 603418 530186 603654
rect 530422 603418 530604 603654
rect 530004 603334 530604 603418
rect 530004 603098 530186 603334
rect 530422 603098 530604 603334
rect 530004 567654 530604 603098
rect 530004 567418 530186 567654
rect 530422 567418 530604 567654
rect 530004 567334 530604 567418
rect 530004 567098 530186 567334
rect 530422 567098 530604 567334
rect 530004 531654 530604 567098
rect 530004 531418 530186 531654
rect 530422 531418 530604 531654
rect 530004 531334 530604 531418
rect 530004 531098 530186 531334
rect 530422 531098 530604 531334
rect 530004 495654 530604 531098
rect 530004 495418 530186 495654
rect 530422 495418 530604 495654
rect 530004 495334 530604 495418
rect 530004 495098 530186 495334
rect 530422 495098 530604 495334
rect 530004 459654 530604 495098
rect 530004 459418 530186 459654
rect 530422 459418 530604 459654
rect 530004 459334 530604 459418
rect 530004 459098 530186 459334
rect 530422 459098 530604 459334
rect 530004 423654 530604 459098
rect 530004 423418 530186 423654
rect 530422 423418 530604 423654
rect 530004 423334 530604 423418
rect 530004 423098 530186 423334
rect 530422 423098 530604 423334
rect 530004 387654 530604 423098
rect 530004 387418 530186 387654
rect 530422 387418 530604 387654
rect 530004 387334 530604 387418
rect 530004 387098 530186 387334
rect 530422 387098 530604 387334
rect 530004 351654 530604 387098
rect 530004 351418 530186 351654
rect 530422 351418 530604 351654
rect 530004 351334 530604 351418
rect 530004 351098 530186 351334
rect 530422 351098 530604 351334
rect 530004 315654 530604 351098
rect 530004 315418 530186 315654
rect 530422 315418 530604 315654
rect 530004 315334 530604 315418
rect 530004 315098 530186 315334
rect 530422 315098 530604 315334
rect 530004 279654 530604 315098
rect 530004 279418 530186 279654
rect 530422 279418 530604 279654
rect 530004 279334 530604 279418
rect 530004 279098 530186 279334
rect 530422 279098 530604 279334
rect 530004 243654 530604 279098
rect 530004 243418 530186 243654
rect 530422 243418 530604 243654
rect 530004 243334 530604 243418
rect 530004 243098 530186 243334
rect 530422 243098 530604 243334
rect 530004 207654 530604 243098
rect 530004 207418 530186 207654
rect 530422 207418 530604 207654
rect 530004 207334 530604 207418
rect 530004 207098 530186 207334
rect 530422 207098 530604 207334
rect 530004 171654 530604 207098
rect 530004 171418 530186 171654
rect 530422 171418 530604 171654
rect 530004 171334 530604 171418
rect 530004 171098 530186 171334
rect 530422 171098 530604 171334
rect 530004 135654 530604 171098
rect 530004 135418 530186 135654
rect 530422 135418 530604 135654
rect 530004 135334 530604 135418
rect 530004 135098 530186 135334
rect 530422 135098 530604 135334
rect 530004 99654 530604 135098
rect 530004 99418 530186 99654
rect 530422 99418 530604 99654
rect 530004 99334 530604 99418
rect 530004 99098 530186 99334
rect 530422 99098 530604 99334
rect 530004 63654 530604 99098
rect 530004 63418 530186 63654
rect 530422 63418 530604 63654
rect 530004 63334 530604 63418
rect 530004 63098 530186 63334
rect 530422 63098 530604 63334
rect 530004 27654 530604 63098
rect 530004 27418 530186 27654
rect 530422 27418 530604 27654
rect 530004 27334 530604 27418
rect 530004 27098 530186 27334
rect 530422 27098 530604 27334
rect 530004 -5046 530604 27098
rect 530004 -5282 530186 -5046
rect 530422 -5282 530604 -5046
rect 530004 -5366 530604 -5282
rect 530004 -5602 530186 -5366
rect 530422 -5602 530604 -5366
rect 530004 -5624 530604 -5602
rect 533604 679254 534204 710862
rect 551604 710478 552204 711440
rect 551604 710242 551786 710478
rect 552022 710242 552204 710478
rect 551604 710158 552204 710242
rect 551604 709922 551786 710158
rect 552022 709922 552204 710158
rect 548004 708598 548604 709560
rect 548004 708362 548186 708598
rect 548422 708362 548604 708598
rect 548004 708278 548604 708362
rect 548004 708042 548186 708278
rect 548422 708042 548604 708278
rect 544404 706718 545004 707680
rect 544404 706482 544586 706718
rect 544822 706482 545004 706718
rect 544404 706398 545004 706482
rect 544404 706162 544586 706398
rect 544822 706162 545004 706398
rect 533604 679018 533786 679254
rect 534022 679018 534204 679254
rect 533604 678934 534204 679018
rect 533604 678698 533786 678934
rect 534022 678698 534204 678934
rect 533604 643254 534204 678698
rect 533604 643018 533786 643254
rect 534022 643018 534204 643254
rect 533604 642934 534204 643018
rect 533604 642698 533786 642934
rect 534022 642698 534204 642934
rect 533604 607254 534204 642698
rect 533604 607018 533786 607254
rect 534022 607018 534204 607254
rect 533604 606934 534204 607018
rect 533604 606698 533786 606934
rect 534022 606698 534204 606934
rect 533604 571254 534204 606698
rect 533604 571018 533786 571254
rect 534022 571018 534204 571254
rect 533604 570934 534204 571018
rect 533604 570698 533786 570934
rect 534022 570698 534204 570934
rect 533604 535254 534204 570698
rect 533604 535018 533786 535254
rect 534022 535018 534204 535254
rect 533604 534934 534204 535018
rect 533604 534698 533786 534934
rect 534022 534698 534204 534934
rect 533604 499254 534204 534698
rect 533604 499018 533786 499254
rect 534022 499018 534204 499254
rect 533604 498934 534204 499018
rect 533604 498698 533786 498934
rect 534022 498698 534204 498934
rect 533604 463254 534204 498698
rect 533604 463018 533786 463254
rect 534022 463018 534204 463254
rect 533604 462934 534204 463018
rect 533604 462698 533786 462934
rect 534022 462698 534204 462934
rect 533604 427254 534204 462698
rect 533604 427018 533786 427254
rect 534022 427018 534204 427254
rect 533604 426934 534204 427018
rect 533604 426698 533786 426934
rect 534022 426698 534204 426934
rect 533604 391254 534204 426698
rect 533604 391018 533786 391254
rect 534022 391018 534204 391254
rect 533604 390934 534204 391018
rect 533604 390698 533786 390934
rect 534022 390698 534204 390934
rect 533604 355254 534204 390698
rect 533604 355018 533786 355254
rect 534022 355018 534204 355254
rect 533604 354934 534204 355018
rect 533604 354698 533786 354934
rect 534022 354698 534204 354934
rect 533604 319254 534204 354698
rect 533604 319018 533786 319254
rect 534022 319018 534204 319254
rect 533604 318934 534204 319018
rect 533604 318698 533786 318934
rect 534022 318698 534204 318934
rect 533604 283254 534204 318698
rect 533604 283018 533786 283254
rect 534022 283018 534204 283254
rect 533604 282934 534204 283018
rect 533604 282698 533786 282934
rect 534022 282698 534204 282934
rect 533604 247254 534204 282698
rect 533604 247018 533786 247254
rect 534022 247018 534204 247254
rect 533604 246934 534204 247018
rect 533604 246698 533786 246934
rect 534022 246698 534204 246934
rect 533604 211254 534204 246698
rect 533604 211018 533786 211254
rect 534022 211018 534204 211254
rect 533604 210934 534204 211018
rect 533604 210698 533786 210934
rect 534022 210698 534204 210934
rect 533604 175254 534204 210698
rect 533604 175018 533786 175254
rect 534022 175018 534204 175254
rect 533604 174934 534204 175018
rect 533604 174698 533786 174934
rect 534022 174698 534204 174934
rect 533604 139254 534204 174698
rect 533604 139018 533786 139254
rect 534022 139018 534204 139254
rect 533604 138934 534204 139018
rect 533604 138698 533786 138934
rect 534022 138698 534204 138934
rect 533604 103254 534204 138698
rect 533604 103018 533786 103254
rect 534022 103018 534204 103254
rect 533604 102934 534204 103018
rect 533604 102698 533786 102934
rect 534022 102698 534204 102934
rect 533604 67254 534204 102698
rect 533604 67018 533786 67254
rect 534022 67018 534204 67254
rect 533604 66934 534204 67018
rect 533604 66698 533786 66934
rect 534022 66698 534204 66934
rect 533604 31254 534204 66698
rect 533604 31018 533786 31254
rect 534022 31018 534204 31254
rect 533604 30934 534204 31018
rect 533604 30698 533786 30934
rect 534022 30698 534204 30934
rect 515604 -6222 515786 -5986
rect 516022 -6222 516204 -5986
rect 515604 -6306 516204 -6222
rect 515604 -6542 515786 -6306
rect 516022 -6542 516204 -6306
rect 515604 -7504 516204 -6542
rect 533604 -6926 534204 30698
rect 540804 704838 541404 705800
rect 540804 704602 540986 704838
rect 541222 704602 541404 704838
rect 540804 704518 541404 704602
rect 540804 704282 540986 704518
rect 541222 704282 541404 704518
rect 540804 686454 541404 704282
rect 540804 686218 540986 686454
rect 541222 686218 541404 686454
rect 540804 686134 541404 686218
rect 540804 685898 540986 686134
rect 541222 685898 541404 686134
rect 540804 650454 541404 685898
rect 540804 650218 540986 650454
rect 541222 650218 541404 650454
rect 540804 650134 541404 650218
rect 540804 649898 540986 650134
rect 541222 649898 541404 650134
rect 540804 614454 541404 649898
rect 540804 614218 540986 614454
rect 541222 614218 541404 614454
rect 540804 614134 541404 614218
rect 540804 613898 540986 614134
rect 541222 613898 541404 614134
rect 540804 578454 541404 613898
rect 540804 578218 540986 578454
rect 541222 578218 541404 578454
rect 540804 578134 541404 578218
rect 540804 577898 540986 578134
rect 541222 577898 541404 578134
rect 540804 542454 541404 577898
rect 540804 542218 540986 542454
rect 541222 542218 541404 542454
rect 540804 542134 541404 542218
rect 540804 541898 540986 542134
rect 541222 541898 541404 542134
rect 540804 506454 541404 541898
rect 540804 506218 540986 506454
rect 541222 506218 541404 506454
rect 540804 506134 541404 506218
rect 540804 505898 540986 506134
rect 541222 505898 541404 506134
rect 540804 470454 541404 505898
rect 540804 470218 540986 470454
rect 541222 470218 541404 470454
rect 540804 470134 541404 470218
rect 540804 469898 540986 470134
rect 541222 469898 541404 470134
rect 540804 434454 541404 469898
rect 540804 434218 540986 434454
rect 541222 434218 541404 434454
rect 540804 434134 541404 434218
rect 540804 433898 540986 434134
rect 541222 433898 541404 434134
rect 540804 398454 541404 433898
rect 540804 398218 540986 398454
rect 541222 398218 541404 398454
rect 540804 398134 541404 398218
rect 540804 397898 540986 398134
rect 541222 397898 541404 398134
rect 540804 362454 541404 397898
rect 540804 362218 540986 362454
rect 541222 362218 541404 362454
rect 540804 362134 541404 362218
rect 540804 361898 540986 362134
rect 541222 361898 541404 362134
rect 540804 326454 541404 361898
rect 540804 326218 540986 326454
rect 541222 326218 541404 326454
rect 540804 326134 541404 326218
rect 540804 325898 540986 326134
rect 541222 325898 541404 326134
rect 540804 290454 541404 325898
rect 540804 290218 540986 290454
rect 541222 290218 541404 290454
rect 540804 290134 541404 290218
rect 540804 289898 540986 290134
rect 541222 289898 541404 290134
rect 540804 254454 541404 289898
rect 540804 254218 540986 254454
rect 541222 254218 541404 254454
rect 540804 254134 541404 254218
rect 540804 253898 540986 254134
rect 541222 253898 541404 254134
rect 540804 218454 541404 253898
rect 540804 218218 540986 218454
rect 541222 218218 541404 218454
rect 540804 218134 541404 218218
rect 540804 217898 540986 218134
rect 541222 217898 541404 218134
rect 540804 182454 541404 217898
rect 540804 182218 540986 182454
rect 541222 182218 541404 182454
rect 540804 182134 541404 182218
rect 540804 181898 540986 182134
rect 541222 181898 541404 182134
rect 540804 146454 541404 181898
rect 540804 146218 540986 146454
rect 541222 146218 541404 146454
rect 540804 146134 541404 146218
rect 540804 145898 540986 146134
rect 541222 145898 541404 146134
rect 540804 110454 541404 145898
rect 540804 110218 540986 110454
rect 541222 110218 541404 110454
rect 540804 110134 541404 110218
rect 540804 109898 540986 110134
rect 541222 109898 541404 110134
rect 540804 74454 541404 109898
rect 540804 74218 540986 74454
rect 541222 74218 541404 74454
rect 540804 74134 541404 74218
rect 540804 73898 540986 74134
rect 541222 73898 541404 74134
rect 540804 38454 541404 73898
rect 540804 38218 540986 38454
rect 541222 38218 541404 38454
rect 540804 38134 541404 38218
rect 540804 37898 540986 38134
rect 541222 37898 541404 38134
rect 540804 2454 541404 37898
rect 540804 2218 540986 2454
rect 541222 2218 541404 2454
rect 540804 2134 541404 2218
rect 540804 1898 540986 2134
rect 541222 1898 541404 2134
rect 540804 -346 541404 1898
rect 540804 -582 540986 -346
rect 541222 -582 541404 -346
rect 540804 -666 541404 -582
rect 540804 -902 540986 -666
rect 541222 -902 541404 -666
rect 540804 -1864 541404 -902
rect 544404 690054 545004 706162
rect 544404 689818 544586 690054
rect 544822 689818 545004 690054
rect 544404 689734 545004 689818
rect 544404 689498 544586 689734
rect 544822 689498 545004 689734
rect 544404 654054 545004 689498
rect 544404 653818 544586 654054
rect 544822 653818 545004 654054
rect 544404 653734 545004 653818
rect 544404 653498 544586 653734
rect 544822 653498 545004 653734
rect 544404 618054 545004 653498
rect 544404 617818 544586 618054
rect 544822 617818 545004 618054
rect 544404 617734 545004 617818
rect 544404 617498 544586 617734
rect 544822 617498 545004 617734
rect 544404 582054 545004 617498
rect 544404 581818 544586 582054
rect 544822 581818 545004 582054
rect 544404 581734 545004 581818
rect 544404 581498 544586 581734
rect 544822 581498 545004 581734
rect 544404 546054 545004 581498
rect 544404 545818 544586 546054
rect 544822 545818 545004 546054
rect 544404 545734 545004 545818
rect 544404 545498 544586 545734
rect 544822 545498 545004 545734
rect 544404 510054 545004 545498
rect 544404 509818 544586 510054
rect 544822 509818 545004 510054
rect 544404 509734 545004 509818
rect 544404 509498 544586 509734
rect 544822 509498 545004 509734
rect 544404 474054 545004 509498
rect 544404 473818 544586 474054
rect 544822 473818 545004 474054
rect 544404 473734 545004 473818
rect 544404 473498 544586 473734
rect 544822 473498 545004 473734
rect 544404 438054 545004 473498
rect 544404 437818 544586 438054
rect 544822 437818 545004 438054
rect 544404 437734 545004 437818
rect 544404 437498 544586 437734
rect 544822 437498 545004 437734
rect 544404 402054 545004 437498
rect 544404 401818 544586 402054
rect 544822 401818 545004 402054
rect 544404 401734 545004 401818
rect 544404 401498 544586 401734
rect 544822 401498 545004 401734
rect 544404 366054 545004 401498
rect 544404 365818 544586 366054
rect 544822 365818 545004 366054
rect 544404 365734 545004 365818
rect 544404 365498 544586 365734
rect 544822 365498 545004 365734
rect 544404 330054 545004 365498
rect 544404 329818 544586 330054
rect 544822 329818 545004 330054
rect 544404 329734 545004 329818
rect 544404 329498 544586 329734
rect 544822 329498 545004 329734
rect 544404 294054 545004 329498
rect 544404 293818 544586 294054
rect 544822 293818 545004 294054
rect 544404 293734 545004 293818
rect 544404 293498 544586 293734
rect 544822 293498 545004 293734
rect 544404 258054 545004 293498
rect 544404 257818 544586 258054
rect 544822 257818 545004 258054
rect 544404 257734 545004 257818
rect 544404 257498 544586 257734
rect 544822 257498 545004 257734
rect 544404 222054 545004 257498
rect 544404 221818 544586 222054
rect 544822 221818 545004 222054
rect 544404 221734 545004 221818
rect 544404 221498 544586 221734
rect 544822 221498 545004 221734
rect 544404 186054 545004 221498
rect 544404 185818 544586 186054
rect 544822 185818 545004 186054
rect 544404 185734 545004 185818
rect 544404 185498 544586 185734
rect 544822 185498 545004 185734
rect 544404 150054 545004 185498
rect 544404 149818 544586 150054
rect 544822 149818 545004 150054
rect 544404 149734 545004 149818
rect 544404 149498 544586 149734
rect 544822 149498 545004 149734
rect 544404 114054 545004 149498
rect 544404 113818 544586 114054
rect 544822 113818 545004 114054
rect 544404 113734 545004 113818
rect 544404 113498 544586 113734
rect 544822 113498 545004 113734
rect 544404 78054 545004 113498
rect 544404 77818 544586 78054
rect 544822 77818 545004 78054
rect 544404 77734 545004 77818
rect 544404 77498 544586 77734
rect 544822 77498 545004 77734
rect 544404 42054 545004 77498
rect 544404 41818 544586 42054
rect 544822 41818 545004 42054
rect 544404 41734 545004 41818
rect 544404 41498 544586 41734
rect 544822 41498 545004 41734
rect 544404 6054 545004 41498
rect 544404 5818 544586 6054
rect 544822 5818 545004 6054
rect 544404 5734 545004 5818
rect 544404 5498 544586 5734
rect 544822 5498 545004 5734
rect 544404 -2226 545004 5498
rect 544404 -2462 544586 -2226
rect 544822 -2462 545004 -2226
rect 544404 -2546 545004 -2462
rect 544404 -2782 544586 -2546
rect 544822 -2782 545004 -2546
rect 544404 -3744 545004 -2782
rect 548004 693654 548604 708042
rect 548004 693418 548186 693654
rect 548422 693418 548604 693654
rect 548004 693334 548604 693418
rect 548004 693098 548186 693334
rect 548422 693098 548604 693334
rect 548004 657654 548604 693098
rect 548004 657418 548186 657654
rect 548422 657418 548604 657654
rect 548004 657334 548604 657418
rect 548004 657098 548186 657334
rect 548422 657098 548604 657334
rect 548004 621654 548604 657098
rect 548004 621418 548186 621654
rect 548422 621418 548604 621654
rect 548004 621334 548604 621418
rect 548004 621098 548186 621334
rect 548422 621098 548604 621334
rect 548004 585654 548604 621098
rect 548004 585418 548186 585654
rect 548422 585418 548604 585654
rect 548004 585334 548604 585418
rect 548004 585098 548186 585334
rect 548422 585098 548604 585334
rect 548004 549654 548604 585098
rect 548004 549418 548186 549654
rect 548422 549418 548604 549654
rect 548004 549334 548604 549418
rect 548004 549098 548186 549334
rect 548422 549098 548604 549334
rect 548004 513654 548604 549098
rect 548004 513418 548186 513654
rect 548422 513418 548604 513654
rect 548004 513334 548604 513418
rect 548004 513098 548186 513334
rect 548422 513098 548604 513334
rect 548004 477654 548604 513098
rect 548004 477418 548186 477654
rect 548422 477418 548604 477654
rect 548004 477334 548604 477418
rect 548004 477098 548186 477334
rect 548422 477098 548604 477334
rect 548004 441654 548604 477098
rect 548004 441418 548186 441654
rect 548422 441418 548604 441654
rect 548004 441334 548604 441418
rect 548004 441098 548186 441334
rect 548422 441098 548604 441334
rect 548004 405654 548604 441098
rect 548004 405418 548186 405654
rect 548422 405418 548604 405654
rect 548004 405334 548604 405418
rect 548004 405098 548186 405334
rect 548422 405098 548604 405334
rect 548004 369654 548604 405098
rect 548004 369418 548186 369654
rect 548422 369418 548604 369654
rect 548004 369334 548604 369418
rect 548004 369098 548186 369334
rect 548422 369098 548604 369334
rect 548004 333654 548604 369098
rect 548004 333418 548186 333654
rect 548422 333418 548604 333654
rect 548004 333334 548604 333418
rect 548004 333098 548186 333334
rect 548422 333098 548604 333334
rect 548004 297654 548604 333098
rect 548004 297418 548186 297654
rect 548422 297418 548604 297654
rect 548004 297334 548604 297418
rect 548004 297098 548186 297334
rect 548422 297098 548604 297334
rect 548004 261654 548604 297098
rect 548004 261418 548186 261654
rect 548422 261418 548604 261654
rect 548004 261334 548604 261418
rect 548004 261098 548186 261334
rect 548422 261098 548604 261334
rect 548004 225654 548604 261098
rect 548004 225418 548186 225654
rect 548422 225418 548604 225654
rect 548004 225334 548604 225418
rect 548004 225098 548186 225334
rect 548422 225098 548604 225334
rect 548004 189654 548604 225098
rect 548004 189418 548186 189654
rect 548422 189418 548604 189654
rect 548004 189334 548604 189418
rect 548004 189098 548186 189334
rect 548422 189098 548604 189334
rect 548004 153654 548604 189098
rect 548004 153418 548186 153654
rect 548422 153418 548604 153654
rect 548004 153334 548604 153418
rect 548004 153098 548186 153334
rect 548422 153098 548604 153334
rect 548004 117654 548604 153098
rect 548004 117418 548186 117654
rect 548422 117418 548604 117654
rect 548004 117334 548604 117418
rect 548004 117098 548186 117334
rect 548422 117098 548604 117334
rect 548004 81654 548604 117098
rect 548004 81418 548186 81654
rect 548422 81418 548604 81654
rect 548004 81334 548604 81418
rect 548004 81098 548186 81334
rect 548422 81098 548604 81334
rect 548004 45654 548604 81098
rect 548004 45418 548186 45654
rect 548422 45418 548604 45654
rect 548004 45334 548604 45418
rect 548004 45098 548186 45334
rect 548422 45098 548604 45334
rect 548004 9654 548604 45098
rect 548004 9418 548186 9654
rect 548422 9418 548604 9654
rect 548004 9334 548604 9418
rect 548004 9098 548186 9334
rect 548422 9098 548604 9334
rect 548004 -4106 548604 9098
rect 548004 -4342 548186 -4106
rect 548422 -4342 548604 -4106
rect 548004 -4426 548604 -4342
rect 548004 -4662 548186 -4426
rect 548422 -4662 548604 -4426
rect 548004 -5624 548604 -4662
rect 551604 697254 552204 709922
rect 569604 711418 570204 711440
rect 569604 711182 569786 711418
rect 570022 711182 570204 711418
rect 569604 711098 570204 711182
rect 569604 710862 569786 711098
rect 570022 710862 570204 711098
rect 566004 709538 566604 709560
rect 566004 709302 566186 709538
rect 566422 709302 566604 709538
rect 566004 709218 566604 709302
rect 566004 708982 566186 709218
rect 566422 708982 566604 709218
rect 562404 707658 563004 707680
rect 562404 707422 562586 707658
rect 562822 707422 563004 707658
rect 562404 707338 563004 707422
rect 562404 707102 562586 707338
rect 562822 707102 563004 707338
rect 551604 697018 551786 697254
rect 552022 697018 552204 697254
rect 551604 696934 552204 697018
rect 551604 696698 551786 696934
rect 552022 696698 552204 696934
rect 551604 661254 552204 696698
rect 551604 661018 551786 661254
rect 552022 661018 552204 661254
rect 551604 660934 552204 661018
rect 551604 660698 551786 660934
rect 552022 660698 552204 660934
rect 551604 625254 552204 660698
rect 551604 625018 551786 625254
rect 552022 625018 552204 625254
rect 551604 624934 552204 625018
rect 551604 624698 551786 624934
rect 552022 624698 552204 624934
rect 551604 589254 552204 624698
rect 551604 589018 551786 589254
rect 552022 589018 552204 589254
rect 551604 588934 552204 589018
rect 551604 588698 551786 588934
rect 552022 588698 552204 588934
rect 551604 553254 552204 588698
rect 551604 553018 551786 553254
rect 552022 553018 552204 553254
rect 551604 552934 552204 553018
rect 551604 552698 551786 552934
rect 552022 552698 552204 552934
rect 551604 517254 552204 552698
rect 551604 517018 551786 517254
rect 552022 517018 552204 517254
rect 551604 516934 552204 517018
rect 551604 516698 551786 516934
rect 552022 516698 552204 516934
rect 551604 481254 552204 516698
rect 551604 481018 551786 481254
rect 552022 481018 552204 481254
rect 551604 480934 552204 481018
rect 551604 480698 551786 480934
rect 552022 480698 552204 480934
rect 551604 445254 552204 480698
rect 551604 445018 551786 445254
rect 552022 445018 552204 445254
rect 551604 444934 552204 445018
rect 551604 444698 551786 444934
rect 552022 444698 552204 444934
rect 551604 409254 552204 444698
rect 551604 409018 551786 409254
rect 552022 409018 552204 409254
rect 551604 408934 552204 409018
rect 551604 408698 551786 408934
rect 552022 408698 552204 408934
rect 551604 373254 552204 408698
rect 551604 373018 551786 373254
rect 552022 373018 552204 373254
rect 551604 372934 552204 373018
rect 551604 372698 551786 372934
rect 552022 372698 552204 372934
rect 551604 337254 552204 372698
rect 551604 337018 551786 337254
rect 552022 337018 552204 337254
rect 551604 336934 552204 337018
rect 551604 336698 551786 336934
rect 552022 336698 552204 336934
rect 551604 301254 552204 336698
rect 551604 301018 551786 301254
rect 552022 301018 552204 301254
rect 551604 300934 552204 301018
rect 551604 300698 551786 300934
rect 552022 300698 552204 300934
rect 551604 265254 552204 300698
rect 551604 265018 551786 265254
rect 552022 265018 552204 265254
rect 551604 264934 552204 265018
rect 551604 264698 551786 264934
rect 552022 264698 552204 264934
rect 551604 229254 552204 264698
rect 551604 229018 551786 229254
rect 552022 229018 552204 229254
rect 551604 228934 552204 229018
rect 551604 228698 551786 228934
rect 552022 228698 552204 228934
rect 551604 193254 552204 228698
rect 551604 193018 551786 193254
rect 552022 193018 552204 193254
rect 551604 192934 552204 193018
rect 551604 192698 551786 192934
rect 552022 192698 552204 192934
rect 551604 157254 552204 192698
rect 551604 157018 551786 157254
rect 552022 157018 552204 157254
rect 551604 156934 552204 157018
rect 551604 156698 551786 156934
rect 552022 156698 552204 156934
rect 551604 121254 552204 156698
rect 551604 121018 551786 121254
rect 552022 121018 552204 121254
rect 551604 120934 552204 121018
rect 551604 120698 551786 120934
rect 552022 120698 552204 120934
rect 551604 85254 552204 120698
rect 551604 85018 551786 85254
rect 552022 85018 552204 85254
rect 551604 84934 552204 85018
rect 551604 84698 551786 84934
rect 552022 84698 552204 84934
rect 551604 49254 552204 84698
rect 551604 49018 551786 49254
rect 552022 49018 552204 49254
rect 551604 48934 552204 49018
rect 551604 48698 551786 48934
rect 552022 48698 552204 48934
rect 551604 13254 552204 48698
rect 551604 13018 551786 13254
rect 552022 13018 552204 13254
rect 551604 12934 552204 13018
rect 551604 12698 551786 12934
rect 552022 12698 552204 12934
rect 533604 -7162 533786 -6926
rect 534022 -7162 534204 -6926
rect 533604 -7246 534204 -7162
rect 533604 -7482 533786 -7246
rect 534022 -7482 534204 -7246
rect 533604 -7504 534204 -7482
rect 551604 -5986 552204 12698
rect 558804 705778 559404 705800
rect 558804 705542 558986 705778
rect 559222 705542 559404 705778
rect 558804 705458 559404 705542
rect 558804 705222 558986 705458
rect 559222 705222 559404 705458
rect 558804 668454 559404 705222
rect 558804 668218 558986 668454
rect 559222 668218 559404 668454
rect 558804 668134 559404 668218
rect 558804 667898 558986 668134
rect 559222 667898 559404 668134
rect 558804 632454 559404 667898
rect 558804 632218 558986 632454
rect 559222 632218 559404 632454
rect 558804 632134 559404 632218
rect 558804 631898 558986 632134
rect 559222 631898 559404 632134
rect 558804 596454 559404 631898
rect 558804 596218 558986 596454
rect 559222 596218 559404 596454
rect 558804 596134 559404 596218
rect 558804 595898 558986 596134
rect 559222 595898 559404 596134
rect 558804 560454 559404 595898
rect 558804 560218 558986 560454
rect 559222 560218 559404 560454
rect 558804 560134 559404 560218
rect 558804 559898 558986 560134
rect 559222 559898 559404 560134
rect 558804 524454 559404 559898
rect 558804 524218 558986 524454
rect 559222 524218 559404 524454
rect 558804 524134 559404 524218
rect 558804 523898 558986 524134
rect 559222 523898 559404 524134
rect 558804 488454 559404 523898
rect 558804 488218 558986 488454
rect 559222 488218 559404 488454
rect 558804 488134 559404 488218
rect 558804 487898 558986 488134
rect 559222 487898 559404 488134
rect 558804 452454 559404 487898
rect 558804 452218 558986 452454
rect 559222 452218 559404 452454
rect 558804 452134 559404 452218
rect 558804 451898 558986 452134
rect 559222 451898 559404 452134
rect 558804 416454 559404 451898
rect 558804 416218 558986 416454
rect 559222 416218 559404 416454
rect 558804 416134 559404 416218
rect 558804 415898 558986 416134
rect 559222 415898 559404 416134
rect 558804 380454 559404 415898
rect 558804 380218 558986 380454
rect 559222 380218 559404 380454
rect 558804 380134 559404 380218
rect 558804 379898 558986 380134
rect 559222 379898 559404 380134
rect 558804 344454 559404 379898
rect 558804 344218 558986 344454
rect 559222 344218 559404 344454
rect 558804 344134 559404 344218
rect 558804 343898 558986 344134
rect 559222 343898 559404 344134
rect 558804 308454 559404 343898
rect 558804 308218 558986 308454
rect 559222 308218 559404 308454
rect 558804 308134 559404 308218
rect 558804 307898 558986 308134
rect 559222 307898 559404 308134
rect 558804 272454 559404 307898
rect 558804 272218 558986 272454
rect 559222 272218 559404 272454
rect 558804 272134 559404 272218
rect 558804 271898 558986 272134
rect 559222 271898 559404 272134
rect 558804 236454 559404 271898
rect 558804 236218 558986 236454
rect 559222 236218 559404 236454
rect 558804 236134 559404 236218
rect 558804 235898 558986 236134
rect 559222 235898 559404 236134
rect 558804 200454 559404 235898
rect 558804 200218 558986 200454
rect 559222 200218 559404 200454
rect 558804 200134 559404 200218
rect 558804 199898 558986 200134
rect 559222 199898 559404 200134
rect 558804 164454 559404 199898
rect 558804 164218 558986 164454
rect 559222 164218 559404 164454
rect 558804 164134 559404 164218
rect 558804 163898 558986 164134
rect 559222 163898 559404 164134
rect 558804 128454 559404 163898
rect 558804 128218 558986 128454
rect 559222 128218 559404 128454
rect 558804 128134 559404 128218
rect 558804 127898 558986 128134
rect 559222 127898 559404 128134
rect 558804 92454 559404 127898
rect 558804 92218 558986 92454
rect 559222 92218 559404 92454
rect 558804 92134 559404 92218
rect 558804 91898 558986 92134
rect 559222 91898 559404 92134
rect 558804 56454 559404 91898
rect 558804 56218 558986 56454
rect 559222 56218 559404 56454
rect 558804 56134 559404 56218
rect 558804 55898 558986 56134
rect 559222 55898 559404 56134
rect 558804 20454 559404 55898
rect 558804 20218 558986 20454
rect 559222 20218 559404 20454
rect 558804 20134 559404 20218
rect 558804 19898 558986 20134
rect 559222 19898 559404 20134
rect 558804 -1286 559404 19898
rect 558804 -1522 558986 -1286
rect 559222 -1522 559404 -1286
rect 558804 -1606 559404 -1522
rect 558804 -1842 558986 -1606
rect 559222 -1842 559404 -1606
rect 558804 -1864 559404 -1842
rect 562404 672054 563004 707102
rect 562404 671818 562586 672054
rect 562822 671818 563004 672054
rect 562404 671734 563004 671818
rect 562404 671498 562586 671734
rect 562822 671498 563004 671734
rect 562404 636054 563004 671498
rect 562404 635818 562586 636054
rect 562822 635818 563004 636054
rect 562404 635734 563004 635818
rect 562404 635498 562586 635734
rect 562822 635498 563004 635734
rect 562404 600054 563004 635498
rect 562404 599818 562586 600054
rect 562822 599818 563004 600054
rect 562404 599734 563004 599818
rect 562404 599498 562586 599734
rect 562822 599498 563004 599734
rect 562404 564054 563004 599498
rect 562404 563818 562586 564054
rect 562822 563818 563004 564054
rect 562404 563734 563004 563818
rect 562404 563498 562586 563734
rect 562822 563498 563004 563734
rect 562404 528054 563004 563498
rect 562404 527818 562586 528054
rect 562822 527818 563004 528054
rect 562404 527734 563004 527818
rect 562404 527498 562586 527734
rect 562822 527498 563004 527734
rect 562404 492054 563004 527498
rect 562404 491818 562586 492054
rect 562822 491818 563004 492054
rect 562404 491734 563004 491818
rect 562404 491498 562586 491734
rect 562822 491498 563004 491734
rect 562404 456054 563004 491498
rect 562404 455818 562586 456054
rect 562822 455818 563004 456054
rect 562404 455734 563004 455818
rect 562404 455498 562586 455734
rect 562822 455498 563004 455734
rect 562404 420054 563004 455498
rect 562404 419818 562586 420054
rect 562822 419818 563004 420054
rect 562404 419734 563004 419818
rect 562404 419498 562586 419734
rect 562822 419498 563004 419734
rect 562404 384054 563004 419498
rect 562404 383818 562586 384054
rect 562822 383818 563004 384054
rect 562404 383734 563004 383818
rect 562404 383498 562586 383734
rect 562822 383498 563004 383734
rect 562404 348054 563004 383498
rect 562404 347818 562586 348054
rect 562822 347818 563004 348054
rect 562404 347734 563004 347818
rect 562404 347498 562586 347734
rect 562822 347498 563004 347734
rect 562404 312054 563004 347498
rect 562404 311818 562586 312054
rect 562822 311818 563004 312054
rect 562404 311734 563004 311818
rect 562404 311498 562586 311734
rect 562822 311498 563004 311734
rect 562404 276054 563004 311498
rect 562404 275818 562586 276054
rect 562822 275818 563004 276054
rect 562404 275734 563004 275818
rect 562404 275498 562586 275734
rect 562822 275498 563004 275734
rect 562404 240054 563004 275498
rect 562404 239818 562586 240054
rect 562822 239818 563004 240054
rect 562404 239734 563004 239818
rect 562404 239498 562586 239734
rect 562822 239498 563004 239734
rect 562404 204054 563004 239498
rect 562404 203818 562586 204054
rect 562822 203818 563004 204054
rect 562404 203734 563004 203818
rect 562404 203498 562586 203734
rect 562822 203498 563004 203734
rect 562404 168054 563004 203498
rect 562404 167818 562586 168054
rect 562822 167818 563004 168054
rect 562404 167734 563004 167818
rect 562404 167498 562586 167734
rect 562822 167498 563004 167734
rect 562404 132054 563004 167498
rect 562404 131818 562586 132054
rect 562822 131818 563004 132054
rect 562404 131734 563004 131818
rect 562404 131498 562586 131734
rect 562822 131498 563004 131734
rect 562404 96054 563004 131498
rect 562404 95818 562586 96054
rect 562822 95818 563004 96054
rect 562404 95734 563004 95818
rect 562404 95498 562586 95734
rect 562822 95498 563004 95734
rect 562404 60054 563004 95498
rect 562404 59818 562586 60054
rect 562822 59818 563004 60054
rect 562404 59734 563004 59818
rect 562404 59498 562586 59734
rect 562822 59498 563004 59734
rect 562404 24054 563004 59498
rect 562404 23818 562586 24054
rect 562822 23818 563004 24054
rect 562404 23734 563004 23818
rect 562404 23498 562586 23734
rect 562822 23498 563004 23734
rect 562404 -3166 563004 23498
rect 562404 -3402 562586 -3166
rect 562822 -3402 563004 -3166
rect 562404 -3486 563004 -3402
rect 562404 -3722 562586 -3486
rect 562822 -3722 563004 -3486
rect 562404 -3744 563004 -3722
rect 566004 675654 566604 708982
rect 566004 675418 566186 675654
rect 566422 675418 566604 675654
rect 566004 675334 566604 675418
rect 566004 675098 566186 675334
rect 566422 675098 566604 675334
rect 566004 639654 566604 675098
rect 566004 639418 566186 639654
rect 566422 639418 566604 639654
rect 566004 639334 566604 639418
rect 566004 639098 566186 639334
rect 566422 639098 566604 639334
rect 566004 603654 566604 639098
rect 566004 603418 566186 603654
rect 566422 603418 566604 603654
rect 566004 603334 566604 603418
rect 566004 603098 566186 603334
rect 566422 603098 566604 603334
rect 566004 567654 566604 603098
rect 566004 567418 566186 567654
rect 566422 567418 566604 567654
rect 566004 567334 566604 567418
rect 566004 567098 566186 567334
rect 566422 567098 566604 567334
rect 566004 531654 566604 567098
rect 566004 531418 566186 531654
rect 566422 531418 566604 531654
rect 566004 531334 566604 531418
rect 566004 531098 566186 531334
rect 566422 531098 566604 531334
rect 566004 495654 566604 531098
rect 566004 495418 566186 495654
rect 566422 495418 566604 495654
rect 566004 495334 566604 495418
rect 566004 495098 566186 495334
rect 566422 495098 566604 495334
rect 566004 459654 566604 495098
rect 566004 459418 566186 459654
rect 566422 459418 566604 459654
rect 566004 459334 566604 459418
rect 566004 459098 566186 459334
rect 566422 459098 566604 459334
rect 566004 423654 566604 459098
rect 566004 423418 566186 423654
rect 566422 423418 566604 423654
rect 566004 423334 566604 423418
rect 566004 423098 566186 423334
rect 566422 423098 566604 423334
rect 566004 387654 566604 423098
rect 566004 387418 566186 387654
rect 566422 387418 566604 387654
rect 566004 387334 566604 387418
rect 566004 387098 566186 387334
rect 566422 387098 566604 387334
rect 566004 351654 566604 387098
rect 566004 351418 566186 351654
rect 566422 351418 566604 351654
rect 566004 351334 566604 351418
rect 566004 351098 566186 351334
rect 566422 351098 566604 351334
rect 566004 315654 566604 351098
rect 566004 315418 566186 315654
rect 566422 315418 566604 315654
rect 566004 315334 566604 315418
rect 566004 315098 566186 315334
rect 566422 315098 566604 315334
rect 566004 279654 566604 315098
rect 566004 279418 566186 279654
rect 566422 279418 566604 279654
rect 566004 279334 566604 279418
rect 566004 279098 566186 279334
rect 566422 279098 566604 279334
rect 566004 243654 566604 279098
rect 566004 243418 566186 243654
rect 566422 243418 566604 243654
rect 566004 243334 566604 243418
rect 566004 243098 566186 243334
rect 566422 243098 566604 243334
rect 566004 207654 566604 243098
rect 566004 207418 566186 207654
rect 566422 207418 566604 207654
rect 566004 207334 566604 207418
rect 566004 207098 566186 207334
rect 566422 207098 566604 207334
rect 566004 171654 566604 207098
rect 566004 171418 566186 171654
rect 566422 171418 566604 171654
rect 566004 171334 566604 171418
rect 566004 171098 566186 171334
rect 566422 171098 566604 171334
rect 566004 135654 566604 171098
rect 566004 135418 566186 135654
rect 566422 135418 566604 135654
rect 566004 135334 566604 135418
rect 566004 135098 566186 135334
rect 566422 135098 566604 135334
rect 566004 99654 566604 135098
rect 566004 99418 566186 99654
rect 566422 99418 566604 99654
rect 566004 99334 566604 99418
rect 566004 99098 566186 99334
rect 566422 99098 566604 99334
rect 566004 63654 566604 99098
rect 566004 63418 566186 63654
rect 566422 63418 566604 63654
rect 566004 63334 566604 63418
rect 566004 63098 566186 63334
rect 566422 63098 566604 63334
rect 566004 27654 566604 63098
rect 566004 27418 566186 27654
rect 566422 27418 566604 27654
rect 566004 27334 566604 27418
rect 566004 27098 566186 27334
rect 566422 27098 566604 27334
rect 566004 -5046 566604 27098
rect 566004 -5282 566186 -5046
rect 566422 -5282 566604 -5046
rect 566004 -5366 566604 -5282
rect 566004 -5602 566186 -5366
rect 566422 -5602 566604 -5366
rect 566004 -5624 566604 -5602
rect 569604 679254 570204 710862
rect 591900 711418 592500 711440
rect 591900 711182 592082 711418
rect 592318 711182 592500 711418
rect 591900 711098 592500 711182
rect 591900 710862 592082 711098
rect 592318 710862 592500 711098
rect 590960 710478 591560 710500
rect 590960 710242 591142 710478
rect 591378 710242 591560 710478
rect 590960 710158 591560 710242
rect 590960 709922 591142 710158
rect 591378 709922 591560 710158
rect 590020 709538 590620 709560
rect 590020 709302 590202 709538
rect 590438 709302 590620 709538
rect 590020 709218 590620 709302
rect 590020 708982 590202 709218
rect 590438 708982 590620 709218
rect 589080 708598 589680 708620
rect 589080 708362 589262 708598
rect 589498 708362 589680 708598
rect 589080 708278 589680 708362
rect 589080 708042 589262 708278
rect 589498 708042 589680 708278
rect 580404 706718 581004 707680
rect 588140 707658 588740 707680
rect 588140 707422 588322 707658
rect 588558 707422 588740 707658
rect 588140 707338 588740 707422
rect 588140 707102 588322 707338
rect 588558 707102 588740 707338
rect 580404 706482 580586 706718
rect 580822 706482 581004 706718
rect 580404 706398 581004 706482
rect 580404 706162 580586 706398
rect 580822 706162 581004 706398
rect 569604 679018 569786 679254
rect 570022 679018 570204 679254
rect 569604 678934 570204 679018
rect 569604 678698 569786 678934
rect 570022 678698 570204 678934
rect 569604 643254 570204 678698
rect 569604 643018 569786 643254
rect 570022 643018 570204 643254
rect 569604 642934 570204 643018
rect 569604 642698 569786 642934
rect 570022 642698 570204 642934
rect 569604 607254 570204 642698
rect 569604 607018 569786 607254
rect 570022 607018 570204 607254
rect 569604 606934 570204 607018
rect 569604 606698 569786 606934
rect 570022 606698 570204 606934
rect 569604 571254 570204 606698
rect 569604 571018 569786 571254
rect 570022 571018 570204 571254
rect 569604 570934 570204 571018
rect 569604 570698 569786 570934
rect 570022 570698 570204 570934
rect 569604 535254 570204 570698
rect 569604 535018 569786 535254
rect 570022 535018 570204 535254
rect 569604 534934 570204 535018
rect 569604 534698 569786 534934
rect 570022 534698 570204 534934
rect 569604 499254 570204 534698
rect 569604 499018 569786 499254
rect 570022 499018 570204 499254
rect 569604 498934 570204 499018
rect 569604 498698 569786 498934
rect 570022 498698 570204 498934
rect 569604 463254 570204 498698
rect 569604 463018 569786 463254
rect 570022 463018 570204 463254
rect 569604 462934 570204 463018
rect 569604 462698 569786 462934
rect 570022 462698 570204 462934
rect 569604 427254 570204 462698
rect 569604 427018 569786 427254
rect 570022 427018 570204 427254
rect 569604 426934 570204 427018
rect 569604 426698 569786 426934
rect 570022 426698 570204 426934
rect 569604 391254 570204 426698
rect 569604 391018 569786 391254
rect 570022 391018 570204 391254
rect 569604 390934 570204 391018
rect 569604 390698 569786 390934
rect 570022 390698 570204 390934
rect 569604 355254 570204 390698
rect 569604 355018 569786 355254
rect 570022 355018 570204 355254
rect 569604 354934 570204 355018
rect 569604 354698 569786 354934
rect 570022 354698 570204 354934
rect 569604 319254 570204 354698
rect 569604 319018 569786 319254
rect 570022 319018 570204 319254
rect 569604 318934 570204 319018
rect 569604 318698 569786 318934
rect 570022 318698 570204 318934
rect 569604 283254 570204 318698
rect 569604 283018 569786 283254
rect 570022 283018 570204 283254
rect 569604 282934 570204 283018
rect 569604 282698 569786 282934
rect 570022 282698 570204 282934
rect 569604 247254 570204 282698
rect 569604 247018 569786 247254
rect 570022 247018 570204 247254
rect 569604 246934 570204 247018
rect 569604 246698 569786 246934
rect 570022 246698 570204 246934
rect 569604 211254 570204 246698
rect 569604 211018 569786 211254
rect 570022 211018 570204 211254
rect 569604 210934 570204 211018
rect 569604 210698 569786 210934
rect 570022 210698 570204 210934
rect 569604 175254 570204 210698
rect 569604 175018 569786 175254
rect 570022 175018 570204 175254
rect 569604 174934 570204 175018
rect 569604 174698 569786 174934
rect 570022 174698 570204 174934
rect 569604 139254 570204 174698
rect 569604 139018 569786 139254
rect 570022 139018 570204 139254
rect 569604 138934 570204 139018
rect 569604 138698 569786 138934
rect 570022 138698 570204 138934
rect 569604 103254 570204 138698
rect 569604 103018 569786 103254
rect 570022 103018 570204 103254
rect 569604 102934 570204 103018
rect 569604 102698 569786 102934
rect 570022 102698 570204 102934
rect 569604 67254 570204 102698
rect 569604 67018 569786 67254
rect 570022 67018 570204 67254
rect 569604 66934 570204 67018
rect 569604 66698 569786 66934
rect 570022 66698 570204 66934
rect 569604 31254 570204 66698
rect 569604 31018 569786 31254
rect 570022 31018 570204 31254
rect 569604 30934 570204 31018
rect 569604 30698 569786 30934
rect 570022 30698 570204 30934
rect 551604 -6222 551786 -5986
rect 552022 -6222 552204 -5986
rect 551604 -6306 552204 -6222
rect 551604 -6542 551786 -6306
rect 552022 -6542 552204 -6306
rect 551604 -7504 552204 -6542
rect 569604 -6926 570204 30698
rect 576804 704838 577404 705800
rect 576804 704602 576986 704838
rect 577222 704602 577404 704838
rect 576804 704518 577404 704602
rect 576804 704282 576986 704518
rect 577222 704282 577404 704518
rect 576804 686454 577404 704282
rect 576804 686218 576986 686454
rect 577222 686218 577404 686454
rect 576804 686134 577404 686218
rect 576804 685898 576986 686134
rect 577222 685898 577404 686134
rect 576804 650454 577404 685898
rect 576804 650218 576986 650454
rect 577222 650218 577404 650454
rect 576804 650134 577404 650218
rect 576804 649898 576986 650134
rect 577222 649898 577404 650134
rect 576804 614454 577404 649898
rect 576804 614218 576986 614454
rect 577222 614218 577404 614454
rect 576804 614134 577404 614218
rect 576804 613898 576986 614134
rect 577222 613898 577404 614134
rect 576804 578454 577404 613898
rect 576804 578218 576986 578454
rect 577222 578218 577404 578454
rect 576804 578134 577404 578218
rect 576804 577898 576986 578134
rect 577222 577898 577404 578134
rect 576804 542454 577404 577898
rect 576804 542218 576986 542454
rect 577222 542218 577404 542454
rect 576804 542134 577404 542218
rect 576804 541898 576986 542134
rect 577222 541898 577404 542134
rect 576804 506454 577404 541898
rect 576804 506218 576986 506454
rect 577222 506218 577404 506454
rect 576804 506134 577404 506218
rect 576804 505898 576986 506134
rect 577222 505898 577404 506134
rect 576804 470454 577404 505898
rect 576804 470218 576986 470454
rect 577222 470218 577404 470454
rect 576804 470134 577404 470218
rect 576804 469898 576986 470134
rect 577222 469898 577404 470134
rect 576804 434454 577404 469898
rect 576804 434218 576986 434454
rect 577222 434218 577404 434454
rect 576804 434134 577404 434218
rect 576804 433898 576986 434134
rect 577222 433898 577404 434134
rect 576804 398454 577404 433898
rect 576804 398218 576986 398454
rect 577222 398218 577404 398454
rect 576804 398134 577404 398218
rect 576804 397898 576986 398134
rect 577222 397898 577404 398134
rect 576804 362454 577404 397898
rect 576804 362218 576986 362454
rect 577222 362218 577404 362454
rect 576804 362134 577404 362218
rect 576804 361898 576986 362134
rect 577222 361898 577404 362134
rect 576804 326454 577404 361898
rect 576804 326218 576986 326454
rect 577222 326218 577404 326454
rect 576804 326134 577404 326218
rect 576804 325898 576986 326134
rect 577222 325898 577404 326134
rect 576804 290454 577404 325898
rect 576804 290218 576986 290454
rect 577222 290218 577404 290454
rect 576804 290134 577404 290218
rect 576804 289898 576986 290134
rect 577222 289898 577404 290134
rect 576804 254454 577404 289898
rect 576804 254218 576986 254454
rect 577222 254218 577404 254454
rect 576804 254134 577404 254218
rect 576804 253898 576986 254134
rect 577222 253898 577404 254134
rect 576804 218454 577404 253898
rect 576804 218218 576986 218454
rect 577222 218218 577404 218454
rect 576804 218134 577404 218218
rect 576804 217898 576986 218134
rect 577222 217898 577404 218134
rect 576804 182454 577404 217898
rect 576804 182218 576986 182454
rect 577222 182218 577404 182454
rect 576804 182134 577404 182218
rect 576804 181898 576986 182134
rect 577222 181898 577404 182134
rect 576804 146454 577404 181898
rect 576804 146218 576986 146454
rect 577222 146218 577404 146454
rect 576804 146134 577404 146218
rect 576804 145898 576986 146134
rect 577222 145898 577404 146134
rect 576804 110454 577404 145898
rect 576804 110218 576986 110454
rect 577222 110218 577404 110454
rect 576804 110134 577404 110218
rect 576804 109898 576986 110134
rect 577222 109898 577404 110134
rect 576804 74454 577404 109898
rect 576804 74218 576986 74454
rect 577222 74218 577404 74454
rect 576804 74134 577404 74218
rect 576804 73898 576986 74134
rect 577222 73898 577404 74134
rect 576804 38454 577404 73898
rect 576804 38218 576986 38454
rect 577222 38218 577404 38454
rect 576804 38134 577404 38218
rect 576804 37898 576986 38134
rect 577222 37898 577404 38134
rect 576804 2454 577404 37898
rect 576804 2218 576986 2454
rect 577222 2218 577404 2454
rect 576804 2134 577404 2218
rect 576804 1898 576986 2134
rect 577222 1898 577404 2134
rect 576804 -346 577404 1898
rect 576804 -582 576986 -346
rect 577222 -582 577404 -346
rect 576804 -666 577404 -582
rect 576804 -902 576986 -666
rect 577222 -902 577404 -666
rect 576804 -1864 577404 -902
rect 580404 690054 581004 706162
rect 587200 706718 587800 706740
rect 587200 706482 587382 706718
rect 587618 706482 587800 706718
rect 587200 706398 587800 706482
rect 587200 706162 587382 706398
rect 587618 706162 587800 706398
rect 586260 705778 586860 705800
rect 586260 705542 586442 705778
rect 586678 705542 586860 705778
rect 586260 705458 586860 705542
rect 586260 705222 586442 705458
rect 586678 705222 586860 705458
rect 580404 689818 580586 690054
rect 580822 689818 581004 690054
rect 580404 689734 581004 689818
rect 580404 689498 580586 689734
rect 580822 689498 581004 689734
rect 580404 654054 581004 689498
rect 580404 653818 580586 654054
rect 580822 653818 581004 654054
rect 580404 653734 581004 653818
rect 580404 653498 580586 653734
rect 580822 653498 581004 653734
rect 580404 618054 581004 653498
rect 580404 617818 580586 618054
rect 580822 617818 581004 618054
rect 580404 617734 581004 617818
rect 580404 617498 580586 617734
rect 580822 617498 581004 617734
rect 580404 582054 581004 617498
rect 580404 581818 580586 582054
rect 580822 581818 581004 582054
rect 580404 581734 581004 581818
rect 580404 581498 580586 581734
rect 580822 581498 581004 581734
rect 580404 546054 581004 581498
rect 580404 545818 580586 546054
rect 580822 545818 581004 546054
rect 580404 545734 581004 545818
rect 580404 545498 580586 545734
rect 580822 545498 581004 545734
rect 580404 510054 581004 545498
rect 580404 509818 580586 510054
rect 580822 509818 581004 510054
rect 580404 509734 581004 509818
rect 580404 509498 580586 509734
rect 580822 509498 581004 509734
rect 580404 474054 581004 509498
rect 580404 473818 580586 474054
rect 580822 473818 581004 474054
rect 580404 473734 581004 473818
rect 580404 473498 580586 473734
rect 580822 473498 581004 473734
rect 580404 438054 581004 473498
rect 580404 437818 580586 438054
rect 580822 437818 581004 438054
rect 580404 437734 581004 437818
rect 580404 437498 580586 437734
rect 580822 437498 581004 437734
rect 580404 402054 581004 437498
rect 580404 401818 580586 402054
rect 580822 401818 581004 402054
rect 580404 401734 581004 401818
rect 580404 401498 580586 401734
rect 580822 401498 581004 401734
rect 580404 366054 581004 401498
rect 580404 365818 580586 366054
rect 580822 365818 581004 366054
rect 580404 365734 581004 365818
rect 580404 365498 580586 365734
rect 580822 365498 581004 365734
rect 580404 330054 581004 365498
rect 580404 329818 580586 330054
rect 580822 329818 581004 330054
rect 580404 329734 581004 329818
rect 580404 329498 580586 329734
rect 580822 329498 581004 329734
rect 580404 294054 581004 329498
rect 580404 293818 580586 294054
rect 580822 293818 581004 294054
rect 580404 293734 581004 293818
rect 580404 293498 580586 293734
rect 580822 293498 581004 293734
rect 580404 258054 581004 293498
rect 580404 257818 580586 258054
rect 580822 257818 581004 258054
rect 580404 257734 581004 257818
rect 580404 257498 580586 257734
rect 580822 257498 581004 257734
rect 580404 222054 581004 257498
rect 580404 221818 580586 222054
rect 580822 221818 581004 222054
rect 580404 221734 581004 221818
rect 580404 221498 580586 221734
rect 580822 221498 581004 221734
rect 580404 186054 581004 221498
rect 580404 185818 580586 186054
rect 580822 185818 581004 186054
rect 580404 185734 581004 185818
rect 580404 185498 580586 185734
rect 580822 185498 581004 185734
rect 580404 150054 581004 185498
rect 580404 149818 580586 150054
rect 580822 149818 581004 150054
rect 580404 149734 581004 149818
rect 580404 149498 580586 149734
rect 580822 149498 581004 149734
rect 580404 114054 581004 149498
rect 580404 113818 580586 114054
rect 580822 113818 581004 114054
rect 580404 113734 581004 113818
rect 580404 113498 580586 113734
rect 580822 113498 581004 113734
rect 580404 78054 581004 113498
rect 580404 77818 580586 78054
rect 580822 77818 581004 78054
rect 580404 77734 581004 77818
rect 580404 77498 580586 77734
rect 580822 77498 581004 77734
rect 580404 42054 581004 77498
rect 580404 41818 580586 42054
rect 580822 41818 581004 42054
rect 580404 41734 581004 41818
rect 580404 41498 580586 41734
rect 580822 41498 581004 41734
rect 580404 6054 581004 41498
rect 580404 5818 580586 6054
rect 580822 5818 581004 6054
rect 580404 5734 581004 5818
rect 580404 5498 580586 5734
rect 580822 5498 581004 5734
rect 580404 -2226 581004 5498
rect 585320 704838 585920 704860
rect 585320 704602 585502 704838
rect 585738 704602 585920 704838
rect 585320 704518 585920 704602
rect 585320 704282 585502 704518
rect 585738 704282 585920 704518
rect 585320 686454 585920 704282
rect 585320 686218 585502 686454
rect 585738 686218 585920 686454
rect 585320 686134 585920 686218
rect 585320 685898 585502 686134
rect 585738 685898 585920 686134
rect 585320 650454 585920 685898
rect 585320 650218 585502 650454
rect 585738 650218 585920 650454
rect 585320 650134 585920 650218
rect 585320 649898 585502 650134
rect 585738 649898 585920 650134
rect 585320 614454 585920 649898
rect 585320 614218 585502 614454
rect 585738 614218 585920 614454
rect 585320 614134 585920 614218
rect 585320 613898 585502 614134
rect 585738 613898 585920 614134
rect 585320 578454 585920 613898
rect 585320 578218 585502 578454
rect 585738 578218 585920 578454
rect 585320 578134 585920 578218
rect 585320 577898 585502 578134
rect 585738 577898 585920 578134
rect 585320 542454 585920 577898
rect 585320 542218 585502 542454
rect 585738 542218 585920 542454
rect 585320 542134 585920 542218
rect 585320 541898 585502 542134
rect 585738 541898 585920 542134
rect 585320 506454 585920 541898
rect 585320 506218 585502 506454
rect 585738 506218 585920 506454
rect 585320 506134 585920 506218
rect 585320 505898 585502 506134
rect 585738 505898 585920 506134
rect 585320 470454 585920 505898
rect 585320 470218 585502 470454
rect 585738 470218 585920 470454
rect 585320 470134 585920 470218
rect 585320 469898 585502 470134
rect 585738 469898 585920 470134
rect 585320 434454 585920 469898
rect 585320 434218 585502 434454
rect 585738 434218 585920 434454
rect 585320 434134 585920 434218
rect 585320 433898 585502 434134
rect 585738 433898 585920 434134
rect 585320 398454 585920 433898
rect 585320 398218 585502 398454
rect 585738 398218 585920 398454
rect 585320 398134 585920 398218
rect 585320 397898 585502 398134
rect 585738 397898 585920 398134
rect 585320 362454 585920 397898
rect 585320 362218 585502 362454
rect 585738 362218 585920 362454
rect 585320 362134 585920 362218
rect 585320 361898 585502 362134
rect 585738 361898 585920 362134
rect 585320 326454 585920 361898
rect 585320 326218 585502 326454
rect 585738 326218 585920 326454
rect 585320 326134 585920 326218
rect 585320 325898 585502 326134
rect 585738 325898 585920 326134
rect 585320 290454 585920 325898
rect 585320 290218 585502 290454
rect 585738 290218 585920 290454
rect 585320 290134 585920 290218
rect 585320 289898 585502 290134
rect 585738 289898 585920 290134
rect 585320 254454 585920 289898
rect 585320 254218 585502 254454
rect 585738 254218 585920 254454
rect 585320 254134 585920 254218
rect 585320 253898 585502 254134
rect 585738 253898 585920 254134
rect 585320 218454 585920 253898
rect 585320 218218 585502 218454
rect 585738 218218 585920 218454
rect 585320 218134 585920 218218
rect 585320 217898 585502 218134
rect 585738 217898 585920 218134
rect 585320 182454 585920 217898
rect 585320 182218 585502 182454
rect 585738 182218 585920 182454
rect 585320 182134 585920 182218
rect 585320 181898 585502 182134
rect 585738 181898 585920 182134
rect 585320 146454 585920 181898
rect 585320 146218 585502 146454
rect 585738 146218 585920 146454
rect 585320 146134 585920 146218
rect 585320 145898 585502 146134
rect 585738 145898 585920 146134
rect 585320 110454 585920 145898
rect 585320 110218 585502 110454
rect 585738 110218 585920 110454
rect 585320 110134 585920 110218
rect 585320 109898 585502 110134
rect 585738 109898 585920 110134
rect 585320 74454 585920 109898
rect 585320 74218 585502 74454
rect 585738 74218 585920 74454
rect 585320 74134 585920 74218
rect 585320 73898 585502 74134
rect 585738 73898 585920 74134
rect 585320 38454 585920 73898
rect 585320 38218 585502 38454
rect 585738 38218 585920 38454
rect 585320 38134 585920 38218
rect 585320 37898 585502 38134
rect 585738 37898 585920 38134
rect 585320 2454 585920 37898
rect 585320 2218 585502 2454
rect 585738 2218 585920 2454
rect 585320 2134 585920 2218
rect 585320 1898 585502 2134
rect 585738 1898 585920 2134
rect 585320 -346 585920 1898
rect 585320 -582 585502 -346
rect 585738 -582 585920 -346
rect 585320 -666 585920 -582
rect 585320 -902 585502 -666
rect 585738 -902 585920 -666
rect 585320 -924 585920 -902
rect 586260 668454 586860 705222
rect 586260 668218 586442 668454
rect 586678 668218 586860 668454
rect 586260 668134 586860 668218
rect 586260 667898 586442 668134
rect 586678 667898 586860 668134
rect 586260 632454 586860 667898
rect 586260 632218 586442 632454
rect 586678 632218 586860 632454
rect 586260 632134 586860 632218
rect 586260 631898 586442 632134
rect 586678 631898 586860 632134
rect 586260 596454 586860 631898
rect 586260 596218 586442 596454
rect 586678 596218 586860 596454
rect 586260 596134 586860 596218
rect 586260 595898 586442 596134
rect 586678 595898 586860 596134
rect 586260 560454 586860 595898
rect 586260 560218 586442 560454
rect 586678 560218 586860 560454
rect 586260 560134 586860 560218
rect 586260 559898 586442 560134
rect 586678 559898 586860 560134
rect 586260 524454 586860 559898
rect 586260 524218 586442 524454
rect 586678 524218 586860 524454
rect 586260 524134 586860 524218
rect 586260 523898 586442 524134
rect 586678 523898 586860 524134
rect 586260 488454 586860 523898
rect 586260 488218 586442 488454
rect 586678 488218 586860 488454
rect 586260 488134 586860 488218
rect 586260 487898 586442 488134
rect 586678 487898 586860 488134
rect 586260 452454 586860 487898
rect 586260 452218 586442 452454
rect 586678 452218 586860 452454
rect 586260 452134 586860 452218
rect 586260 451898 586442 452134
rect 586678 451898 586860 452134
rect 586260 416454 586860 451898
rect 586260 416218 586442 416454
rect 586678 416218 586860 416454
rect 586260 416134 586860 416218
rect 586260 415898 586442 416134
rect 586678 415898 586860 416134
rect 586260 380454 586860 415898
rect 586260 380218 586442 380454
rect 586678 380218 586860 380454
rect 586260 380134 586860 380218
rect 586260 379898 586442 380134
rect 586678 379898 586860 380134
rect 586260 344454 586860 379898
rect 586260 344218 586442 344454
rect 586678 344218 586860 344454
rect 586260 344134 586860 344218
rect 586260 343898 586442 344134
rect 586678 343898 586860 344134
rect 586260 308454 586860 343898
rect 586260 308218 586442 308454
rect 586678 308218 586860 308454
rect 586260 308134 586860 308218
rect 586260 307898 586442 308134
rect 586678 307898 586860 308134
rect 586260 272454 586860 307898
rect 586260 272218 586442 272454
rect 586678 272218 586860 272454
rect 586260 272134 586860 272218
rect 586260 271898 586442 272134
rect 586678 271898 586860 272134
rect 586260 236454 586860 271898
rect 586260 236218 586442 236454
rect 586678 236218 586860 236454
rect 586260 236134 586860 236218
rect 586260 235898 586442 236134
rect 586678 235898 586860 236134
rect 586260 200454 586860 235898
rect 586260 200218 586442 200454
rect 586678 200218 586860 200454
rect 586260 200134 586860 200218
rect 586260 199898 586442 200134
rect 586678 199898 586860 200134
rect 586260 164454 586860 199898
rect 586260 164218 586442 164454
rect 586678 164218 586860 164454
rect 586260 164134 586860 164218
rect 586260 163898 586442 164134
rect 586678 163898 586860 164134
rect 586260 128454 586860 163898
rect 586260 128218 586442 128454
rect 586678 128218 586860 128454
rect 586260 128134 586860 128218
rect 586260 127898 586442 128134
rect 586678 127898 586860 128134
rect 586260 92454 586860 127898
rect 586260 92218 586442 92454
rect 586678 92218 586860 92454
rect 586260 92134 586860 92218
rect 586260 91898 586442 92134
rect 586678 91898 586860 92134
rect 586260 56454 586860 91898
rect 586260 56218 586442 56454
rect 586678 56218 586860 56454
rect 586260 56134 586860 56218
rect 586260 55898 586442 56134
rect 586678 55898 586860 56134
rect 586260 20454 586860 55898
rect 586260 20218 586442 20454
rect 586678 20218 586860 20454
rect 586260 20134 586860 20218
rect 586260 19898 586442 20134
rect 586678 19898 586860 20134
rect 586260 -1286 586860 19898
rect 586260 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect 586260 -1606 586860 -1522
rect 586260 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect 586260 -1864 586860 -1842
rect 587200 690054 587800 706162
rect 587200 689818 587382 690054
rect 587618 689818 587800 690054
rect 587200 689734 587800 689818
rect 587200 689498 587382 689734
rect 587618 689498 587800 689734
rect 587200 654054 587800 689498
rect 587200 653818 587382 654054
rect 587618 653818 587800 654054
rect 587200 653734 587800 653818
rect 587200 653498 587382 653734
rect 587618 653498 587800 653734
rect 587200 618054 587800 653498
rect 587200 617818 587382 618054
rect 587618 617818 587800 618054
rect 587200 617734 587800 617818
rect 587200 617498 587382 617734
rect 587618 617498 587800 617734
rect 587200 582054 587800 617498
rect 587200 581818 587382 582054
rect 587618 581818 587800 582054
rect 587200 581734 587800 581818
rect 587200 581498 587382 581734
rect 587618 581498 587800 581734
rect 587200 546054 587800 581498
rect 587200 545818 587382 546054
rect 587618 545818 587800 546054
rect 587200 545734 587800 545818
rect 587200 545498 587382 545734
rect 587618 545498 587800 545734
rect 587200 510054 587800 545498
rect 587200 509818 587382 510054
rect 587618 509818 587800 510054
rect 587200 509734 587800 509818
rect 587200 509498 587382 509734
rect 587618 509498 587800 509734
rect 587200 474054 587800 509498
rect 587200 473818 587382 474054
rect 587618 473818 587800 474054
rect 587200 473734 587800 473818
rect 587200 473498 587382 473734
rect 587618 473498 587800 473734
rect 587200 438054 587800 473498
rect 587200 437818 587382 438054
rect 587618 437818 587800 438054
rect 587200 437734 587800 437818
rect 587200 437498 587382 437734
rect 587618 437498 587800 437734
rect 587200 402054 587800 437498
rect 587200 401818 587382 402054
rect 587618 401818 587800 402054
rect 587200 401734 587800 401818
rect 587200 401498 587382 401734
rect 587618 401498 587800 401734
rect 587200 366054 587800 401498
rect 587200 365818 587382 366054
rect 587618 365818 587800 366054
rect 587200 365734 587800 365818
rect 587200 365498 587382 365734
rect 587618 365498 587800 365734
rect 587200 330054 587800 365498
rect 587200 329818 587382 330054
rect 587618 329818 587800 330054
rect 587200 329734 587800 329818
rect 587200 329498 587382 329734
rect 587618 329498 587800 329734
rect 587200 294054 587800 329498
rect 587200 293818 587382 294054
rect 587618 293818 587800 294054
rect 587200 293734 587800 293818
rect 587200 293498 587382 293734
rect 587618 293498 587800 293734
rect 587200 258054 587800 293498
rect 587200 257818 587382 258054
rect 587618 257818 587800 258054
rect 587200 257734 587800 257818
rect 587200 257498 587382 257734
rect 587618 257498 587800 257734
rect 587200 222054 587800 257498
rect 587200 221818 587382 222054
rect 587618 221818 587800 222054
rect 587200 221734 587800 221818
rect 587200 221498 587382 221734
rect 587618 221498 587800 221734
rect 587200 186054 587800 221498
rect 587200 185818 587382 186054
rect 587618 185818 587800 186054
rect 587200 185734 587800 185818
rect 587200 185498 587382 185734
rect 587618 185498 587800 185734
rect 587200 150054 587800 185498
rect 587200 149818 587382 150054
rect 587618 149818 587800 150054
rect 587200 149734 587800 149818
rect 587200 149498 587382 149734
rect 587618 149498 587800 149734
rect 587200 114054 587800 149498
rect 587200 113818 587382 114054
rect 587618 113818 587800 114054
rect 587200 113734 587800 113818
rect 587200 113498 587382 113734
rect 587618 113498 587800 113734
rect 587200 78054 587800 113498
rect 587200 77818 587382 78054
rect 587618 77818 587800 78054
rect 587200 77734 587800 77818
rect 587200 77498 587382 77734
rect 587618 77498 587800 77734
rect 587200 42054 587800 77498
rect 587200 41818 587382 42054
rect 587618 41818 587800 42054
rect 587200 41734 587800 41818
rect 587200 41498 587382 41734
rect 587618 41498 587800 41734
rect 587200 6054 587800 41498
rect 587200 5818 587382 6054
rect 587618 5818 587800 6054
rect 587200 5734 587800 5818
rect 587200 5498 587382 5734
rect 587618 5498 587800 5734
rect 580404 -2462 580586 -2226
rect 580822 -2462 581004 -2226
rect 580404 -2546 581004 -2462
rect 580404 -2782 580586 -2546
rect 580822 -2782 581004 -2546
rect 580404 -3744 581004 -2782
rect 587200 -2226 587800 5498
rect 587200 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect 587200 -2546 587800 -2462
rect 587200 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect 587200 -2804 587800 -2782
rect 588140 672054 588740 707102
rect 588140 671818 588322 672054
rect 588558 671818 588740 672054
rect 588140 671734 588740 671818
rect 588140 671498 588322 671734
rect 588558 671498 588740 671734
rect 588140 636054 588740 671498
rect 588140 635818 588322 636054
rect 588558 635818 588740 636054
rect 588140 635734 588740 635818
rect 588140 635498 588322 635734
rect 588558 635498 588740 635734
rect 588140 600054 588740 635498
rect 588140 599818 588322 600054
rect 588558 599818 588740 600054
rect 588140 599734 588740 599818
rect 588140 599498 588322 599734
rect 588558 599498 588740 599734
rect 588140 564054 588740 599498
rect 588140 563818 588322 564054
rect 588558 563818 588740 564054
rect 588140 563734 588740 563818
rect 588140 563498 588322 563734
rect 588558 563498 588740 563734
rect 588140 528054 588740 563498
rect 588140 527818 588322 528054
rect 588558 527818 588740 528054
rect 588140 527734 588740 527818
rect 588140 527498 588322 527734
rect 588558 527498 588740 527734
rect 588140 492054 588740 527498
rect 588140 491818 588322 492054
rect 588558 491818 588740 492054
rect 588140 491734 588740 491818
rect 588140 491498 588322 491734
rect 588558 491498 588740 491734
rect 588140 456054 588740 491498
rect 588140 455818 588322 456054
rect 588558 455818 588740 456054
rect 588140 455734 588740 455818
rect 588140 455498 588322 455734
rect 588558 455498 588740 455734
rect 588140 420054 588740 455498
rect 588140 419818 588322 420054
rect 588558 419818 588740 420054
rect 588140 419734 588740 419818
rect 588140 419498 588322 419734
rect 588558 419498 588740 419734
rect 588140 384054 588740 419498
rect 588140 383818 588322 384054
rect 588558 383818 588740 384054
rect 588140 383734 588740 383818
rect 588140 383498 588322 383734
rect 588558 383498 588740 383734
rect 588140 348054 588740 383498
rect 588140 347818 588322 348054
rect 588558 347818 588740 348054
rect 588140 347734 588740 347818
rect 588140 347498 588322 347734
rect 588558 347498 588740 347734
rect 588140 312054 588740 347498
rect 588140 311818 588322 312054
rect 588558 311818 588740 312054
rect 588140 311734 588740 311818
rect 588140 311498 588322 311734
rect 588558 311498 588740 311734
rect 588140 276054 588740 311498
rect 588140 275818 588322 276054
rect 588558 275818 588740 276054
rect 588140 275734 588740 275818
rect 588140 275498 588322 275734
rect 588558 275498 588740 275734
rect 588140 240054 588740 275498
rect 588140 239818 588322 240054
rect 588558 239818 588740 240054
rect 588140 239734 588740 239818
rect 588140 239498 588322 239734
rect 588558 239498 588740 239734
rect 588140 204054 588740 239498
rect 588140 203818 588322 204054
rect 588558 203818 588740 204054
rect 588140 203734 588740 203818
rect 588140 203498 588322 203734
rect 588558 203498 588740 203734
rect 588140 168054 588740 203498
rect 588140 167818 588322 168054
rect 588558 167818 588740 168054
rect 588140 167734 588740 167818
rect 588140 167498 588322 167734
rect 588558 167498 588740 167734
rect 588140 132054 588740 167498
rect 588140 131818 588322 132054
rect 588558 131818 588740 132054
rect 588140 131734 588740 131818
rect 588140 131498 588322 131734
rect 588558 131498 588740 131734
rect 588140 96054 588740 131498
rect 588140 95818 588322 96054
rect 588558 95818 588740 96054
rect 588140 95734 588740 95818
rect 588140 95498 588322 95734
rect 588558 95498 588740 95734
rect 588140 60054 588740 95498
rect 588140 59818 588322 60054
rect 588558 59818 588740 60054
rect 588140 59734 588740 59818
rect 588140 59498 588322 59734
rect 588558 59498 588740 59734
rect 588140 24054 588740 59498
rect 588140 23818 588322 24054
rect 588558 23818 588740 24054
rect 588140 23734 588740 23818
rect 588140 23498 588322 23734
rect 588558 23498 588740 23734
rect 588140 -3166 588740 23498
rect 588140 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect 588140 -3486 588740 -3402
rect 588140 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect 588140 -3744 588740 -3722
rect 589080 693654 589680 708042
rect 589080 693418 589262 693654
rect 589498 693418 589680 693654
rect 589080 693334 589680 693418
rect 589080 693098 589262 693334
rect 589498 693098 589680 693334
rect 589080 657654 589680 693098
rect 589080 657418 589262 657654
rect 589498 657418 589680 657654
rect 589080 657334 589680 657418
rect 589080 657098 589262 657334
rect 589498 657098 589680 657334
rect 589080 621654 589680 657098
rect 589080 621418 589262 621654
rect 589498 621418 589680 621654
rect 589080 621334 589680 621418
rect 589080 621098 589262 621334
rect 589498 621098 589680 621334
rect 589080 585654 589680 621098
rect 589080 585418 589262 585654
rect 589498 585418 589680 585654
rect 589080 585334 589680 585418
rect 589080 585098 589262 585334
rect 589498 585098 589680 585334
rect 589080 549654 589680 585098
rect 589080 549418 589262 549654
rect 589498 549418 589680 549654
rect 589080 549334 589680 549418
rect 589080 549098 589262 549334
rect 589498 549098 589680 549334
rect 589080 513654 589680 549098
rect 589080 513418 589262 513654
rect 589498 513418 589680 513654
rect 589080 513334 589680 513418
rect 589080 513098 589262 513334
rect 589498 513098 589680 513334
rect 589080 477654 589680 513098
rect 589080 477418 589262 477654
rect 589498 477418 589680 477654
rect 589080 477334 589680 477418
rect 589080 477098 589262 477334
rect 589498 477098 589680 477334
rect 589080 441654 589680 477098
rect 589080 441418 589262 441654
rect 589498 441418 589680 441654
rect 589080 441334 589680 441418
rect 589080 441098 589262 441334
rect 589498 441098 589680 441334
rect 589080 405654 589680 441098
rect 589080 405418 589262 405654
rect 589498 405418 589680 405654
rect 589080 405334 589680 405418
rect 589080 405098 589262 405334
rect 589498 405098 589680 405334
rect 589080 369654 589680 405098
rect 589080 369418 589262 369654
rect 589498 369418 589680 369654
rect 589080 369334 589680 369418
rect 589080 369098 589262 369334
rect 589498 369098 589680 369334
rect 589080 333654 589680 369098
rect 589080 333418 589262 333654
rect 589498 333418 589680 333654
rect 589080 333334 589680 333418
rect 589080 333098 589262 333334
rect 589498 333098 589680 333334
rect 589080 297654 589680 333098
rect 589080 297418 589262 297654
rect 589498 297418 589680 297654
rect 589080 297334 589680 297418
rect 589080 297098 589262 297334
rect 589498 297098 589680 297334
rect 589080 261654 589680 297098
rect 589080 261418 589262 261654
rect 589498 261418 589680 261654
rect 589080 261334 589680 261418
rect 589080 261098 589262 261334
rect 589498 261098 589680 261334
rect 589080 225654 589680 261098
rect 589080 225418 589262 225654
rect 589498 225418 589680 225654
rect 589080 225334 589680 225418
rect 589080 225098 589262 225334
rect 589498 225098 589680 225334
rect 589080 189654 589680 225098
rect 589080 189418 589262 189654
rect 589498 189418 589680 189654
rect 589080 189334 589680 189418
rect 589080 189098 589262 189334
rect 589498 189098 589680 189334
rect 589080 153654 589680 189098
rect 589080 153418 589262 153654
rect 589498 153418 589680 153654
rect 589080 153334 589680 153418
rect 589080 153098 589262 153334
rect 589498 153098 589680 153334
rect 589080 117654 589680 153098
rect 589080 117418 589262 117654
rect 589498 117418 589680 117654
rect 589080 117334 589680 117418
rect 589080 117098 589262 117334
rect 589498 117098 589680 117334
rect 589080 81654 589680 117098
rect 589080 81418 589262 81654
rect 589498 81418 589680 81654
rect 589080 81334 589680 81418
rect 589080 81098 589262 81334
rect 589498 81098 589680 81334
rect 589080 45654 589680 81098
rect 589080 45418 589262 45654
rect 589498 45418 589680 45654
rect 589080 45334 589680 45418
rect 589080 45098 589262 45334
rect 589498 45098 589680 45334
rect 589080 9654 589680 45098
rect 589080 9418 589262 9654
rect 589498 9418 589680 9654
rect 589080 9334 589680 9418
rect 589080 9098 589262 9334
rect 589498 9098 589680 9334
rect 589080 -4106 589680 9098
rect 589080 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect 589080 -4426 589680 -4342
rect 589080 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect 589080 -4684 589680 -4662
rect 590020 675654 590620 708982
rect 590020 675418 590202 675654
rect 590438 675418 590620 675654
rect 590020 675334 590620 675418
rect 590020 675098 590202 675334
rect 590438 675098 590620 675334
rect 590020 639654 590620 675098
rect 590020 639418 590202 639654
rect 590438 639418 590620 639654
rect 590020 639334 590620 639418
rect 590020 639098 590202 639334
rect 590438 639098 590620 639334
rect 590020 603654 590620 639098
rect 590020 603418 590202 603654
rect 590438 603418 590620 603654
rect 590020 603334 590620 603418
rect 590020 603098 590202 603334
rect 590438 603098 590620 603334
rect 590020 567654 590620 603098
rect 590020 567418 590202 567654
rect 590438 567418 590620 567654
rect 590020 567334 590620 567418
rect 590020 567098 590202 567334
rect 590438 567098 590620 567334
rect 590020 531654 590620 567098
rect 590020 531418 590202 531654
rect 590438 531418 590620 531654
rect 590020 531334 590620 531418
rect 590020 531098 590202 531334
rect 590438 531098 590620 531334
rect 590020 495654 590620 531098
rect 590020 495418 590202 495654
rect 590438 495418 590620 495654
rect 590020 495334 590620 495418
rect 590020 495098 590202 495334
rect 590438 495098 590620 495334
rect 590020 459654 590620 495098
rect 590020 459418 590202 459654
rect 590438 459418 590620 459654
rect 590020 459334 590620 459418
rect 590020 459098 590202 459334
rect 590438 459098 590620 459334
rect 590020 423654 590620 459098
rect 590020 423418 590202 423654
rect 590438 423418 590620 423654
rect 590020 423334 590620 423418
rect 590020 423098 590202 423334
rect 590438 423098 590620 423334
rect 590020 387654 590620 423098
rect 590020 387418 590202 387654
rect 590438 387418 590620 387654
rect 590020 387334 590620 387418
rect 590020 387098 590202 387334
rect 590438 387098 590620 387334
rect 590020 351654 590620 387098
rect 590020 351418 590202 351654
rect 590438 351418 590620 351654
rect 590020 351334 590620 351418
rect 590020 351098 590202 351334
rect 590438 351098 590620 351334
rect 590020 315654 590620 351098
rect 590020 315418 590202 315654
rect 590438 315418 590620 315654
rect 590020 315334 590620 315418
rect 590020 315098 590202 315334
rect 590438 315098 590620 315334
rect 590020 279654 590620 315098
rect 590020 279418 590202 279654
rect 590438 279418 590620 279654
rect 590020 279334 590620 279418
rect 590020 279098 590202 279334
rect 590438 279098 590620 279334
rect 590020 243654 590620 279098
rect 590020 243418 590202 243654
rect 590438 243418 590620 243654
rect 590020 243334 590620 243418
rect 590020 243098 590202 243334
rect 590438 243098 590620 243334
rect 590020 207654 590620 243098
rect 590020 207418 590202 207654
rect 590438 207418 590620 207654
rect 590020 207334 590620 207418
rect 590020 207098 590202 207334
rect 590438 207098 590620 207334
rect 590020 171654 590620 207098
rect 590020 171418 590202 171654
rect 590438 171418 590620 171654
rect 590020 171334 590620 171418
rect 590020 171098 590202 171334
rect 590438 171098 590620 171334
rect 590020 135654 590620 171098
rect 590020 135418 590202 135654
rect 590438 135418 590620 135654
rect 590020 135334 590620 135418
rect 590020 135098 590202 135334
rect 590438 135098 590620 135334
rect 590020 99654 590620 135098
rect 590020 99418 590202 99654
rect 590438 99418 590620 99654
rect 590020 99334 590620 99418
rect 590020 99098 590202 99334
rect 590438 99098 590620 99334
rect 590020 63654 590620 99098
rect 590020 63418 590202 63654
rect 590438 63418 590620 63654
rect 590020 63334 590620 63418
rect 590020 63098 590202 63334
rect 590438 63098 590620 63334
rect 590020 27654 590620 63098
rect 590020 27418 590202 27654
rect 590438 27418 590620 27654
rect 590020 27334 590620 27418
rect 590020 27098 590202 27334
rect 590438 27098 590620 27334
rect 590020 -5046 590620 27098
rect 590020 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect 590020 -5366 590620 -5282
rect 590020 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect 590020 -5624 590620 -5602
rect 590960 697254 591560 709922
rect 590960 697018 591142 697254
rect 591378 697018 591560 697254
rect 590960 696934 591560 697018
rect 590960 696698 591142 696934
rect 591378 696698 591560 696934
rect 590960 661254 591560 696698
rect 590960 661018 591142 661254
rect 591378 661018 591560 661254
rect 590960 660934 591560 661018
rect 590960 660698 591142 660934
rect 591378 660698 591560 660934
rect 590960 625254 591560 660698
rect 590960 625018 591142 625254
rect 591378 625018 591560 625254
rect 590960 624934 591560 625018
rect 590960 624698 591142 624934
rect 591378 624698 591560 624934
rect 590960 589254 591560 624698
rect 590960 589018 591142 589254
rect 591378 589018 591560 589254
rect 590960 588934 591560 589018
rect 590960 588698 591142 588934
rect 591378 588698 591560 588934
rect 590960 553254 591560 588698
rect 590960 553018 591142 553254
rect 591378 553018 591560 553254
rect 590960 552934 591560 553018
rect 590960 552698 591142 552934
rect 591378 552698 591560 552934
rect 590960 517254 591560 552698
rect 590960 517018 591142 517254
rect 591378 517018 591560 517254
rect 590960 516934 591560 517018
rect 590960 516698 591142 516934
rect 591378 516698 591560 516934
rect 590960 481254 591560 516698
rect 590960 481018 591142 481254
rect 591378 481018 591560 481254
rect 590960 480934 591560 481018
rect 590960 480698 591142 480934
rect 591378 480698 591560 480934
rect 590960 445254 591560 480698
rect 590960 445018 591142 445254
rect 591378 445018 591560 445254
rect 590960 444934 591560 445018
rect 590960 444698 591142 444934
rect 591378 444698 591560 444934
rect 590960 409254 591560 444698
rect 590960 409018 591142 409254
rect 591378 409018 591560 409254
rect 590960 408934 591560 409018
rect 590960 408698 591142 408934
rect 591378 408698 591560 408934
rect 590960 373254 591560 408698
rect 590960 373018 591142 373254
rect 591378 373018 591560 373254
rect 590960 372934 591560 373018
rect 590960 372698 591142 372934
rect 591378 372698 591560 372934
rect 590960 337254 591560 372698
rect 590960 337018 591142 337254
rect 591378 337018 591560 337254
rect 590960 336934 591560 337018
rect 590960 336698 591142 336934
rect 591378 336698 591560 336934
rect 590960 301254 591560 336698
rect 590960 301018 591142 301254
rect 591378 301018 591560 301254
rect 590960 300934 591560 301018
rect 590960 300698 591142 300934
rect 591378 300698 591560 300934
rect 590960 265254 591560 300698
rect 590960 265018 591142 265254
rect 591378 265018 591560 265254
rect 590960 264934 591560 265018
rect 590960 264698 591142 264934
rect 591378 264698 591560 264934
rect 590960 229254 591560 264698
rect 590960 229018 591142 229254
rect 591378 229018 591560 229254
rect 590960 228934 591560 229018
rect 590960 228698 591142 228934
rect 591378 228698 591560 228934
rect 590960 193254 591560 228698
rect 590960 193018 591142 193254
rect 591378 193018 591560 193254
rect 590960 192934 591560 193018
rect 590960 192698 591142 192934
rect 591378 192698 591560 192934
rect 590960 157254 591560 192698
rect 590960 157018 591142 157254
rect 591378 157018 591560 157254
rect 590960 156934 591560 157018
rect 590960 156698 591142 156934
rect 591378 156698 591560 156934
rect 590960 121254 591560 156698
rect 590960 121018 591142 121254
rect 591378 121018 591560 121254
rect 590960 120934 591560 121018
rect 590960 120698 591142 120934
rect 591378 120698 591560 120934
rect 590960 85254 591560 120698
rect 590960 85018 591142 85254
rect 591378 85018 591560 85254
rect 590960 84934 591560 85018
rect 590960 84698 591142 84934
rect 591378 84698 591560 84934
rect 590960 49254 591560 84698
rect 590960 49018 591142 49254
rect 591378 49018 591560 49254
rect 590960 48934 591560 49018
rect 590960 48698 591142 48934
rect 591378 48698 591560 48934
rect 590960 13254 591560 48698
rect 590960 13018 591142 13254
rect 591378 13018 591560 13254
rect 590960 12934 591560 13018
rect 590960 12698 591142 12934
rect 591378 12698 591560 12934
rect 590960 -5986 591560 12698
rect 590960 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect 590960 -6306 591560 -6222
rect 590960 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect 590960 -6564 591560 -6542
rect 591900 679254 592500 710862
rect 591900 679018 592082 679254
rect 592318 679018 592500 679254
rect 591900 678934 592500 679018
rect 591900 678698 592082 678934
rect 592318 678698 592500 678934
rect 591900 643254 592500 678698
rect 591900 643018 592082 643254
rect 592318 643018 592500 643254
rect 591900 642934 592500 643018
rect 591900 642698 592082 642934
rect 592318 642698 592500 642934
rect 591900 607254 592500 642698
rect 591900 607018 592082 607254
rect 592318 607018 592500 607254
rect 591900 606934 592500 607018
rect 591900 606698 592082 606934
rect 592318 606698 592500 606934
rect 591900 571254 592500 606698
rect 591900 571018 592082 571254
rect 592318 571018 592500 571254
rect 591900 570934 592500 571018
rect 591900 570698 592082 570934
rect 592318 570698 592500 570934
rect 591900 535254 592500 570698
rect 591900 535018 592082 535254
rect 592318 535018 592500 535254
rect 591900 534934 592500 535018
rect 591900 534698 592082 534934
rect 592318 534698 592500 534934
rect 591900 499254 592500 534698
rect 591900 499018 592082 499254
rect 592318 499018 592500 499254
rect 591900 498934 592500 499018
rect 591900 498698 592082 498934
rect 592318 498698 592500 498934
rect 591900 463254 592500 498698
rect 591900 463018 592082 463254
rect 592318 463018 592500 463254
rect 591900 462934 592500 463018
rect 591900 462698 592082 462934
rect 592318 462698 592500 462934
rect 591900 427254 592500 462698
rect 591900 427018 592082 427254
rect 592318 427018 592500 427254
rect 591900 426934 592500 427018
rect 591900 426698 592082 426934
rect 592318 426698 592500 426934
rect 591900 391254 592500 426698
rect 591900 391018 592082 391254
rect 592318 391018 592500 391254
rect 591900 390934 592500 391018
rect 591900 390698 592082 390934
rect 592318 390698 592500 390934
rect 591900 355254 592500 390698
rect 591900 355018 592082 355254
rect 592318 355018 592500 355254
rect 591900 354934 592500 355018
rect 591900 354698 592082 354934
rect 592318 354698 592500 354934
rect 591900 319254 592500 354698
rect 591900 319018 592082 319254
rect 592318 319018 592500 319254
rect 591900 318934 592500 319018
rect 591900 318698 592082 318934
rect 592318 318698 592500 318934
rect 591900 283254 592500 318698
rect 591900 283018 592082 283254
rect 592318 283018 592500 283254
rect 591900 282934 592500 283018
rect 591900 282698 592082 282934
rect 592318 282698 592500 282934
rect 591900 247254 592500 282698
rect 591900 247018 592082 247254
rect 592318 247018 592500 247254
rect 591900 246934 592500 247018
rect 591900 246698 592082 246934
rect 592318 246698 592500 246934
rect 591900 211254 592500 246698
rect 591900 211018 592082 211254
rect 592318 211018 592500 211254
rect 591900 210934 592500 211018
rect 591900 210698 592082 210934
rect 592318 210698 592500 210934
rect 591900 175254 592500 210698
rect 591900 175018 592082 175254
rect 592318 175018 592500 175254
rect 591900 174934 592500 175018
rect 591900 174698 592082 174934
rect 592318 174698 592500 174934
rect 591900 139254 592500 174698
rect 591900 139018 592082 139254
rect 592318 139018 592500 139254
rect 591900 138934 592500 139018
rect 591900 138698 592082 138934
rect 592318 138698 592500 138934
rect 591900 103254 592500 138698
rect 591900 103018 592082 103254
rect 592318 103018 592500 103254
rect 591900 102934 592500 103018
rect 591900 102698 592082 102934
rect 592318 102698 592500 102934
rect 591900 67254 592500 102698
rect 591900 67018 592082 67254
rect 592318 67018 592500 67254
rect 591900 66934 592500 67018
rect 591900 66698 592082 66934
rect 592318 66698 592500 66934
rect 591900 31254 592500 66698
rect 591900 31018 592082 31254
rect 592318 31018 592500 31254
rect 591900 30934 592500 31018
rect 591900 30698 592082 30934
rect 592318 30698 592500 30934
rect 569604 -7162 569786 -6926
rect 570022 -7162 570204 -6926
rect 569604 -7246 570204 -7162
rect 569604 -7482 569786 -7246
rect 570022 -7482 570204 -7246
rect 569604 -7504 570204 -7482
rect 591900 -6926 592500 30698
rect 591900 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect 591900 -7246 592500 -7162
rect 591900 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect 591900 -7504 592500 -7482
<< via4 >>
rect -8394 711182 -8158 711418
rect -8394 710862 -8158 711098
rect -8394 679018 -8158 679254
rect -8394 678698 -8158 678934
rect -8394 643018 -8158 643254
rect -8394 642698 -8158 642934
rect -8394 607018 -8158 607254
rect -8394 606698 -8158 606934
rect -8394 571018 -8158 571254
rect -8394 570698 -8158 570934
rect -8394 535018 -8158 535254
rect -8394 534698 -8158 534934
rect -8394 499018 -8158 499254
rect -8394 498698 -8158 498934
rect -8394 463018 -8158 463254
rect -8394 462698 -8158 462934
rect -8394 427018 -8158 427254
rect -8394 426698 -8158 426934
rect -8394 391018 -8158 391254
rect -8394 390698 -8158 390934
rect -8394 355018 -8158 355254
rect -8394 354698 -8158 354934
rect -8394 319018 -8158 319254
rect -8394 318698 -8158 318934
rect -8394 283018 -8158 283254
rect -8394 282698 -8158 282934
rect -8394 247018 -8158 247254
rect -8394 246698 -8158 246934
rect -8394 211018 -8158 211254
rect -8394 210698 -8158 210934
rect -8394 175018 -8158 175254
rect -8394 174698 -8158 174934
rect -8394 139018 -8158 139254
rect -8394 138698 -8158 138934
rect -8394 103018 -8158 103254
rect -8394 102698 -8158 102934
rect -8394 67018 -8158 67254
rect -8394 66698 -8158 66934
rect -8394 31018 -8158 31254
rect -8394 30698 -8158 30934
rect -7454 710242 -7218 710478
rect -7454 709922 -7218 710158
rect 11786 710242 12022 710478
rect 11786 709922 12022 710158
rect -7454 697018 -7218 697254
rect -7454 696698 -7218 696934
rect -7454 661018 -7218 661254
rect -7454 660698 -7218 660934
rect -7454 625018 -7218 625254
rect -7454 624698 -7218 624934
rect -7454 589018 -7218 589254
rect -7454 588698 -7218 588934
rect -7454 553018 -7218 553254
rect -7454 552698 -7218 552934
rect -7454 517018 -7218 517254
rect -7454 516698 -7218 516934
rect -7454 481018 -7218 481254
rect -7454 480698 -7218 480934
rect -7454 445018 -7218 445254
rect -7454 444698 -7218 444934
rect -7454 409018 -7218 409254
rect -7454 408698 -7218 408934
rect -7454 373018 -7218 373254
rect -7454 372698 -7218 372934
rect -7454 337018 -7218 337254
rect -7454 336698 -7218 336934
rect -7454 301018 -7218 301254
rect -7454 300698 -7218 300934
rect -7454 265018 -7218 265254
rect -7454 264698 -7218 264934
rect -7454 229018 -7218 229254
rect -7454 228698 -7218 228934
rect -7454 193018 -7218 193254
rect -7454 192698 -7218 192934
rect -7454 157018 -7218 157254
rect -7454 156698 -7218 156934
rect -7454 121018 -7218 121254
rect -7454 120698 -7218 120934
rect -7454 85018 -7218 85254
rect -7454 84698 -7218 84934
rect -7454 49018 -7218 49254
rect -7454 48698 -7218 48934
rect -7454 13018 -7218 13254
rect -7454 12698 -7218 12934
rect -6514 709302 -6278 709538
rect -6514 708982 -6278 709218
rect -6514 675418 -6278 675654
rect -6514 675098 -6278 675334
rect -6514 639418 -6278 639654
rect -6514 639098 -6278 639334
rect -6514 603418 -6278 603654
rect -6514 603098 -6278 603334
rect -6514 567418 -6278 567654
rect -6514 567098 -6278 567334
rect -6514 531418 -6278 531654
rect -6514 531098 -6278 531334
rect -6514 495418 -6278 495654
rect -6514 495098 -6278 495334
rect -6514 459418 -6278 459654
rect -6514 459098 -6278 459334
rect -6514 423418 -6278 423654
rect -6514 423098 -6278 423334
rect -6514 387418 -6278 387654
rect -6514 387098 -6278 387334
rect -6514 351418 -6278 351654
rect -6514 351098 -6278 351334
rect -6514 315418 -6278 315654
rect -6514 315098 -6278 315334
rect -6514 279418 -6278 279654
rect -6514 279098 -6278 279334
rect -6514 243418 -6278 243654
rect -6514 243098 -6278 243334
rect -6514 207418 -6278 207654
rect -6514 207098 -6278 207334
rect -6514 171418 -6278 171654
rect -6514 171098 -6278 171334
rect -6514 135418 -6278 135654
rect -6514 135098 -6278 135334
rect -6514 99418 -6278 99654
rect -6514 99098 -6278 99334
rect -6514 63418 -6278 63654
rect -6514 63098 -6278 63334
rect -6514 27418 -6278 27654
rect -6514 27098 -6278 27334
rect -5574 708362 -5338 708598
rect -5574 708042 -5338 708278
rect 8186 708362 8422 708598
rect 8186 708042 8422 708278
rect -5574 693418 -5338 693654
rect -5574 693098 -5338 693334
rect -5574 657418 -5338 657654
rect -5574 657098 -5338 657334
rect -5574 621418 -5338 621654
rect -5574 621098 -5338 621334
rect -5574 585418 -5338 585654
rect -5574 585098 -5338 585334
rect -5574 549418 -5338 549654
rect -5574 549098 -5338 549334
rect -5574 513418 -5338 513654
rect -5574 513098 -5338 513334
rect -5574 477418 -5338 477654
rect -5574 477098 -5338 477334
rect -5574 441418 -5338 441654
rect -5574 441098 -5338 441334
rect -5574 405418 -5338 405654
rect -5574 405098 -5338 405334
rect -5574 369418 -5338 369654
rect -5574 369098 -5338 369334
rect -5574 333418 -5338 333654
rect -5574 333098 -5338 333334
rect -5574 297418 -5338 297654
rect -5574 297098 -5338 297334
rect -5574 261418 -5338 261654
rect -5574 261098 -5338 261334
rect -5574 225418 -5338 225654
rect -5574 225098 -5338 225334
rect -5574 189418 -5338 189654
rect -5574 189098 -5338 189334
rect -5574 153418 -5338 153654
rect -5574 153098 -5338 153334
rect -5574 117418 -5338 117654
rect -5574 117098 -5338 117334
rect -5574 81418 -5338 81654
rect -5574 81098 -5338 81334
rect -5574 45418 -5338 45654
rect -5574 45098 -5338 45334
rect -5574 9418 -5338 9654
rect -5574 9098 -5338 9334
rect -4634 707422 -4398 707658
rect -4634 707102 -4398 707338
rect -4634 671818 -4398 672054
rect -4634 671498 -4398 671734
rect -4634 635818 -4398 636054
rect -4634 635498 -4398 635734
rect -4634 599818 -4398 600054
rect -4634 599498 -4398 599734
rect -4634 563818 -4398 564054
rect -4634 563498 -4398 563734
rect -4634 527818 -4398 528054
rect -4634 527498 -4398 527734
rect -4634 491818 -4398 492054
rect -4634 491498 -4398 491734
rect -4634 455818 -4398 456054
rect -4634 455498 -4398 455734
rect -4634 419818 -4398 420054
rect -4634 419498 -4398 419734
rect -4634 383818 -4398 384054
rect -4634 383498 -4398 383734
rect -4634 347818 -4398 348054
rect -4634 347498 -4398 347734
rect -4634 311818 -4398 312054
rect -4634 311498 -4398 311734
rect -4634 275818 -4398 276054
rect -4634 275498 -4398 275734
rect -4634 239818 -4398 240054
rect -4634 239498 -4398 239734
rect -4634 203818 -4398 204054
rect -4634 203498 -4398 203734
rect -4634 167818 -4398 168054
rect -4634 167498 -4398 167734
rect -4634 131818 -4398 132054
rect -4634 131498 -4398 131734
rect -4634 95818 -4398 96054
rect -4634 95498 -4398 95734
rect -4634 59818 -4398 60054
rect -4634 59498 -4398 59734
rect -4634 23818 -4398 24054
rect -4634 23498 -4398 23734
rect -3694 706482 -3458 706718
rect -3694 706162 -3458 706398
rect 4586 706482 4822 706718
rect 4586 706162 4822 706398
rect -3694 689818 -3458 690054
rect -3694 689498 -3458 689734
rect -3694 653818 -3458 654054
rect -3694 653498 -3458 653734
rect -3694 617818 -3458 618054
rect -3694 617498 -3458 617734
rect -3694 581818 -3458 582054
rect -3694 581498 -3458 581734
rect -3694 545818 -3458 546054
rect -3694 545498 -3458 545734
rect -3694 509818 -3458 510054
rect -3694 509498 -3458 509734
rect -3694 473818 -3458 474054
rect -3694 473498 -3458 473734
rect -3694 437818 -3458 438054
rect -3694 437498 -3458 437734
rect -3694 401818 -3458 402054
rect -3694 401498 -3458 401734
rect -3694 365818 -3458 366054
rect -3694 365498 -3458 365734
rect -3694 329818 -3458 330054
rect -3694 329498 -3458 329734
rect -3694 293818 -3458 294054
rect -3694 293498 -3458 293734
rect -3694 257818 -3458 258054
rect -3694 257498 -3458 257734
rect -3694 221818 -3458 222054
rect -3694 221498 -3458 221734
rect -3694 185818 -3458 186054
rect -3694 185498 -3458 185734
rect -3694 149818 -3458 150054
rect -3694 149498 -3458 149734
rect -3694 113818 -3458 114054
rect -3694 113498 -3458 113734
rect -3694 77818 -3458 78054
rect -3694 77498 -3458 77734
rect -3694 41818 -3458 42054
rect -3694 41498 -3458 41734
rect -3694 5818 -3458 6054
rect -3694 5498 -3458 5734
rect -2754 705542 -2518 705778
rect -2754 705222 -2518 705458
rect -2754 668218 -2518 668454
rect -2754 667898 -2518 668134
rect -2754 632218 -2518 632454
rect -2754 631898 -2518 632134
rect -2754 596218 -2518 596454
rect -2754 595898 -2518 596134
rect -2754 560218 -2518 560454
rect -2754 559898 -2518 560134
rect -2754 524218 -2518 524454
rect -2754 523898 -2518 524134
rect -2754 488218 -2518 488454
rect -2754 487898 -2518 488134
rect -2754 452218 -2518 452454
rect -2754 451898 -2518 452134
rect -2754 416218 -2518 416454
rect -2754 415898 -2518 416134
rect -2754 380218 -2518 380454
rect -2754 379898 -2518 380134
rect -2754 344218 -2518 344454
rect -2754 343898 -2518 344134
rect -2754 308218 -2518 308454
rect -2754 307898 -2518 308134
rect -2754 272218 -2518 272454
rect -2754 271898 -2518 272134
rect -2754 236218 -2518 236454
rect -2754 235898 -2518 236134
rect -2754 200218 -2518 200454
rect -2754 199898 -2518 200134
rect -2754 164218 -2518 164454
rect -2754 163898 -2518 164134
rect -2754 128218 -2518 128454
rect -2754 127898 -2518 128134
rect -2754 92218 -2518 92454
rect -2754 91898 -2518 92134
rect -2754 56218 -2518 56454
rect -2754 55898 -2518 56134
rect -2754 20218 -2518 20454
rect -2754 19898 -2518 20134
rect -1814 704602 -1578 704838
rect -1814 704282 -1578 704518
rect -1814 686218 -1578 686454
rect -1814 685898 -1578 686134
rect -1814 650218 -1578 650454
rect -1814 649898 -1578 650134
rect -1814 614218 -1578 614454
rect -1814 613898 -1578 614134
rect -1814 578218 -1578 578454
rect -1814 577898 -1578 578134
rect -1814 542218 -1578 542454
rect -1814 541898 -1578 542134
rect -1814 506218 -1578 506454
rect -1814 505898 -1578 506134
rect -1814 470218 -1578 470454
rect -1814 469898 -1578 470134
rect -1814 434218 -1578 434454
rect -1814 433898 -1578 434134
rect -1814 398218 -1578 398454
rect -1814 397898 -1578 398134
rect -1814 362218 -1578 362454
rect -1814 361898 -1578 362134
rect -1814 326218 -1578 326454
rect -1814 325898 -1578 326134
rect -1814 290218 -1578 290454
rect -1814 289898 -1578 290134
rect -1814 254218 -1578 254454
rect -1814 253898 -1578 254134
rect -1814 218218 -1578 218454
rect -1814 217898 -1578 218134
rect -1814 182218 -1578 182454
rect -1814 181898 -1578 182134
rect -1814 146218 -1578 146454
rect -1814 145898 -1578 146134
rect -1814 110218 -1578 110454
rect -1814 109898 -1578 110134
rect -1814 74218 -1578 74454
rect -1814 73898 -1578 74134
rect -1814 38218 -1578 38454
rect -1814 37898 -1578 38134
rect -1814 2218 -1578 2454
rect -1814 1898 -1578 2134
rect -1814 -582 -1578 -346
rect -1814 -902 -1578 -666
rect 986 704602 1222 704838
rect 986 704282 1222 704518
rect 986 686218 1222 686454
rect 986 685898 1222 686134
rect 986 650218 1222 650454
rect 986 649898 1222 650134
rect 986 614218 1222 614454
rect 986 613898 1222 614134
rect 986 578218 1222 578454
rect 986 577898 1222 578134
rect 986 542218 1222 542454
rect 986 541898 1222 542134
rect 986 506218 1222 506454
rect 986 505898 1222 506134
rect 986 470218 1222 470454
rect 986 469898 1222 470134
rect 986 434218 1222 434454
rect 986 433898 1222 434134
rect 986 398218 1222 398454
rect 986 397898 1222 398134
rect 986 362218 1222 362454
rect 986 361898 1222 362134
rect 986 326218 1222 326454
rect 986 325898 1222 326134
rect 986 290218 1222 290454
rect 986 289898 1222 290134
rect 986 254218 1222 254454
rect 986 253898 1222 254134
rect 986 218218 1222 218454
rect 986 217898 1222 218134
rect 986 182218 1222 182454
rect 986 181898 1222 182134
rect 986 146218 1222 146454
rect 986 145898 1222 146134
rect 986 110218 1222 110454
rect 986 109898 1222 110134
rect 986 74218 1222 74454
rect 986 73898 1222 74134
rect 986 38218 1222 38454
rect 986 37898 1222 38134
rect 986 2218 1222 2454
rect 986 1898 1222 2134
rect 986 -582 1222 -346
rect 986 -902 1222 -666
rect -2754 -1522 -2518 -1286
rect -2754 -1842 -2518 -1606
rect 4586 689818 4822 690054
rect 4586 689498 4822 689734
rect 4586 653818 4822 654054
rect 4586 653498 4822 653734
rect 4586 617818 4822 618054
rect 4586 617498 4822 617734
rect 4586 581818 4822 582054
rect 4586 581498 4822 581734
rect 4586 545818 4822 546054
rect 4586 545498 4822 545734
rect 4586 509818 4822 510054
rect 4586 509498 4822 509734
rect 4586 473818 4822 474054
rect 4586 473498 4822 473734
rect 4586 437818 4822 438054
rect 4586 437498 4822 437734
rect 4586 401818 4822 402054
rect 4586 401498 4822 401734
rect 4586 365818 4822 366054
rect 4586 365498 4822 365734
rect 4586 329818 4822 330054
rect 4586 329498 4822 329734
rect 4586 293818 4822 294054
rect 4586 293498 4822 293734
rect 4586 257818 4822 258054
rect 4586 257498 4822 257734
rect 4586 221818 4822 222054
rect 4586 221498 4822 221734
rect 4586 185818 4822 186054
rect 4586 185498 4822 185734
rect 4586 149818 4822 150054
rect 4586 149498 4822 149734
rect 4586 113818 4822 114054
rect 4586 113498 4822 113734
rect 4586 77818 4822 78054
rect 4586 77498 4822 77734
rect 4586 41818 4822 42054
rect 4586 41498 4822 41734
rect 4586 5818 4822 6054
rect 4586 5498 4822 5734
rect -3694 -2462 -3458 -2226
rect -3694 -2782 -3458 -2546
rect 4586 -2462 4822 -2226
rect 4586 -2782 4822 -2546
rect -4634 -3402 -4398 -3166
rect -4634 -3722 -4398 -3486
rect 8186 693418 8422 693654
rect 8186 693098 8422 693334
rect 8186 657418 8422 657654
rect 8186 657098 8422 657334
rect 8186 621418 8422 621654
rect 8186 621098 8422 621334
rect 8186 585418 8422 585654
rect 8186 585098 8422 585334
rect 8186 549418 8422 549654
rect 8186 549098 8422 549334
rect 8186 513418 8422 513654
rect 8186 513098 8422 513334
rect 8186 477418 8422 477654
rect 8186 477098 8422 477334
rect 8186 441418 8422 441654
rect 8186 441098 8422 441334
rect 8186 405418 8422 405654
rect 8186 405098 8422 405334
rect 8186 369418 8422 369654
rect 8186 369098 8422 369334
rect 8186 333418 8422 333654
rect 8186 333098 8422 333334
rect 8186 297418 8422 297654
rect 8186 297098 8422 297334
rect 8186 261418 8422 261654
rect 8186 261098 8422 261334
rect 8186 225418 8422 225654
rect 8186 225098 8422 225334
rect 8186 189418 8422 189654
rect 8186 189098 8422 189334
rect 8186 153418 8422 153654
rect 8186 153098 8422 153334
rect 8186 117418 8422 117654
rect 8186 117098 8422 117334
rect 8186 81418 8422 81654
rect 8186 81098 8422 81334
rect 8186 45418 8422 45654
rect 8186 45098 8422 45334
rect 8186 9418 8422 9654
rect 8186 9098 8422 9334
rect -5574 -4342 -5338 -4106
rect -5574 -4662 -5338 -4426
rect 8186 -4342 8422 -4106
rect 8186 -4662 8422 -4426
rect -6514 -5282 -6278 -5046
rect -6514 -5602 -6278 -5366
rect 29786 711182 30022 711418
rect 29786 710862 30022 711098
rect 26186 709302 26422 709538
rect 26186 708982 26422 709218
rect 22586 707422 22822 707658
rect 22586 707102 22822 707338
rect 11786 697018 12022 697254
rect 11786 696698 12022 696934
rect 11786 661018 12022 661254
rect 11786 660698 12022 660934
rect 11786 625018 12022 625254
rect 11786 624698 12022 624934
rect 11786 589018 12022 589254
rect 11786 588698 12022 588934
rect 11786 553018 12022 553254
rect 11786 552698 12022 552934
rect 11786 517018 12022 517254
rect 11786 516698 12022 516934
rect 11786 481018 12022 481254
rect 11786 480698 12022 480934
rect 11786 445018 12022 445254
rect 11786 444698 12022 444934
rect 11786 409018 12022 409254
rect 11786 408698 12022 408934
rect 11786 373018 12022 373254
rect 11786 372698 12022 372934
rect 11786 337018 12022 337254
rect 11786 336698 12022 336934
rect 11786 301018 12022 301254
rect 11786 300698 12022 300934
rect 11786 265018 12022 265254
rect 11786 264698 12022 264934
rect 11786 229018 12022 229254
rect 11786 228698 12022 228934
rect 11786 193018 12022 193254
rect 11786 192698 12022 192934
rect 11786 157018 12022 157254
rect 11786 156698 12022 156934
rect 11786 121018 12022 121254
rect 11786 120698 12022 120934
rect 11786 85018 12022 85254
rect 11786 84698 12022 84934
rect 11786 49018 12022 49254
rect 11786 48698 12022 48934
rect 11786 13018 12022 13254
rect 11786 12698 12022 12934
rect -7454 -6222 -7218 -5986
rect -7454 -6542 -7218 -6306
rect 18986 705542 19222 705778
rect 18986 705222 19222 705458
rect 18986 668218 19222 668454
rect 18986 667898 19222 668134
rect 18986 632218 19222 632454
rect 18986 631898 19222 632134
rect 18986 596218 19222 596454
rect 18986 595898 19222 596134
rect 18986 560218 19222 560454
rect 18986 559898 19222 560134
rect 18986 524218 19222 524454
rect 18986 523898 19222 524134
rect 18986 488218 19222 488454
rect 18986 487898 19222 488134
rect 18986 452218 19222 452454
rect 18986 451898 19222 452134
rect 18986 416218 19222 416454
rect 18986 415898 19222 416134
rect 18986 380218 19222 380454
rect 18986 379898 19222 380134
rect 18986 344218 19222 344454
rect 18986 343898 19222 344134
rect 18986 308218 19222 308454
rect 18986 307898 19222 308134
rect 18986 272218 19222 272454
rect 18986 271898 19222 272134
rect 18986 236218 19222 236454
rect 18986 235898 19222 236134
rect 18986 200218 19222 200454
rect 18986 199898 19222 200134
rect 18986 164218 19222 164454
rect 18986 163898 19222 164134
rect 18986 128218 19222 128454
rect 18986 127898 19222 128134
rect 18986 92218 19222 92454
rect 18986 91898 19222 92134
rect 18986 56218 19222 56454
rect 18986 55898 19222 56134
rect 18986 20218 19222 20454
rect 18986 19898 19222 20134
rect 18986 -1522 19222 -1286
rect 18986 -1842 19222 -1606
rect 22586 671818 22822 672054
rect 22586 671498 22822 671734
rect 22586 635818 22822 636054
rect 22586 635498 22822 635734
rect 22586 599818 22822 600054
rect 22586 599498 22822 599734
rect 22586 563818 22822 564054
rect 22586 563498 22822 563734
rect 22586 527818 22822 528054
rect 22586 527498 22822 527734
rect 22586 491818 22822 492054
rect 22586 491498 22822 491734
rect 22586 455818 22822 456054
rect 22586 455498 22822 455734
rect 22586 419818 22822 420054
rect 22586 419498 22822 419734
rect 22586 383818 22822 384054
rect 22586 383498 22822 383734
rect 22586 347818 22822 348054
rect 22586 347498 22822 347734
rect 22586 311818 22822 312054
rect 22586 311498 22822 311734
rect 22586 275818 22822 276054
rect 22586 275498 22822 275734
rect 22586 239818 22822 240054
rect 22586 239498 22822 239734
rect 22586 203818 22822 204054
rect 22586 203498 22822 203734
rect 22586 167818 22822 168054
rect 22586 167498 22822 167734
rect 22586 131818 22822 132054
rect 22586 131498 22822 131734
rect 22586 95818 22822 96054
rect 22586 95498 22822 95734
rect 22586 59818 22822 60054
rect 22586 59498 22822 59734
rect 22586 23818 22822 24054
rect 22586 23498 22822 23734
rect 22586 -3402 22822 -3166
rect 22586 -3722 22822 -3486
rect 26186 675418 26422 675654
rect 26186 675098 26422 675334
rect 26186 639418 26422 639654
rect 26186 639098 26422 639334
rect 26186 603418 26422 603654
rect 26186 603098 26422 603334
rect 26186 567418 26422 567654
rect 26186 567098 26422 567334
rect 26186 531418 26422 531654
rect 26186 531098 26422 531334
rect 26186 495418 26422 495654
rect 26186 495098 26422 495334
rect 26186 459418 26422 459654
rect 26186 459098 26422 459334
rect 26186 423418 26422 423654
rect 26186 423098 26422 423334
rect 26186 387418 26422 387654
rect 26186 387098 26422 387334
rect 26186 351418 26422 351654
rect 26186 351098 26422 351334
rect 26186 315418 26422 315654
rect 26186 315098 26422 315334
rect 26186 279418 26422 279654
rect 26186 279098 26422 279334
rect 26186 243418 26422 243654
rect 26186 243098 26422 243334
rect 26186 207418 26422 207654
rect 26186 207098 26422 207334
rect 26186 171418 26422 171654
rect 26186 171098 26422 171334
rect 26186 135418 26422 135654
rect 26186 135098 26422 135334
rect 26186 99418 26422 99654
rect 26186 99098 26422 99334
rect 26186 63418 26422 63654
rect 26186 63098 26422 63334
rect 26186 27418 26422 27654
rect 26186 27098 26422 27334
rect 26186 -5282 26422 -5046
rect 26186 -5602 26422 -5366
rect 47786 710242 48022 710478
rect 47786 709922 48022 710158
rect 44186 708362 44422 708598
rect 44186 708042 44422 708278
rect 40586 706482 40822 706718
rect 40586 706162 40822 706398
rect 29786 679018 30022 679254
rect 29786 678698 30022 678934
rect 29786 643018 30022 643254
rect 29786 642698 30022 642934
rect 29786 607018 30022 607254
rect 29786 606698 30022 606934
rect 29786 571018 30022 571254
rect 29786 570698 30022 570934
rect 29786 535018 30022 535254
rect 29786 534698 30022 534934
rect 29786 499018 30022 499254
rect 29786 498698 30022 498934
rect 29786 463018 30022 463254
rect 29786 462698 30022 462934
rect 29786 427018 30022 427254
rect 29786 426698 30022 426934
rect 29786 391018 30022 391254
rect 29786 390698 30022 390934
rect 29786 355018 30022 355254
rect 29786 354698 30022 354934
rect 29786 319018 30022 319254
rect 29786 318698 30022 318934
rect 29786 283018 30022 283254
rect 29786 282698 30022 282934
rect 29786 247018 30022 247254
rect 29786 246698 30022 246934
rect 29786 211018 30022 211254
rect 29786 210698 30022 210934
rect 29786 175018 30022 175254
rect 29786 174698 30022 174934
rect 29786 139018 30022 139254
rect 29786 138698 30022 138934
rect 29786 103018 30022 103254
rect 29786 102698 30022 102934
rect 29786 67018 30022 67254
rect 29786 66698 30022 66934
rect 29786 31018 30022 31254
rect 29786 30698 30022 30934
rect 11786 -6222 12022 -5986
rect 11786 -6542 12022 -6306
rect -8394 -7162 -8158 -6926
rect -8394 -7482 -8158 -7246
rect 36986 704602 37222 704838
rect 36986 704282 37222 704518
rect 36986 686218 37222 686454
rect 36986 685898 37222 686134
rect 36986 650218 37222 650454
rect 36986 649898 37222 650134
rect 36986 614218 37222 614454
rect 36986 613898 37222 614134
rect 36986 578218 37222 578454
rect 36986 577898 37222 578134
rect 36986 542218 37222 542454
rect 36986 541898 37222 542134
rect 36986 506218 37222 506454
rect 36986 505898 37222 506134
rect 36986 470218 37222 470454
rect 36986 469898 37222 470134
rect 36986 434218 37222 434454
rect 36986 433898 37222 434134
rect 36986 398218 37222 398454
rect 36986 397898 37222 398134
rect 36986 362218 37222 362454
rect 36986 361898 37222 362134
rect 36986 326218 37222 326454
rect 36986 325898 37222 326134
rect 36986 290218 37222 290454
rect 36986 289898 37222 290134
rect 36986 254218 37222 254454
rect 36986 253898 37222 254134
rect 36986 218218 37222 218454
rect 36986 217898 37222 218134
rect 36986 182218 37222 182454
rect 36986 181898 37222 182134
rect 36986 146218 37222 146454
rect 36986 145898 37222 146134
rect 36986 110218 37222 110454
rect 36986 109898 37222 110134
rect 36986 74218 37222 74454
rect 36986 73898 37222 74134
rect 36986 38218 37222 38454
rect 36986 37898 37222 38134
rect 36986 2218 37222 2454
rect 36986 1898 37222 2134
rect 36986 -582 37222 -346
rect 36986 -902 37222 -666
rect 40586 689818 40822 690054
rect 40586 689498 40822 689734
rect 40586 653818 40822 654054
rect 40586 653498 40822 653734
rect 40586 617818 40822 618054
rect 40586 617498 40822 617734
rect 40586 581818 40822 582054
rect 40586 581498 40822 581734
rect 40586 545818 40822 546054
rect 40586 545498 40822 545734
rect 40586 509818 40822 510054
rect 40586 509498 40822 509734
rect 40586 473818 40822 474054
rect 40586 473498 40822 473734
rect 40586 437818 40822 438054
rect 40586 437498 40822 437734
rect 40586 401818 40822 402054
rect 40586 401498 40822 401734
rect 40586 365818 40822 366054
rect 40586 365498 40822 365734
rect 40586 329818 40822 330054
rect 40586 329498 40822 329734
rect 40586 293818 40822 294054
rect 40586 293498 40822 293734
rect 40586 257818 40822 258054
rect 40586 257498 40822 257734
rect 40586 221818 40822 222054
rect 40586 221498 40822 221734
rect 40586 185818 40822 186054
rect 40586 185498 40822 185734
rect 40586 149818 40822 150054
rect 40586 149498 40822 149734
rect 40586 113818 40822 114054
rect 40586 113498 40822 113734
rect 40586 77818 40822 78054
rect 40586 77498 40822 77734
rect 40586 41818 40822 42054
rect 40586 41498 40822 41734
rect 40586 5818 40822 6054
rect 40586 5498 40822 5734
rect 40586 -2462 40822 -2226
rect 40586 -2782 40822 -2546
rect 44186 693418 44422 693654
rect 44186 693098 44422 693334
rect 44186 657418 44422 657654
rect 44186 657098 44422 657334
rect 44186 621418 44422 621654
rect 44186 621098 44422 621334
rect 44186 585418 44422 585654
rect 44186 585098 44422 585334
rect 44186 549418 44422 549654
rect 44186 549098 44422 549334
rect 44186 513418 44422 513654
rect 44186 513098 44422 513334
rect 44186 477418 44422 477654
rect 44186 477098 44422 477334
rect 44186 441418 44422 441654
rect 44186 441098 44422 441334
rect 44186 405418 44422 405654
rect 44186 405098 44422 405334
rect 44186 369418 44422 369654
rect 44186 369098 44422 369334
rect 44186 333418 44422 333654
rect 44186 333098 44422 333334
rect 44186 297418 44422 297654
rect 44186 297098 44422 297334
rect 44186 261418 44422 261654
rect 44186 261098 44422 261334
rect 44186 225418 44422 225654
rect 44186 225098 44422 225334
rect 44186 189418 44422 189654
rect 44186 189098 44422 189334
rect 44186 153418 44422 153654
rect 44186 153098 44422 153334
rect 44186 117418 44422 117654
rect 44186 117098 44422 117334
rect 44186 81418 44422 81654
rect 44186 81098 44422 81334
rect 44186 45418 44422 45654
rect 44186 45098 44422 45334
rect 44186 9418 44422 9654
rect 44186 9098 44422 9334
rect 44186 -4342 44422 -4106
rect 44186 -4662 44422 -4426
rect 65786 711182 66022 711418
rect 65786 710862 66022 711098
rect 62186 709302 62422 709538
rect 62186 708982 62422 709218
rect 58586 707422 58822 707658
rect 58586 707102 58822 707338
rect 47786 697018 48022 697254
rect 47786 696698 48022 696934
rect 47786 661018 48022 661254
rect 47786 660698 48022 660934
rect 47786 625018 48022 625254
rect 47786 624698 48022 624934
rect 47786 589018 48022 589254
rect 47786 588698 48022 588934
rect 47786 553018 48022 553254
rect 47786 552698 48022 552934
rect 47786 517018 48022 517254
rect 47786 516698 48022 516934
rect 47786 481018 48022 481254
rect 47786 480698 48022 480934
rect 47786 445018 48022 445254
rect 47786 444698 48022 444934
rect 47786 409018 48022 409254
rect 47786 408698 48022 408934
rect 47786 373018 48022 373254
rect 47786 372698 48022 372934
rect 47786 337018 48022 337254
rect 47786 336698 48022 336934
rect 47786 301018 48022 301254
rect 47786 300698 48022 300934
rect 47786 265018 48022 265254
rect 47786 264698 48022 264934
rect 47786 229018 48022 229254
rect 47786 228698 48022 228934
rect 47786 193018 48022 193254
rect 47786 192698 48022 192934
rect 47786 157018 48022 157254
rect 47786 156698 48022 156934
rect 47786 121018 48022 121254
rect 47786 120698 48022 120934
rect 47786 85018 48022 85254
rect 47786 84698 48022 84934
rect 47786 49018 48022 49254
rect 47786 48698 48022 48934
rect 47786 13018 48022 13254
rect 47786 12698 48022 12934
rect 29786 -7162 30022 -6926
rect 29786 -7482 30022 -7246
rect 54986 705542 55222 705778
rect 54986 705222 55222 705458
rect 54986 668218 55222 668454
rect 54986 667898 55222 668134
rect 54986 632218 55222 632454
rect 54986 631898 55222 632134
rect 54986 596218 55222 596454
rect 54986 595898 55222 596134
rect 54986 560218 55222 560454
rect 54986 559898 55222 560134
rect 54986 524218 55222 524454
rect 54986 523898 55222 524134
rect 54986 488218 55222 488454
rect 54986 487898 55222 488134
rect 54986 452218 55222 452454
rect 54986 451898 55222 452134
rect 54986 416218 55222 416454
rect 54986 415898 55222 416134
rect 54986 380218 55222 380454
rect 54986 379898 55222 380134
rect 54986 344218 55222 344454
rect 54986 343898 55222 344134
rect 54986 308218 55222 308454
rect 54986 307898 55222 308134
rect 54986 272218 55222 272454
rect 54986 271898 55222 272134
rect 54986 236218 55222 236454
rect 54986 235898 55222 236134
rect 54986 200218 55222 200454
rect 54986 199898 55222 200134
rect 54986 164218 55222 164454
rect 54986 163898 55222 164134
rect 54986 128218 55222 128454
rect 54986 127898 55222 128134
rect 54986 92218 55222 92454
rect 54986 91898 55222 92134
rect 54986 56218 55222 56454
rect 54986 55898 55222 56134
rect 54986 20218 55222 20454
rect 54986 19898 55222 20134
rect 54986 -1522 55222 -1286
rect 54986 -1842 55222 -1606
rect 58586 671818 58822 672054
rect 58586 671498 58822 671734
rect 58586 635818 58822 636054
rect 58586 635498 58822 635734
rect 58586 599818 58822 600054
rect 58586 599498 58822 599734
rect 58586 563818 58822 564054
rect 58586 563498 58822 563734
rect 58586 527818 58822 528054
rect 58586 527498 58822 527734
rect 58586 491818 58822 492054
rect 58586 491498 58822 491734
rect 58586 455818 58822 456054
rect 58586 455498 58822 455734
rect 58586 419818 58822 420054
rect 58586 419498 58822 419734
rect 58586 383818 58822 384054
rect 58586 383498 58822 383734
rect 58586 347818 58822 348054
rect 58586 347498 58822 347734
rect 58586 311818 58822 312054
rect 58586 311498 58822 311734
rect 58586 275818 58822 276054
rect 58586 275498 58822 275734
rect 58586 239818 58822 240054
rect 58586 239498 58822 239734
rect 58586 203818 58822 204054
rect 58586 203498 58822 203734
rect 58586 167818 58822 168054
rect 58586 167498 58822 167734
rect 58586 131818 58822 132054
rect 58586 131498 58822 131734
rect 58586 95818 58822 96054
rect 58586 95498 58822 95734
rect 58586 59818 58822 60054
rect 58586 59498 58822 59734
rect 58586 23818 58822 24054
rect 58586 23498 58822 23734
rect 58586 -3402 58822 -3166
rect 58586 -3722 58822 -3486
rect 62186 675418 62422 675654
rect 62186 675098 62422 675334
rect 62186 639418 62422 639654
rect 62186 639098 62422 639334
rect 62186 603418 62422 603654
rect 62186 603098 62422 603334
rect 62186 567418 62422 567654
rect 62186 567098 62422 567334
rect 62186 531418 62422 531654
rect 62186 531098 62422 531334
rect 62186 495418 62422 495654
rect 62186 495098 62422 495334
rect 62186 459418 62422 459654
rect 62186 459098 62422 459334
rect 62186 423418 62422 423654
rect 62186 423098 62422 423334
rect 62186 387418 62422 387654
rect 62186 387098 62422 387334
rect 62186 351418 62422 351654
rect 62186 351098 62422 351334
rect 62186 315418 62422 315654
rect 62186 315098 62422 315334
rect 62186 279418 62422 279654
rect 62186 279098 62422 279334
rect 62186 243418 62422 243654
rect 62186 243098 62422 243334
rect 62186 207418 62422 207654
rect 62186 207098 62422 207334
rect 62186 171418 62422 171654
rect 62186 171098 62422 171334
rect 62186 135418 62422 135654
rect 62186 135098 62422 135334
rect 62186 99418 62422 99654
rect 62186 99098 62422 99334
rect 62186 63418 62422 63654
rect 62186 63098 62422 63334
rect 62186 27418 62422 27654
rect 62186 27098 62422 27334
rect 62186 -5282 62422 -5046
rect 62186 -5602 62422 -5366
rect 83786 710242 84022 710478
rect 83786 709922 84022 710158
rect 80186 708362 80422 708598
rect 80186 708042 80422 708278
rect 76586 706482 76822 706718
rect 76586 706162 76822 706398
rect 65786 679018 66022 679254
rect 65786 678698 66022 678934
rect 65786 643018 66022 643254
rect 65786 642698 66022 642934
rect 65786 607018 66022 607254
rect 65786 606698 66022 606934
rect 65786 571018 66022 571254
rect 65786 570698 66022 570934
rect 65786 535018 66022 535254
rect 65786 534698 66022 534934
rect 65786 499018 66022 499254
rect 65786 498698 66022 498934
rect 65786 463018 66022 463254
rect 65786 462698 66022 462934
rect 65786 427018 66022 427254
rect 65786 426698 66022 426934
rect 65786 391018 66022 391254
rect 65786 390698 66022 390934
rect 65786 355018 66022 355254
rect 65786 354698 66022 354934
rect 65786 319018 66022 319254
rect 65786 318698 66022 318934
rect 65786 283018 66022 283254
rect 65786 282698 66022 282934
rect 65786 247018 66022 247254
rect 65786 246698 66022 246934
rect 65786 211018 66022 211254
rect 65786 210698 66022 210934
rect 65786 175018 66022 175254
rect 65786 174698 66022 174934
rect 65786 139018 66022 139254
rect 65786 138698 66022 138934
rect 65786 103018 66022 103254
rect 65786 102698 66022 102934
rect 65786 67018 66022 67254
rect 65786 66698 66022 66934
rect 65786 31018 66022 31254
rect 65786 30698 66022 30934
rect 47786 -6222 48022 -5986
rect 47786 -6542 48022 -6306
rect 72986 704602 73222 704838
rect 72986 704282 73222 704518
rect 72986 686218 73222 686454
rect 72986 685898 73222 686134
rect 72986 650218 73222 650454
rect 72986 649898 73222 650134
rect 72986 614218 73222 614454
rect 72986 613898 73222 614134
rect 72986 578218 73222 578454
rect 72986 577898 73222 578134
rect 72986 542218 73222 542454
rect 72986 541898 73222 542134
rect 72986 506218 73222 506454
rect 72986 505898 73222 506134
rect 72986 470218 73222 470454
rect 72986 469898 73222 470134
rect 72986 434218 73222 434454
rect 72986 433898 73222 434134
rect 72986 398218 73222 398454
rect 72986 397898 73222 398134
rect 72986 362218 73222 362454
rect 72986 361898 73222 362134
rect 72986 326218 73222 326454
rect 72986 325898 73222 326134
rect 72986 290218 73222 290454
rect 72986 289898 73222 290134
rect 72986 254218 73222 254454
rect 72986 253898 73222 254134
rect 72986 218218 73222 218454
rect 72986 217898 73222 218134
rect 72986 182218 73222 182454
rect 72986 181898 73222 182134
rect 72986 146218 73222 146454
rect 72986 145898 73222 146134
rect 72986 110218 73222 110454
rect 72986 109898 73222 110134
rect 72986 74218 73222 74454
rect 72986 73898 73222 74134
rect 72986 38218 73222 38454
rect 72986 37898 73222 38134
rect 72986 2218 73222 2454
rect 72986 1898 73222 2134
rect 72986 -582 73222 -346
rect 72986 -902 73222 -666
rect 76586 689818 76822 690054
rect 76586 689498 76822 689734
rect 76586 653818 76822 654054
rect 76586 653498 76822 653734
rect 76586 617818 76822 618054
rect 76586 617498 76822 617734
rect 76586 581818 76822 582054
rect 76586 581498 76822 581734
rect 76586 545818 76822 546054
rect 76586 545498 76822 545734
rect 76586 509818 76822 510054
rect 76586 509498 76822 509734
rect 76586 473818 76822 474054
rect 76586 473498 76822 473734
rect 76586 437818 76822 438054
rect 76586 437498 76822 437734
rect 76586 401818 76822 402054
rect 76586 401498 76822 401734
rect 76586 365818 76822 366054
rect 76586 365498 76822 365734
rect 76586 329818 76822 330054
rect 76586 329498 76822 329734
rect 76586 293818 76822 294054
rect 76586 293498 76822 293734
rect 76586 257818 76822 258054
rect 76586 257498 76822 257734
rect 76586 221818 76822 222054
rect 76586 221498 76822 221734
rect 76586 185818 76822 186054
rect 76586 185498 76822 185734
rect 76586 149818 76822 150054
rect 76586 149498 76822 149734
rect 76586 113818 76822 114054
rect 76586 113498 76822 113734
rect 76586 77818 76822 78054
rect 76586 77498 76822 77734
rect 76586 41818 76822 42054
rect 76586 41498 76822 41734
rect 76586 5818 76822 6054
rect 76586 5498 76822 5734
rect 76586 -2462 76822 -2226
rect 76586 -2782 76822 -2546
rect 80186 693418 80422 693654
rect 80186 693098 80422 693334
rect 80186 657418 80422 657654
rect 80186 657098 80422 657334
rect 80186 621418 80422 621654
rect 80186 621098 80422 621334
rect 80186 585418 80422 585654
rect 80186 585098 80422 585334
rect 80186 549418 80422 549654
rect 80186 549098 80422 549334
rect 80186 513418 80422 513654
rect 80186 513098 80422 513334
rect 80186 477418 80422 477654
rect 80186 477098 80422 477334
rect 80186 441418 80422 441654
rect 80186 441098 80422 441334
rect 80186 405418 80422 405654
rect 80186 405098 80422 405334
rect 80186 369418 80422 369654
rect 80186 369098 80422 369334
rect 80186 333418 80422 333654
rect 80186 333098 80422 333334
rect 80186 297418 80422 297654
rect 80186 297098 80422 297334
rect 80186 261418 80422 261654
rect 80186 261098 80422 261334
rect 80186 225418 80422 225654
rect 80186 225098 80422 225334
rect 80186 189418 80422 189654
rect 80186 189098 80422 189334
rect 80186 153418 80422 153654
rect 80186 153098 80422 153334
rect 80186 117418 80422 117654
rect 80186 117098 80422 117334
rect 80186 81418 80422 81654
rect 80186 81098 80422 81334
rect 80186 45418 80422 45654
rect 80186 45098 80422 45334
rect 80186 9418 80422 9654
rect 80186 9098 80422 9334
rect 80186 -4342 80422 -4106
rect 80186 -4662 80422 -4426
rect 101786 711182 102022 711418
rect 101786 710862 102022 711098
rect 98186 709302 98422 709538
rect 98186 708982 98422 709218
rect 94586 707422 94822 707658
rect 94586 707102 94822 707338
rect 83786 697018 84022 697254
rect 83786 696698 84022 696934
rect 83786 661018 84022 661254
rect 83786 660698 84022 660934
rect 83786 625018 84022 625254
rect 83786 624698 84022 624934
rect 83786 589018 84022 589254
rect 83786 588698 84022 588934
rect 83786 553018 84022 553254
rect 83786 552698 84022 552934
rect 83786 517018 84022 517254
rect 83786 516698 84022 516934
rect 83786 481018 84022 481254
rect 83786 480698 84022 480934
rect 83786 445018 84022 445254
rect 83786 444698 84022 444934
rect 83786 409018 84022 409254
rect 83786 408698 84022 408934
rect 83786 373018 84022 373254
rect 83786 372698 84022 372934
rect 83786 337018 84022 337254
rect 83786 336698 84022 336934
rect 83786 301018 84022 301254
rect 83786 300698 84022 300934
rect 83786 265018 84022 265254
rect 83786 264698 84022 264934
rect 83786 229018 84022 229254
rect 83786 228698 84022 228934
rect 83786 193018 84022 193254
rect 83786 192698 84022 192934
rect 83786 157018 84022 157254
rect 83786 156698 84022 156934
rect 83786 121018 84022 121254
rect 83786 120698 84022 120934
rect 83786 85018 84022 85254
rect 83786 84698 84022 84934
rect 83786 49018 84022 49254
rect 83786 48698 84022 48934
rect 83786 13018 84022 13254
rect 83786 12698 84022 12934
rect 65786 -7162 66022 -6926
rect 65786 -7482 66022 -7246
rect 90986 705542 91222 705778
rect 90986 705222 91222 705458
rect 90986 668218 91222 668454
rect 90986 667898 91222 668134
rect 90986 632218 91222 632454
rect 90986 631898 91222 632134
rect 90986 596218 91222 596454
rect 90986 595898 91222 596134
rect 90986 560218 91222 560454
rect 90986 559898 91222 560134
rect 90986 524218 91222 524454
rect 90986 523898 91222 524134
rect 90986 488218 91222 488454
rect 90986 487898 91222 488134
rect 90986 452218 91222 452454
rect 90986 451898 91222 452134
rect 90986 416218 91222 416454
rect 90986 415898 91222 416134
rect 90986 380218 91222 380454
rect 90986 379898 91222 380134
rect 90986 344218 91222 344454
rect 90986 343898 91222 344134
rect 90986 308218 91222 308454
rect 90986 307898 91222 308134
rect 90986 272218 91222 272454
rect 90986 271898 91222 272134
rect 90986 236218 91222 236454
rect 90986 235898 91222 236134
rect 90986 200218 91222 200454
rect 90986 199898 91222 200134
rect 90986 164218 91222 164454
rect 90986 163898 91222 164134
rect 90986 128218 91222 128454
rect 90986 127898 91222 128134
rect 90986 92218 91222 92454
rect 90986 91898 91222 92134
rect 90986 56218 91222 56454
rect 90986 55898 91222 56134
rect 90986 20218 91222 20454
rect 90986 19898 91222 20134
rect 90986 -1522 91222 -1286
rect 90986 -1842 91222 -1606
rect 94586 671818 94822 672054
rect 94586 671498 94822 671734
rect 94586 635818 94822 636054
rect 94586 635498 94822 635734
rect 94586 599818 94822 600054
rect 94586 599498 94822 599734
rect 94586 563818 94822 564054
rect 94586 563498 94822 563734
rect 94586 527818 94822 528054
rect 94586 527498 94822 527734
rect 94586 491818 94822 492054
rect 94586 491498 94822 491734
rect 94586 455818 94822 456054
rect 94586 455498 94822 455734
rect 94586 419818 94822 420054
rect 94586 419498 94822 419734
rect 94586 383818 94822 384054
rect 94586 383498 94822 383734
rect 94586 347818 94822 348054
rect 94586 347498 94822 347734
rect 94586 311818 94822 312054
rect 94586 311498 94822 311734
rect 94586 275818 94822 276054
rect 94586 275498 94822 275734
rect 94586 239818 94822 240054
rect 94586 239498 94822 239734
rect 94586 203818 94822 204054
rect 94586 203498 94822 203734
rect 94586 167818 94822 168054
rect 94586 167498 94822 167734
rect 94586 131818 94822 132054
rect 94586 131498 94822 131734
rect 94586 95818 94822 96054
rect 94586 95498 94822 95734
rect 94586 59818 94822 60054
rect 94586 59498 94822 59734
rect 94586 23818 94822 24054
rect 94586 23498 94822 23734
rect 94586 -3402 94822 -3166
rect 94586 -3722 94822 -3486
rect 98186 675418 98422 675654
rect 98186 675098 98422 675334
rect 98186 639418 98422 639654
rect 98186 639098 98422 639334
rect 98186 603418 98422 603654
rect 98186 603098 98422 603334
rect 98186 567418 98422 567654
rect 98186 567098 98422 567334
rect 98186 531418 98422 531654
rect 98186 531098 98422 531334
rect 98186 495418 98422 495654
rect 98186 495098 98422 495334
rect 98186 459418 98422 459654
rect 98186 459098 98422 459334
rect 98186 423418 98422 423654
rect 98186 423098 98422 423334
rect 98186 387418 98422 387654
rect 98186 387098 98422 387334
rect 98186 351418 98422 351654
rect 98186 351098 98422 351334
rect 98186 315418 98422 315654
rect 98186 315098 98422 315334
rect 98186 279418 98422 279654
rect 98186 279098 98422 279334
rect 98186 243418 98422 243654
rect 98186 243098 98422 243334
rect 98186 207418 98422 207654
rect 98186 207098 98422 207334
rect 98186 171418 98422 171654
rect 98186 171098 98422 171334
rect 98186 135418 98422 135654
rect 98186 135098 98422 135334
rect 98186 99418 98422 99654
rect 98186 99098 98422 99334
rect 98186 63418 98422 63654
rect 98186 63098 98422 63334
rect 98186 27418 98422 27654
rect 98186 27098 98422 27334
rect 98186 -5282 98422 -5046
rect 98186 -5602 98422 -5366
rect 119786 710242 120022 710478
rect 119786 709922 120022 710158
rect 116186 708362 116422 708598
rect 116186 708042 116422 708278
rect 112586 706482 112822 706718
rect 112586 706162 112822 706398
rect 101786 679018 102022 679254
rect 101786 678698 102022 678934
rect 101786 643018 102022 643254
rect 101786 642698 102022 642934
rect 101786 607018 102022 607254
rect 101786 606698 102022 606934
rect 101786 571018 102022 571254
rect 101786 570698 102022 570934
rect 101786 535018 102022 535254
rect 101786 534698 102022 534934
rect 101786 499018 102022 499254
rect 101786 498698 102022 498934
rect 101786 463018 102022 463254
rect 101786 462698 102022 462934
rect 101786 427018 102022 427254
rect 101786 426698 102022 426934
rect 101786 391018 102022 391254
rect 101786 390698 102022 390934
rect 101786 355018 102022 355254
rect 101786 354698 102022 354934
rect 101786 319018 102022 319254
rect 101786 318698 102022 318934
rect 101786 283018 102022 283254
rect 101786 282698 102022 282934
rect 101786 247018 102022 247254
rect 101786 246698 102022 246934
rect 101786 211018 102022 211254
rect 101786 210698 102022 210934
rect 101786 175018 102022 175254
rect 101786 174698 102022 174934
rect 101786 139018 102022 139254
rect 101786 138698 102022 138934
rect 101786 103018 102022 103254
rect 101786 102698 102022 102934
rect 101786 67018 102022 67254
rect 101786 66698 102022 66934
rect 101786 31018 102022 31254
rect 101786 30698 102022 30934
rect 83786 -6222 84022 -5986
rect 83786 -6542 84022 -6306
rect 108986 704602 109222 704838
rect 108986 704282 109222 704518
rect 108986 686218 109222 686454
rect 108986 685898 109222 686134
rect 108986 650218 109222 650454
rect 108986 649898 109222 650134
rect 108986 614218 109222 614454
rect 108986 613898 109222 614134
rect 108986 578218 109222 578454
rect 108986 577898 109222 578134
rect 108986 542218 109222 542454
rect 108986 541898 109222 542134
rect 108986 506218 109222 506454
rect 108986 505898 109222 506134
rect 108986 470218 109222 470454
rect 108986 469898 109222 470134
rect 108986 434218 109222 434454
rect 108986 433898 109222 434134
rect 108986 398218 109222 398454
rect 108986 397898 109222 398134
rect 108986 362218 109222 362454
rect 108986 361898 109222 362134
rect 108986 326218 109222 326454
rect 108986 325898 109222 326134
rect 108986 290218 109222 290454
rect 108986 289898 109222 290134
rect 108986 254218 109222 254454
rect 108986 253898 109222 254134
rect 108986 218218 109222 218454
rect 108986 217898 109222 218134
rect 108986 182218 109222 182454
rect 108986 181898 109222 182134
rect 108986 146218 109222 146454
rect 108986 145898 109222 146134
rect 108986 110218 109222 110454
rect 108986 109898 109222 110134
rect 108986 74218 109222 74454
rect 108986 73898 109222 74134
rect 108986 38218 109222 38454
rect 108986 37898 109222 38134
rect 108986 2218 109222 2454
rect 108986 1898 109222 2134
rect 108986 -582 109222 -346
rect 108986 -902 109222 -666
rect 112586 689818 112822 690054
rect 112586 689498 112822 689734
rect 112586 653818 112822 654054
rect 112586 653498 112822 653734
rect 112586 617818 112822 618054
rect 112586 617498 112822 617734
rect 112586 581818 112822 582054
rect 112586 581498 112822 581734
rect 112586 545818 112822 546054
rect 112586 545498 112822 545734
rect 112586 509818 112822 510054
rect 112586 509498 112822 509734
rect 112586 473818 112822 474054
rect 112586 473498 112822 473734
rect 112586 437818 112822 438054
rect 112586 437498 112822 437734
rect 112586 401818 112822 402054
rect 112586 401498 112822 401734
rect 112586 365818 112822 366054
rect 112586 365498 112822 365734
rect 112586 329818 112822 330054
rect 112586 329498 112822 329734
rect 112586 293818 112822 294054
rect 112586 293498 112822 293734
rect 112586 257818 112822 258054
rect 112586 257498 112822 257734
rect 112586 221818 112822 222054
rect 112586 221498 112822 221734
rect 112586 185818 112822 186054
rect 112586 185498 112822 185734
rect 112586 149818 112822 150054
rect 112586 149498 112822 149734
rect 112586 113818 112822 114054
rect 112586 113498 112822 113734
rect 112586 77818 112822 78054
rect 112586 77498 112822 77734
rect 112586 41818 112822 42054
rect 112586 41498 112822 41734
rect 112586 5818 112822 6054
rect 112586 5498 112822 5734
rect 112586 -2462 112822 -2226
rect 112586 -2782 112822 -2546
rect 116186 693418 116422 693654
rect 116186 693098 116422 693334
rect 116186 657418 116422 657654
rect 116186 657098 116422 657334
rect 116186 621418 116422 621654
rect 116186 621098 116422 621334
rect 116186 585418 116422 585654
rect 116186 585098 116422 585334
rect 116186 549418 116422 549654
rect 116186 549098 116422 549334
rect 116186 513418 116422 513654
rect 116186 513098 116422 513334
rect 116186 477418 116422 477654
rect 116186 477098 116422 477334
rect 116186 441418 116422 441654
rect 116186 441098 116422 441334
rect 116186 405418 116422 405654
rect 116186 405098 116422 405334
rect 116186 369418 116422 369654
rect 116186 369098 116422 369334
rect 116186 333418 116422 333654
rect 116186 333098 116422 333334
rect 116186 297418 116422 297654
rect 116186 297098 116422 297334
rect 116186 261418 116422 261654
rect 116186 261098 116422 261334
rect 116186 225418 116422 225654
rect 116186 225098 116422 225334
rect 116186 189418 116422 189654
rect 116186 189098 116422 189334
rect 116186 153418 116422 153654
rect 116186 153098 116422 153334
rect 116186 117418 116422 117654
rect 116186 117098 116422 117334
rect 116186 81418 116422 81654
rect 116186 81098 116422 81334
rect 116186 45418 116422 45654
rect 116186 45098 116422 45334
rect 116186 9418 116422 9654
rect 116186 9098 116422 9334
rect 116186 -4342 116422 -4106
rect 116186 -4662 116422 -4426
rect 137786 711182 138022 711418
rect 137786 710862 138022 711098
rect 134186 709302 134422 709538
rect 134186 708982 134422 709218
rect 130586 707422 130822 707658
rect 130586 707102 130822 707338
rect 119786 697018 120022 697254
rect 119786 696698 120022 696934
rect 119786 661018 120022 661254
rect 119786 660698 120022 660934
rect 119786 625018 120022 625254
rect 119786 624698 120022 624934
rect 119786 589018 120022 589254
rect 119786 588698 120022 588934
rect 119786 553018 120022 553254
rect 119786 552698 120022 552934
rect 119786 517018 120022 517254
rect 119786 516698 120022 516934
rect 126986 705542 127222 705778
rect 126986 705222 127222 705458
rect 126986 668218 127222 668454
rect 126986 667898 127222 668134
rect 126986 632218 127222 632454
rect 126986 631898 127222 632134
rect 126986 596218 127222 596454
rect 126986 595898 127222 596134
rect 126986 560218 127222 560454
rect 126986 559898 127222 560134
rect 126986 524218 127222 524454
rect 126986 523898 127222 524134
rect 119786 481018 120022 481254
rect 119786 480698 120022 480934
rect 119786 445018 120022 445254
rect 119786 444698 120022 444934
rect 119786 409018 120022 409254
rect 119786 408698 120022 408934
rect 119786 373018 120022 373254
rect 119786 372698 120022 372934
rect 119786 337018 120022 337254
rect 119786 336698 120022 336934
rect 119786 301018 120022 301254
rect 119786 300698 120022 300934
rect 119786 265018 120022 265254
rect 119786 264698 120022 264934
rect 119786 229018 120022 229254
rect 119786 228698 120022 228934
rect 119786 193018 120022 193254
rect 119786 192698 120022 192934
rect 119786 157018 120022 157254
rect 119786 156698 120022 156934
rect 119786 121018 120022 121254
rect 119786 120698 120022 120934
rect 119786 85018 120022 85254
rect 119786 84698 120022 84934
rect 119786 49018 120022 49254
rect 119786 48698 120022 48934
rect 119786 13018 120022 13254
rect 119786 12698 120022 12934
rect 101786 -7162 102022 -6926
rect 101786 -7482 102022 -7246
rect 126986 488218 127222 488454
rect 126986 487898 127222 488134
rect 126986 452218 127222 452454
rect 126986 451898 127222 452134
rect 126986 416218 127222 416454
rect 126986 415898 127222 416134
rect 126986 380218 127222 380454
rect 126986 379898 127222 380134
rect 126986 344218 127222 344454
rect 126986 343898 127222 344134
rect 126986 308218 127222 308454
rect 126986 307898 127222 308134
rect 126986 272218 127222 272454
rect 126986 271898 127222 272134
rect 126986 236218 127222 236454
rect 126986 235898 127222 236134
rect 126986 200218 127222 200454
rect 126986 199898 127222 200134
rect 126986 164218 127222 164454
rect 126986 163898 127222 164134
rect 126986 128218 127222 128454
rect 126986 127898 127222 128134
rect 126986 92218 127222 92454
rect 126986 91898 127222 92134
rect 126986 56218 127222 56454
rect 126986 55898 127222 56134
rect 126986 20218 127222 20454
rect 126986 19898 127222 20134
rect 126986 -1522 127222 -1286
rect 126986 -1842 127222 -1606
rect 130586 671818 130822 672054
rect 130586 671498 130822 671734
rect 130586 635818 130822 636054
rect 130586 635498 130822 635734
rect 130586 599818 130822 600054
rect 130586 599498 130822 599734
rect 130586 563818 130822 564054
rect 130586 563498 130822 563734
rect 130586 527818 130822 528054
rect 130586 527498 130822 527734
rect 130586 491818 130822 492054
rect 130586 491498 130822 491734
rect 130586 455818 130822 456054
rect 130586 455498 130822 455734
rect 130586 419818 130822 420054
rect 130586 419498 130822 419734
rect 130586 383818 130822 384054
rect 130586 383498 130822 383734
rect 130586 347818 130822 348054
rect 130586 347498 130822 347734
rect 130586 311818 130822 312054
rect 130586 311498 130822 311734
rect 130586 275818 130822 276054
rect 130586 275498 130822 275734
rect 130586 239818 130822 240054
rect 130586 239498 130822 239734
rect 130586 203818 130822 204054
rect 130586 203498 130822 203734
rect 130586 167818 130822 168054
rect 130586 167498 130822 167734
rect 134186 675418 134422 675654
rect 134186 675098 134422 675334
rect 134186 639418 134422 639654
rect 134186 639098 134422 639334
rect 134186 603418 134422 603654
rect 134186 603098 134422 603334
rect 134186 567418 134422 567654
rect 134186 567098 134422 567334
rect 134186 531418 134422 531654
rect 134186 531098 134422 531334
rect 134186 495418 134422 495654
rect 134186 495098 134422 495334
rect 134186 459418 134422 459654
rect 134186 459098 134422 459334
rect 134186 423418 134422 423654
rect 134186 423098 134422 423334
rect 134186 387418 134422 387654
rect 134186 387098 134422 387334
rect 134186 351418 134422 351654
rect 134186 351098 134422 351334
rect 134186 315418 134422 315654
rect 134186 315098 134422 315334
rect 134186 279418 134422 279654
rect 134186 279098 134422 279334
rect 134186 243418 134422 243654
rect 134186 243098 134422 243334
rect 134186 207418 134422 207654
rect 134186 207098 134422 207334
rect 134186 171418 134422 171654
rect 134186 171098 134422 171334
rect 134186 135418 134422 135654
rect 134186 135098 134422 135334
rect 130586 131818 130822 132054
rect 130586 131498 130822 131734
rect 130586 95818 130822 96054
rect 130586 95498 130822 95734
rect 130586 59818 130822 60054
rect 130586 59498 130822 59734
rect 130586 23818 130822 24054
rect 130586 23498 130822 23734
rect 130586 -3402 130822 -3166
rect 130586 -3722 130822 -3486
rect 134186 99418 134422 99654
rect 134186 99098 134422 99334
rect 134186 63418 134422 63654
rect 134186 63098 134422 63334
rect 134186 27418 134422 27654
rect 134186 27098 134422 27334
rect 134186 -5282 134422 -5046
rect 134186 -5602 134422 -5366
rect 155786 710242 156022 710478
rect 155786 709922 156022 710158
rect 152186 708362 152422 708598
rect 152186 708042 152422 708278
rect 148586 706482 148822 706718
rect 148586 706162 148822 706398
rect 137786 679018 138022 679254
rect 137786 678698 138022 678934
rect 137786 643018 138022 643254
rect 137786 642698 138022 642934
rect 137786 607018 138022 607254
rect 137786 606698 138022 606934
rect 137786 571018 138022 571254
rect 137786 570698 138022 570934
rect 137786 535018 138022 535254
rect 137786 534698 138022 534934
rect 137786 499018 138022 499254
rect 137786 498698 138022 498934
rect 137786 463018 138022 463254
rect 137786 462698 138022 462934
rect 137786 427018 138022 427254
rect 137786 426698 138022 426934
rect 137786 391018 138022 391254
rect 137786 390698 138022 390934
rect 137786 355018 138022 355254
rect 137786 354698 138022 354934
rect 137786 319018 138022 319254
rect 137786 318698 138022 318934
rect 137786 283018 138022 283254
rect 137786 282698 138022 282934
rect 137786 247018 138022 247254
rect 137786 246698 138022 246934
rect 137786 211018 138022 211254
rect 137786 210698 138022 210934
rect 137786 175018 138022 175254
rect 137786 174698 138022 174934
rect 137786 139018 138022 139254
rect 137786 138698 138022 138934
rect 137786 103018 138022 103254
rect 137786 102698 138022 102934
rect 137786 67018 138022 67254
rect 137786 66698 138022 66934
rect 137786 31018 138022 31254
rect 137786 30698 138022 30934
rect 119786 -6222 120022 -5986
rect 119786 -6542 120022 -6306
rect 144986 704602 145222 704838
rect 144986 704282 145222 704518
rect 144986 686218 145222 686454
rect 144986 685898 145222 686134
rect 144986 650218 145222 650454
rect 144986 649898 145222 650134
rect 144986 614218 145222 614454
rect 144986 613898 145222 614134
rect 144986 578218 145222 578454
rect 144986 577898 145222 578134
rect 144986 542218 145222 542454
rect 144986 541898 145222 542134
rect 144986 506218 145222 506454
rect 144986 505898 145222 506134
rect 144986 470218 145222 470454
rect 144986 469898 145222 470134
rect 144986 434218 145222 434454
rect 144986 433898 145222 434134
rect 144986 398218 145222 398454
rect 144986 397898 145222 398134
rect 144986 362218 145222 362454
rect 144986 361898 145222 362134
rect 144986 326218 145222 326454
rect 144986 325898 145222 326134
rect 144986 290218 145222 290454
rect 144986 289898 145222 290134
rect 144986 254218 145222 254454
rect 144986 253898 145222 254134
rect 144986 218218 145222 218454
rect 144986 217898 145222 218134
rect 144986 182218 145222 182454
rect 144986 181898 145222 182134
rect 144986 146218 145222 146454
rect 144986 145898 145222 146134
rect 144986 110218 145222 110454
rect 144986 109898 145222 110134
rect 144986 74218 145222 74454
rect 144986 73898 145222 74134
rect 144986 38218 145222 38454
rect 144986 37898 145222 38134
rect 144986 2218 145222 2454
rect 144986 1898 145222 2134
rect 144986 -582 145222 -346
rect 144986 -902 145222 -666
rect 148586 689818 148822 690054
rect 148586 689498 148822 689734
rect 148586 653818 148822 654054
rect 148586 653498 148822 653734
rect 148586 617818 148822 618054
rect 148586 617498 148822 617734
rect 148586 581818 148822 582054
rect 148586 581498 148822 581734
rect 148586 545818 148822 546054
rect 148586 545498 148822 545734
rect 148586 509818 148822 510054
rect 148586 509498 148822 509734
rect 148586 473818 148822 474054
rect 148586 473498 148822 473734
rect 148586 437818 148822 438054
rect 148586 437498 148822 437734
rect 148586 401818 148822 402054
rect 148586 401498 148822 401734
rect 148586 365818 148822 366054
rect 148586 365498 148822 365734
rect 148586 329818 148822 330054
rect 148586 329498 148822 329734
rect 148586 293818 148822 294054
rect 148586 293498 148822 293734
rect 148586 257818 148822 258054
rect 148586 257498 148822 257734
rect 148586 221818 148822 222054
rect 148586 221498 148822 221734
rect 148586 185818 148822 186054
rect 148586 185498 148822 185734
rect 148586 149818 148822 150054
rect 148586 149498 148822 149734
rect 148586 113818 148822 114054
rect 148586 113498 148822 113734
rect 148586 77818 148822 78054
rect 148586 77498 148822 77734
rect 148586 41818 148822 42054
rect 148586 41498 148822 41734
rect 148586 5818 148822 6054
rect 148586 5498 148822 5734
rect 148586 -2462 148822 -2226
rect 148586 -2782 148822 -2546
rect 152186 693418 152422 693654
rect 152186 693098 152422 693334
rect 152186 657418 152422 657654
rect 152186 657098 152422 657334
rect 152186 621418 152422 621654
rect 152186 621098 152422 621334
rect 152186 585418 152422 585654
rect 152186 585098 152422 585334
rect 152186 549418 152422 549654
rect 152186 549098 152422 549334
rect 152186 513418 152422 513654
rect 152186 513098 152422 513334
rect 152186 477418 152422 477654
rect 152186 477098 152422 477334
rect 173786 711182 174022 711418
rect 173786 710862 174022 711098
rect 170186 709302 170422 709538
rect 170186 708982 170422 709218
rect 166586 707422 166822 707658
rect 166586 707102 166822 707338
rect 155786 697018 156022 697254
rect 155786 696698 156022 696934
rect 155786 661018 156022 661254
rect 155786 660698 156022 660934
rect 155786 625018 156022 625254
rect 155786 624698 156022 624934
rect 155786 589018 156022 589254
rect 155786 588698 156022 588934
rect 155786 553018 156022 553254
rect 155786 552698 156022 552934
rect 155786 517018 156022 517254
rect 155786 516698 156022 516934
rect 155786 481018 156022 481254
rect 155786 480698 156022 480934
rect 155786 445018 156022 445254
rect 155786 444698 156022 444934
rect 152186 441418 152422 441654
rect 152186 441098 152422 441334
rect 152186 405418 152422 405654
rect 152186 405098 152422 405334
rect 152186 369418 152422 369654
rect 152186 369098 152422 369334
rect 152186 333418 152422 333654
rect 152186 333098 152422 333334
rect 152186 297418 152422 297654
rect 152186 297098 152422 297334
rect 152186 261418 152422 261654
rect 152186 261098 152422 261334
rect 152186 225418 152422 225654
rect 152186 225098 152422 225334
rect 152186 189418 152422 189654
rect 152186 189098 152422 189334
rect 152186 153418 152422 153654
rect 152186 153098 152422 153334
rect 152186 117418 152422 117654
rect 152186 117098 152422 117334
rect 152186 81418 152422 81654
rect 152186 81098 152422 81334
rect 152186 45418 152422 45654
rect 152186 45098 152422 45334
rect 152186 9418 152422 9654
rect 152186 9098 152422 9334
rect 152186 -4342 152422 -4106
rect 152186 -4662 152422 -4426
rect 155786 409018 156022 409254
rect 155786 408698 156022 408934
rect 155786 373018 156022 373254
rect 155786 372698 156022 372934
rect 155786 337018 156022 337254
rect 155786 336698 156022 336934
rect 155786 301018 156022 301254
rect 155786 300698 156022 300934
rect 155786 265018 156022 265254
rect 155786 264698 156022 264934
rect 155786 229018 156022 229254
rect 155786 228698 156022 228934
rect 155786 193018 156022 193254
rect 155786 192698 156022 192934
rect 155786 157018 156022 157254
rect 155786 156698 156022 156934
rect 155786 121018 156022 121254
rect 155786 120698 156022 120934
rect 155786 85018 156022 85254
rect 155786 84698 156022 84934
rect 155786 49018 156022 49254
rect 155786 48698 156022 48934
rect 155786 13018 156022 13254
rect 155786 12698 156022 12934
rect 137786 -7162 138022 -6926
rect 137786 -7482 138022 -7246
rect 162986 705542 163222 705778
rect 162986 705222 163222 705458
rect 162986 668218 163222 668454
rect 162986 667898 163222 668134
rect 166586 671818 166822 672054
rect 166586 671498 166822 671734
rect 162986 632218 163222 632454
rect 162986 631898 163222 632134
rect 166586 635818 166822 636054
rect 166586 635498 166822 635734
rect 162986 596218 163222 596454
rect 162986 595898 163222 596134
rect 166586 599818 166822 600054
rect 166586 599498 166822 599734
rect 162986 560218 163222 560454
rect 162986 559898 163222 560134
rect 162986 524218 163222 524454
rect 162986 523898 163222 524134
rect 162986 488218 163222 488454
rect 162986 487898 163222 488134
rect 162986 452218 163222 452454
rect 162986 451898 163222 452134
rect 162986 416218 163222 416454
rect 162986 415898 163222 416134
rect 162986 380218 163222 380454
rect 162986 379898 163222 380134
rect 162986 344218 163222 344454
rect 162986 343898 163222 344134
rect 162986 308218 163222 308454
rect 162986 307898 163222 308134
rect 162986 272218 163222 272454
rect 162986 271898 163222 272134
rect 162986 236218 163222 236454
rect 162986 235898 163222 236134
rect 162986 200218 163222 200454
rect 162986 199898 163222 200134
rect 162986 164218 163222 164454
rect 162986 163898 163222 164134
rect 162986 128218 163222 128454
rect 162986 127898 163222 128134
rect 162986 92218 163222 92454
rect 162986 91898 163222 92134
rect 162986 56218 163222 56454
rect 162986 55898 163222 56134
rect 162986 20218 163222 20454
rect 162986 19898 163222 20134
rect 162986 -1522 163222 -1286
rect 162986 -1842 163222 -1606
rect 166586 563818 166822 564054
rect 166586 563498 166822 563734
rect 166586 527818 166822 528054
rect 166586 527498 166822 527734
rect 166586 491818 166822 492054
rect 166586 491498 166822 491734
rect 166586 455818 166822 456054
rect 166586 455498 166822 455734
rect 166586 419818 166822 420054
rect 166586 419498 166822 419734
rect 166586 383818 166822 384054
rect 166586 383498 166822 383734
rect 166586 347818 166822 348054
rect 166586 347498 166822 347734
rect 166586 311818 166822 312054
rect 166586 311498 166822 311734
rect 166586 275818 166822 276054
rect 166586 275498 166822 275734
rect 166586 239818 166822 240054
rect 166586 239498 166822 239734
rect 166586 203818 166822 204054
rect 166586 203498 166822 203734
rect 166586 167818 166822 168054
rect 166586 167498 166822 167734
rect 166586 131818 166822 132054
rect 166586 131498 166822 131734
rect 166586 95818 166822 96054
rect 166586 95498 166822 95734
rect 166586 59818 166822 60054
rect 166586 59498 166822 59734
rect 166586 23818 166822 24054
rect 166586 23498 166822 23734
rect 166586 -3402 166822 -3166
rect 166586 -3722 166822 -3486
rect 170186 675418 170422 675654
rect 170186 675098 170422 675334
rect 170186 639418 170422 639654
rect 170186 639098 170422 639334
rect 170186 603418 170422 603654
rect 170186 603098 170422 603334
rect 170186 567418 170422 567654
rect 170186 567098 170422 567334
rect 170186 531418 170422 531654
rect 170186 531098 170422 531334
rect 170186 495418 170422 495654
rect 170186 495098 170422 495334
rect 170186 459418 170422 459654
rect 170186 459098 170422 459334
rect 170186 423418 170422 423654
rect 170186 423098 170422 423334
rect 170186 387418 170422 387654
rect 170186 387098 170422 387334
rect 170186 351418 170422 351654
rect 170186 351098 170422 351334
rect 170186 315418 170422 315654
rect 170186 315098 170422 315334
rect 170186 279418 170422 279654
rect 170186 279098 170422 279334
rect 170186 243418 170422 243654
rect 170186 243098 170422 243334
rect 170186 207418 170422 207654
rect 170186 207098 170422 207334
rect 170186 171418 170422 171654
rect 170186 171098 170422 171334
rect 170186 135418 170422 135654
rect 170186 135098 170422 135334
rect 170186 99418 170422 99654
rect 170186 99098 170422 99334
rect 170186 63418 170422 63654
rect 170186 63098 170422 63334
rect 170186 27418 170422 27654
rect 170186 27098 170422 27334
rect 170186 -5282 170422 -5046
rect 170186 -5602 170422 -5366
rect 191786 710242 192022 710478
rect 191786 709922 192022 710158
rect 188186 708362 188422 708598
rect 188186 708042 188422 708278
rect 184586 706482 184822 706718
rect 184586 706162 184822 706398
rect 173786 679018 174022 679254
rect 173786 678698 174022 678934
rect 173786 643018 174022 643254
rect 173786 642698 174022 642934
rect 173786 607018 174022 607254
rect 173786 606698 174022 606934
rect 173786 571018 174022 571254
rect 173786 570698 174022 570934
rect 173786 535018 174022 535254
rect 173786 534698 174022 534934
rect 173786 499018 174022 499254
rect 173786 498698 174022 498934
rect 173786 463018 174022 463254
rect 173786 462698 174022 462934
rect 173786 427018 174022 427254
rect 173786 426698 174022 426934
rect 173786 391018 174022 391254
rect 173786 390698 174022 390934
rect 173786 355018 174022 355254
rect 173786 354698 174022 354934
rect 173786 319018 174022 319254
rect 173786 318698 174022 318934
rect 173786 283018 174022 283254
rect 173786 282698 174022 282934
rect 173786 247018 174022 247254
rect 173786 246698 174022 246934
rect 173786 211018 174022 211254
rect 173786 210698 174022 210934
rect 173786 175018 174022 175254
rect 173786 174698 174022 174934
rect 173786 139018 174022 139254
rect 173786 138698 174022 138934
rect 173786 103018 174022 103254
rect 173786 102698 174022 102934
rect 173786 67018 174022 67254
rect 173786 66698 174022 66934
rect 173786 31018 174022 31254
rect 173786 30698 174022 30934
rect 155786 -6222 156022 -5986
rect 155786 -6542 156022 -6306
rect 180986 704602 181222 704838
rect 180986 704282 181222 704518
rect 180986 686218 181222 686454
rect 180986 685898 181222 686134
rect 180986 650218 181222 650454
rect 180986 649898 181222 650134
rect 180986 614218 181222 614454
rect 180986 613898 181222 614134
rect 180986 578218 181222 578454
rect 180986 577898 181222 578134
rect 180986 542218 181222 542454
rect 180986 541898 181222 542134
rect 180986 506218 181222 506454
rect 180986 505898 181222 506134
rect 180986 470218 181222 470454
rect 180986 469898 181222 470134
rect 180986 434218 181222 434454
rect 180986 433898 181222 434134
rect 180986 398218 181222 398454
rect 180986 397898 181222 398134
rect 180986 362218 181222 362454
rect 180986 361898 181222 362134
rect 180986 326218 181222 326454
rect 180986 325898 181222 326134
rect 180986 290218 181222 290454
rect 180986 289898 181222 290134
rect 180986 254218 181222 254454
rect 180986 253898 181222 254134
rect 180986 218218 181222 218454
rect 180986 217898 181222 218134
rect 180986 182218 181222 182454
rect 180986 181898 181222 182134
rect 180986 146218 181222 146454
rect 180986 145898 181222 146134
rect 180986 110218 181222 110454
rect 180986 109898 181222 110134
rect 180986 74218 181222 74454
rect 180986 73898 181222 74134
rect 184586 689818 184822 690054
rect 184586 689498 184822 689734
rect 184586 653818 184822 654054
rect 184586 653498 184822 653734
rect 184586 617818 184822 618054
rect 184586 617498 184822 617734
rect 184586 581818 184822 582054
rect 184586 581498 184822 581734
rect 184586 545818 184822 546054
rect 184586 545498 184822 545734
rect 184586 509818 184822 510054
rect 184586 509498 184822 509734
rect 184586 473818 184822 474054
rect 184586 473498 184822 473734
rect 184586 437818 184822 438054
rect 184586 437498 184822 437734
rect 184586 401818 184822 402054
rect 184586 401498 184822 401734
rect 184586 365818 184822 366054
rect 184586 365498 184822 365734
rect 184586 329818 184822 330054
rect 184586 329498 184822 329734
rect 184586 293818 184822 294054
rect 184586 293498 184822 293734
rect 184586 257818 184822 258054
rect 184586 257498 184822 257734
rect 184586 221818 184822 222054
rect 184586 221498 184822 221734
rect 184586 185818 184822 186054
rect 184586 185498 184822 185734
rect 184586 149818 184822 150054
rect 184586 149498 184822 149734
rect 184586 113818 184822 114054
rect 184586 113498 184822 113734
rect 184586 77818 184822 78054
rect 184586 77498 184822 77734
rect 184586 41818 184822 42054
rect 184586 41498 184822 41734
rect 180986 38218 181222 38454
rect 180986 37898 181222 38134
rect 180986 2218 181222 2454
rect 180986 1898 181222 2134
rect 180986 -582 181222 -346
rect 180986 -902 181222 -666
rect 184586 5818 184822 6054
rect 184586 5498 184822 5734
rect 184586 -2462 184822 -2226
rect 184586 -2782 184822 -2546
rect 188186 693418 188422 693654
rect 188186 693098 188422 693334
rect 188186 657418 188422 657654
rect 188186 657098 188422 657334
rect 188186 621418 188422 621654
rect 188186 621098 188422 621334
rect 188186 585418 188422 585654
rect 188186 585098 188422 585334
rect 188186 549418 188422 549654
rect 188186 549098 188422 549334
rect 188186 513418 188422 513654
rect 188186 513098 188422 513334
rect 188186 477418 188422 477654
rect 188186 477098 188422 477334
rect 188186 441418 188422 441654
rect 188186 441098 188422 441334
rect 188186 405418 188422 405654
rect 188186 405098 188422 405334
rect 188186 369418 188422 369654
rect 188186 369098 188422 369334
rect 188186 333418 188422 333654
rect 188186 333098 188422 333334
rect 188186 297418 188422 297654
rect 188186 297098 188422 297334
rect 188186 261418 188422 261654
rect 188186 261098 188422 261334
rect 188186 225418 188422 225654
rect 188186 225098 188422 225334
rect 188186 189418 188422 189654
rect 188186 189098 188422 189334
rect 188186 153418 188422 153654
rect 188186 153098 188422 153334
rect 188186 117418 188422 117654
rect 188186 117098 188422 117334
rect 188186 81418 188422 81654
rect 188186 81098 188422 81334
rect 188186 45418 188422 45654
rect 188186 45098 188422 45334
rect 188186 9418 188422 9654
rect 188186 9098 188422 9334
rect 188186 -4342 188422 -4106
rect 188186 -4662 188422 -4426
rect 209786 711182 210022 711418
rect 209786 710862 210022 711098
rect 206186 709302 206422 709538
rect 206186 708982 206422 709218
rect 202586 707422 202822 707658
rect 202586 707102 202822 707338
rect 191786 697018 192022 697254
rect 191786 696698 192022 696934
rect 191786 661018 192022 661254
rect 191786 660698 192022 660934
rect 191786 625018 192022 625254
rect 191786 624698 192022 624934
rect 191786 589018 192022 589254
rect 191786 588698 192022 588934
rect 198986 705542 199222 705778
rect 198986 705222 199222 705458
rect 198986 668218 199222 668454
rect 198986 667898 199222 668134
rect 198986 632218 199222 632454
rect 198986 631898 199222 632134
rect 198986 596218 199222 596454
rect 198986 595898 199222 596134
rect 202586 671818 202822 672054
rect 202586 671498 202822 671734
rect 202586 635818 202822 636054
rect 202586 635498 202822 635734
rect 202586 599818 202822 600054
rect 202586 599498 202822 599734
rect 202586 563818 202822 564054
rect 202586 563498 202822 563734
rect 198986 560218 199222 560454
rect 198986 559898 199222 560134
rect 191786 553018 192022 553254
rect 191786 552698 192022 552934
rect 191786 517018 192022 517254
rect 191786 516698 192022 516934
rect 191786 481018 192022 481254
rect 191786 480698 192022 480934
rect 191786 445018 192022 445254
rect 191786 444698 192022 444934
rect 191786 409018 192022 409254
rect 191786 408698 192022 408934
rect 191786 373018 192022 373254
rect 191786 372698 192022 372934
rect 191786 337018 192022 337254
rect 191786 336698 192022 336934
rect 191786 301018 192022 301254
rect 191786 300698 192022 300934
rect 191786 265018 192022 265254
rect 191786 264698 192022 264934
rect 191786 229018 192022 229254
rect 191786 228698 192022 228934
rect 198986 524218 199222 524454
rect 198986 523898 199222 524134
rect 198986 488218 199222 488454
rect 198986 487898 199222 488134
rect 198986 452218 199222 452454
rect 198986 451898 199222 452134
rect 198986 416218 199222 416454
rect 198986 415898 199222 416134
rect 198986 380218 199222 380454
rect 198986 379898 199222 380134
rect 198986 344218 199222 344454
rect 198986 343898 199222 344134
rect 198986 308218 199222 308454
rect 198986 307898 199222 308134
rect 198986 272218 199222 272454
rect 198986 271898 199222 272134
rect 198986 236218 199222 236454
rect 198986 235898 199222 236134
rect 191786 193018 192022 193254
rect 191786 192698 192022 192934
rect 191786 157018 192022 157254
rect 191786 156698 192022 156934
rect 191786 121018 192022 121254
rect 191786 120698 192022 120934
rect 191786 85018 192022 85254
rect 191786 84698 192022 84934
rect 191786 49018 192022 49254
rect 191786 48698 192022 48934
rect 191786 13018 192022 13254
rect 191786 12698 192022 12934
rect 173786 -7162 174022 -6926
rect 173786 -7482 174022 -7246
rect 202586 527818 202822 528054
rect 202586 527498 202822 527734
rect 202586 491818 202822 492054
rect 202586 491498 202822 491734
rect 202586 455818 202822 456054
rect 202586 455498 202822 455734
rect 202586 419818 202822 420054
rect 202586 419498 202822 419734
rect 202586 383818 202822 384054
rect 202586 383498 202822 383734
rect 202586 347818 202822 348054
rect 202586 347498 202822 347734
rect 202586 311818 202822 312054
rect 202586 311498 202822 311734
rect 202586 275818 202822 276054
rect 202586 275498 202822 275734
rect 202586 239818 202822 240054
rect 202586 239498 202822 239734
rect 202586 203818 202822 204054
rect 202586 203498 202822 203734
rect 198986 200218 199222 200454
rect 198986 199898 199222 200134
rect 198986 164218 199222 164454
rect 198986 163898 199222 164134
rect 198986 128218 199222 128454
rect 198986 127898 199222 128134
rect 198986 92218 199222 92454
rect 198986 91898 199222 92134
rect 198986 56218 199222 56454
rect 198986 55898 199222 56134
rect 198986 20218 199222 20454
rect 198986 19898 199222 20134
rect 198986 -1522 199222 -1286
rect 198986 -1842 199222 -1606
rect 202586 167818 202822 168054
rect 202586 167498 202822 167734
rect 202586 131818 202822 132054
rect 202586 131498 202822 131734
rect 202586 95818 202822 96054
rect 202586 95498 202822 95734
rect 202586 59818 202822 60054
rect 202586 59498 202822 59734
rect 202586 23818 202822 24054
rect 202586 23498 202822 23734
rect 202586 -3402 202822 -3166
rect 202586 -3722 202822 -3486
rect 206186 675418 206422 675654
rect 206186 675098 206422 675334
rect 206186 639418 206422 639654
rect 206186 639098 206422 639334
rect 206186 603418 206422 603654
rect 206186 603098 206422 603334
rect 206186 567418 206422 567654
rect 206186 567098 206422 567334
rect 206186 531418 206422 531654
rect 206186 531098 206422 531334
rect 206186 495418 206422 495654
rect 206186 495098 206422 495334
rect 206186 459418 206422 459654
rect 206186 459098 206422 459334
rect 206186 423418 206422 423654
rect 206186 423098 206422 423334
rect 206186 387418 206422 387654
rect 206186 387098 206422 387334
rect 206186 351418 206422 351654
rect 206186 351098 206422 351334
rect 206186 315418 206422 315654
rect 206186 315098 206422 315334
rect 206186 279418 206422 279654
rect 206186 279098 206422 279334
rect 206186 243418 206422 243654
rect 206186 243098 206422 243334
rect 206186 207418 206422 207654
rect 206186 207098 206422 207334
rect 206186 171418 206422 171654
rect 206186 171098 206422 171334
rect 206186 135418 206422 135654
rect 206186 135098 206422 135334
rect 206186 99418 206422 99654
rect 206186 99098 206422 99334
rect 206186 63418 206422 63654
rect 206186 63098 206422 63334
rect 206186 27418 206422 27654
rect 206186 27098 206422 27334
rect 206186 -5282 206422 -5046
rect 206186 -5602 206422 -5366
rect 227786 710242 228022 710478
rect 227786 709922 228022 710158
rect 224186 708362 224422 708598
rect 224186 708042 224422 708278
rect 220586 706482 220822 706718
rect 220586 706162 220822 706398
rect 209786 679018 210022 679254
rect 209786 678698 210022 678934
rect 209786 643018 210022 643254
rect 209786 642698 210022 642934
rect 209786 607018 210022 607254
rect 209786 606698 210022 606934
rect 209786 571018 210022 571254
rect 209786 570698 210022 570934
rect 209786 535018 210022 535254
rect 209786 534698 210022 534934
rect 209786 499018 210022 499254
rect 209786 498698 210022 498934
rect 209786 463018 210022 463254
rect 209786 462698 210022 462934
rect 209786 427018 210022 427254
rect 209786 426698 210022 426934
rect 209786 391018 210022 391254
rect 209786 390698 210022 390934
rect 209786 355018 210022 355254
rect 209786 354698 210022 354934
rect 209786 319018 210022 319254
rect 209786 318698 210022 318934
rect 209786 283018 210022 283254
rect 209786 282698 210022 282934
rect 209786 247018 210022 247254
rect 209786 246698 210022 246934
rect 209786 211018 210022 211254
rect 209786 210698 210022 210934
rect 209786 175018 210022 175254
rect 209786 174698 210022 174934
rect 209786 139018 210022 139254
rect 209786 138698 210022 138934
rect 209786 103018 210022 103254
rect 209786 102698 210022 102934
rect 209786 67018 210022 67254
rect 209786 66698 210022 66934
rect 209786 31018 210022 31254
rect 209786 30698 210022 30934
rect 191786 -6222 192022 -5986
rect 191786 -6542 192022 -6306
rect 216986 704602 217222 704838
rect 216986 704282 217222 704518
rect 216986 686218 217222 686454
rect 216986 685898 217222 686134
rect 216986 650218 217222 650454
rect 216986 649898 217222 650134
rect 216986 614218 217222 614454
rect 216986 613898 217222 614134
rect 216986 578218 217222 578454
rect 216986 577898 217222 578134
rect 216986 542218 217222 542454
rect 216986 541898 217222 542134
rect 216986 506218 217222 506454
rect 216986 505898 217222 506134
rect 216986 470218 217222 470454
rect 216986 469898 217222 470134
rect 216986 434218 217222 434454
rect 216986 433898 217222 434134
rect 216986 398218 217222 398454
rect 216986 397898 217222 398134
rect 216986 362218 217222 362454
rect 216986 361898 217222 362134
rect 216986 326218 217222 326454
rect 216986 325898 217222 326134
rect 216986 290218 217222 290454
rect 216986 289898 217222 290134
rect 216986 254218 217222 254454
rect 216986 253898 217222 254134
rect 216986 218218 217222 218454
rect 216986 217898 217222 218134
rect 216986 182218 217222 182454
rect 216986 181898 217222 182134
rect 216986 146218 217222 146454
rect 216986 145898 217222 146134
rect 216986 110218 217222 110454
rect 216986 109898 217222 110134
rect 216986 74218 217222 74454
rect 216986 73898 217222 74134
rect 216986 38218 217222 38454
rect 216986 37898 217222 38134
rect 216986 2218 217222 2454
rect 216986 1898 217222 2134
rect 216986 -582 217222 -346
rect 216986 -902 217222 -666
rect 220586 689818 220822 690054
rect 220586 689498 220822 689734
rect 220586 653818 220822 654054
rect 220586 653498 220822 653734
rect 220586 617818 220822 618054
rect 220586 617498 220822 617734
rect 220586 581818 220822 582054
rect 220586 581498 220822 581734
rect 220586 545818 220822 546054
rect 220586 545498 220822 545734
rect 220586 509818 220822 510054
rect 220586 509498 220822 509734
rect 220586 473818 220822 474054
rect 220586 473498 220822 473734
rect 220586 437818 220822 438054
rect 220586 437498 220822 437734
rect 220586 401818 220822 402054
rect 220586 401498 220822 401734
rect 220586 365818 220822 366054
rect 220586 365498 220822 365734
rect 220586 329818 220822 330054
rect 220586 329498 220822 329734
rect 220586 293818 220822 294054
rect 220586 293498 220822 293734
rect 220586 257818 220822 258054
rect 220586 257498 220822 257734
rect 220586 221818 220822 222054
rect 220586 221498 220822 221734
rect 220586 185818 220822 186054
rect 220586 185498 220822 185734
rect 220586 149818 220822 150054
rect 220586 149498 220822 149734
rect 220586 113818 220822 114054
rect 220586 113498 220822 113734
rect 220586 77818 220822 78054
rect 220586 77498 220822 77734
rect 220586 41818 220822 42054
rect 220586 41498 220822 41734
rect 220586 5818 220822 6054
rect 220586 5498 220822 5734
rect 220586 -2462 220822 -2226
rect 220586 -2782 220822 -2546
rect 224186 693418 224422 693654
rect 224186 693098 224422 693334
rect 224186 657418 224422 657654
rect 224186 657098 224422 657334
rect 224186 621418 224422 621654
rect 224186 621098 224422 621334
rect 224186 585418 224422 585654
rect 224186 585098 224422 585334
rect 224186 549418 224422 549654
rect 224186 549098 224422 549334
rect 224186 513418 224422 513654
rect 224186 513098 224422 513334
rect 224186 477418 224422 477654
rect 224186 477098 224422 477334
rect 224186 441418 224422 441654
rect 224186 441098 224422 441334
rect 224186 405418 224422 405654
rect 224186 405098 224422 405334
rect 224186 369418 224422 369654
rect 224186 369098 224422 369334
rect 224186 333418 224422 333654
rect 224186 333098 224422 333334
rect 224186 297418 224422 297654
rect 224186 297098 224422 297334
rect 224186 261418 224422 261654
rect 224186 261098 224422 261334
rect 224186 225418 224422 225654
rect 224186 225098 224422 225334
rect 224186 189418 224422 189654
rect 224186 189098 224422 189334
rect 224186 153418 224422 153654
rect 224186 153098 224422 153334
rect 224186 117418 224422 117654
rect 224186 117098 224422 117334
rect 224186 81418 224422 81654
rect 224186 81098 224422 81334
rect 224186 45418 224422 45654
rect 224186 45098 224422 45334
rect 224186 9418 224422 9654
rect 224186 9098 224422 9334
rect 224186 -4342 224422 -4106
rect 224186 -4662 224422 -4426
rect 245786 711182 246022 711418
rect 245786 710862 246022 711098
rect 242186 709302 242422 709538
rect 242186 708982 242422 709218
rect 238586 707422 238822 707658
rect 238586 707102 238822 707338
rect 227786 697018 228022 697254
rect 227786 696698 228022 696934
rect 227786 661018 228022 661254
rect 227786 660698 228022 660934
rect 227786 625018 228022 625254
rect 227786 624698 228022 624934
rect 227786 589018 228022 589254
rect 227786 588698 228022 588934
rect 227786 553018 228022 553254
rect 227786 552698 228022 552934
rect 227786 517018 228022 517254
rect 227786 516698 228022 516934
rect 227786 481018 228022 481254
rect 227786 480698 228022 480934
rect 227786 445018 228022 445254
rect 227786 444698 228022 444934
rect 227786 409018 228022 409254
rect 227786 408698 228022 408934
rect 227786 373018 228022 373254
rect 227786 372698 228022 372934
rect 227786 337018 228022 337254
rect 227786 336698 228022 336934
rect 227786 301018 228022 301254
rect 227786 300698 228022 300934
rect 227786 265018 228022 265254
rect 227786 264698 228022 264934
rect 227786 229018 228022 229254
rect 227786 228698 228022 228934
rect 227786 193018 228022 193254
rect 227786 192698 228022 192934
rect 227786 157018 228022 157254
rect 227786 156698 228022 156934
rect 227786 121018 228022 121254
rect 227786 120698 228022 120934
rect 227786 85018 228022 85254
rect 227786 84698 228022 84934
rect 227786 49018 228022 49254
rect 227786 48698 228022 48934
rect 227786 13018 228022 13254
rect 227786 12698 228022 12934
rect 209786 -7162 210022 -6926
rect 209786 -7482 210022 -7246
rect 234986 705542 235222 705778
rect 234986 705222 235222 705458
rect 234986 668218 235222 668454
rect 234986 667898 235222 668134
rect 234986 632218 235222 632454
rect 234986 631898 235222 632134
rect 234986 596218 235222 596454
rect 234986 595898 235222 596134
rect 234986 560218 235222 560454
rect 234986 559898 235222 560134
rect 234986 524218 235222 524454
rect 234986 523898 235222 524134
rect 234986 488218 235222 488454
rect 234986 487898 235222 488134
rect 234986 452218 235222 452454
rect 234986 451898 235222 452134
rect 234986 416218 235222 416454
rect 234986 415898 235222 416134
rect 234986 380218 235222 380454
rect 234986 379898 235222 380134
rect 234986 344218 235222 344454
rect 234986 343898 235222 344134
rect 234986 308218 235222 308454
rect 234986 307898 235222 308134
rect 234986 272218 235222 272454
rect 234986 271898 235222 272134
rect 234986 236218 235222 236454
rect 234986 235898 235222 236134
rect 234986 200218 235222 200454
rect 234986 199898 235222 200134
rect 234986 164218 235222 164454
rect 234986 163898 235222 164134
rect 234986 128218 235222 128454
rect 234986 127898 235222 128134
rect 234986 92218 235222 92454
rect 234986 91898 235222 92134
rect 234986 56218 235222 56454
rect 234986 55898 235222 56134
rect 234986 20218 235222 20454
rect 234986 19898 235222 20134
rect 234986 -1522 235222 -1286
rect 234986 -1842 235222 -1606
rect 238586 671818 238822 672054
rect 238586 671498 238822 671734
rect 238586 635818 238822 636054
rect 238586 635498 238822 635734
rect 238586 599818 238822 600054
rect 238586 599498 238822 599734
rect 238586 563818 238822 564054
rect 238586 563498 238822 563734
rect 238586 527818 238822 528054
rect 238586 527498 238822 527734
rect 238586 491818 238822 492054
rect 238586 491498 238822 491734
rect 238586 455818 238822 456054
rect 238586 455498 238822 455734
rect 238586 419818 238822 420054
rect 238586 419498 238822 419734
rect 238586 383818 238822 384054
rect 238586 383498 238822 383734
rect 238586 347818 238822 348054
rect 238586 347498 238822 347734
rect 238586 311818 238822 312054
rect 238586 311498 238822 311734
rect 238586 275818 238822 276054
rect 238586 275498 238822 275734
rect 238586 239818 238822 240054
rect 238586 239498 238822 239734
rect 238586 203818 238822 204054
rect 238586 203498 238822 203734
rect 238586 167818 238822 168054
rect 238586 167498 238822 167734
rect 238586 131818 238822 132054
rect 238586 131498 238822 131734
rect 238586 95818 238822 96054
rect 238586 95498 238822 95734
rect 238586 59818 238822 60054
rect 238586 59498 238822 59734
rect 238586 23818 238822 24054
rect 238586 23498 238822 23734
rect 238586 -3402 238822 -3166
rect 238586 -3722 238822 -3486
rect 242186 675418 242422 675654
rect 242186 675098 242422 675334
rect 242186 639418 242422 639654
rect 242186 639098 242422 639334
rect 242186 603418 242422 603654
rect 242186 603098 242422 603334
rect 242186 567418 242422 567654
rect 242186 567098 242422 567334
rect 242186 531418 242422 531654
rect 242186 531098 242422 531334
rect 242186 495418 242422 495654
rect 242186 495098 242422 495334
rect 242186 459418 242422 459654
rect 242186 459098 242422 459334
rect 242186 423418 242422 423654
rect 242186 423098 242422 423334
rect 242186 387418 242422 387654
rect 242186 387098 242422 387334
rect 242186 351418 242422 351654
rect 242186 351098 242422 351334
rect 242186 315418 242422 315654
rect 242186 315098 242422 315334
rect 242186 279418 242422 279654
rect 242186 279098 242422 279334
rect 242186 243418 242422 243654
rect 242186 243098 242422 243334
rect 242186 207418 242422 207654
rect 242186 207098 242422 207334
rect 242186 171418 242422 171654
rect 242186 171098 242422 171334
rect 242186 135418 242422 135654
rect 242186 135098 242422 135334
rect 242186 99418 242422 99654
rect 242186 99098 242422 99334
rect 242186 63418 242422 63654
rect 242186 63098 242422 63334
rect 242186 27418 242422 27654
rect 242186 27098 242422 27334
rect 242186 -5282 242422 -5046
rect 242186 -5602 242422 -5366
rect 263786 710242 264022 710478
rect 263786 709922 264022 710158
rect 260186 708362 260422 708598
rect 260186 708042 260422 708278
rect 256586 706482 256822 706718
rect 256586 706162 256822 706398
rect 245786 679018 246022 679254
rect 245786 678698 246022 678934
rect 245786 643018 246022 643254
rect 245786 642698 246022 642934
rect 245786 607018 246022 607254
rect 245786 606698 246022 606934
rect 245786 571018 246022 571254
rect 245786 570698 246022 570934
rect 245786 535018 246022 535254
rect 245786 534698 246022 534934
rect 245786 499018 246022 499254
rect 245786 498698 246022 498934
rect 245786 463018 246022 463254
rect 245786 462698 246022 462934
rect 245786 427018 246022 427254
rect 245786 426698 246022 426934
rect 245786 391018 246022 391254
rect 245786 390698 246022 390934
rect 245786 355018 246022 355254
rect 245786 354698 246022 354934
rect 245786 319018 246022 319254
rect 245786 318698 246022 318934
rect 245786 283018 246022 283254
rect 245786 282698 246022 282934
rect 245786 247018 246022 247254
rect 245786 246698 246022 246934
rect 245786 211018 246022 211254
rect 245786 210698 246022 210934
rect 245786 175018 246022 175254
rect 245786 174698 246022 174934
rect 245786 139018 246022 139254
rect 245786 138698 246022 138934
rect 245786 103018 246022 103254
rect 245786 102698 246022 102934
rect 245786 67018 246022 67254
rect 245786 66698 246022 66934
rect 245786 31018 246022 31254
rect 245786 30698 246022 30934
rect 227786 -6222 228022 -5986
rect 227786 -6542 228022 -6306
rect 252986 704602 253222 704838
rect 252986 704282 253222 704518
rect 252986 686218 253222 686454
rect 252986 685898 253222 686134
rect 252986 650218 253222 650454
rect 252986 649898 253222 650134
rect 252986 614218 253222 614454
rect 252986 613898 253222 614134
rect 252986 578218 253222 578454
rect 252986 577898 253222 578134
rect 252986 542218 253222 542454
rect 252986 541898 253222 542134
rect 252986 506218 253222 506454
rect 252986 505898 253222 506134
rect 252986 470218 253222 470454
rect 252986 469898 253222 470134
rect 252986 434218 253222 434454
rect 252986 433898 253222 434134
rect 252986 398218 253222 398454
rect 252986 397898 253222 398134
rect 252986 362218 253222 362454
rect 252986 361898 253222 362134
rect 252986 326218 253222 326454
rect 252986 325898 253222 326134
rect 252986 290218 253222 290454
rect 252986 289898 253222 290134
rect 252986 254218 253222 254454
rect 252986 253898 253222 254134
rect 252986 218218 253222 218454
rect 252986 217898 253222 218134
rect 252986 182218 253222 182454
rect 252986 181898 253222 182134
rect 252986 146218 253222 146454
rect 252986 145898 253222 146134
rect 252986 110218 253222 110454
rect 252986 109898 253222 110134
rect 252986 74218 253222 74454
rect 252986 73898 253222 74134
rect 252986 38218 253222 38454
rect 252986 37898 253222 38134
rect 252986 2218 253222 2454
rect 252986 1898 253222 2134
rect 252986 -582 253222 -346
rect 252986 -902 253222 -666
rect 256586 689818 256822 690054
rect 256586 689498 256822 689734
rect 256586 653818 256822 654054
rect 256586 653498 256822 653734
rect 256586 617818 256822 618054
rect 256586 617498 256822 617734
rect 256586 581818 256822 582054
rect 256586 581498 256822 581734
rect 256586 545818 256822 546054
rect 256586 545498 256822 545734
rect 256586 509818 256822 510054
rect 256586 509498 256822 509734
rect 256586 473818 256822 474054
rect 256586 473498 256822 473734
rect 256586 437818 256822 438054
rect 256586 437498 256822 437734
rect 256586 401818 256822 402054
rect 256586 401498 256822 401734
rect 256586 365818 256822 366054
rect 256586 365498 256822 365734
rect 256586 329818 256822 330054
rect 256586 329498 256822 329734
rect 260186 693418 260422 693654
rect 260186 693098 260422 693334
rect 260186 657418 260422 657654
rect 260186 657098 260422 657334
rect 260186 621418 260422 621654
rect 260186 621098 260422 621334
rect 260186 585418 260422 585654
rect 260186 585098 260422 585334
rect 260186 549418 260422 549654
rect 260186 549098 260422 549334
rect 260186 513418 260422 513654
rect 260186 513098 260422 513334
rect 260186 477418 260422 477654
rect 260186 477098 260422 477334
rect 260186 441418 260422 441654
rect 260186 441098 260422 441334
rect 260186 405418 260422 405654
rect 260186 405098 260422 405334
rect 260186 369418 260422 369654
rect 260186 369098 260422 369334
rect 260186 333418 260422 333654
rect 260186 333098 260422 333334
rect 256586 293818 256822 294054
rect 256586 293498 256822 293734
rect 256586 257818 256822 258054
rect 256586 257498 256822 257734
rect 256586 221818 256822 222054
rect 256586 221498 256822 221734
rect 256586 185818 256822 186054
rect 256586 185498 256822 185734
rect 256586 149818 256822 150054
rect 256586 149498 256822 149734
rect 256586 113818 256822 114054
rect 256586 113498 256822 113734
rect 256586 77818 256822 78054
rect 256586 77498 256822 77734
rect 256586 41818 256822 42054
rect 256586 41498 256822 41734
rect 256586 5818 256822 6054
rect 256586 5498 256822 5734
rect 256586 -2462 256822 -2226
rect 256586 -2782 256822 -2546
rect 260186 297418 260422 297654
rect 260186 297098 260422 297334
rect 260186 261418 260422 261654
rect 260186 261098 260422 261334
rect 260186 225418 260422 225654
rect 260186 225098 260422 225334
rect 260186 189418 260422 189654
rect 260186 189098 260422 189334
rect 260186 153418 260422 153654
rect 260186 153098 260422 153334
rect 260186 117418 260422 117654
rect 260186 117098 260422 117334
rect 260186 81418 260422 81654
rect 260186 81098 260422 81334
rect 260186 45418 260422 45654
rect 260186 45098 260422 45334
rect 260186 9418 260422 9654
rect 260186 9098 260422 9334
rect 260186 -4342 260422 -4106
rect 260186 -4662 260422 -4426
rect 281786 711182 282022 711418
rect 281786 710862 282022 711098
rect 278186 709302 278422 709538
rect 278186 708982 278422 709218
rect 274586 707422 274822 707658
rect 274586 707102 274822 707338
rect 263786 697018 264022 697254
rect 263786 696698 264022 696934
rect 263786 661018 264022 661254
rect 263786 660698 264022 660934
rect 263786 625018 264022 625254
rect 263786 624698 264022 624934
rect 263786 589018 264022 589254
rect 263786 588698 264022 588934
rect 263786 553018 264022 553254
rect 263786 552698 264022 552934
rect 263786 517018 264022 517254
rect 263786 516698 264022 516934
rect 263786 481018 264022 481254
rect 263786 480698 264022 480934
rect 263786 445018 264022 445254
rect 263786 444698 264022 444934
rect 270986 705542 271222 705778
rect 270986 705222 271222 705458
rect 270986 668218 271222 668454
rect 270986 667898 271222 668134
rect 270986 632218 271222 632454
rect 270986 631898 271222 632134
rect 270986 596218 271222 596454
rect 270986 595898 271222 596134
rect 270986 560218 271222 560454
rect 270986 559898 271222 560134
rect 270986 524218 271222 524454
rect 270986 523898 271222 524134
rect 270986 488218 271222 488454
rect 270986 487898 271222 488134
rect 270986 452218 271222 452454
rect 270986 451898 271222 452134
rect 270986 416218 271222 416454
rect 270986 415898 271222 416134
rect 263786 409018 264022 409254
rect 263786 408698 264022 408934
rect 263786 373018 264022 373254
rect 263786 372698 264022 372934
rect 263786 337018 264022 337254
rect 263786 336698 264022 336934
rect 263786 301018 264022 301254
rect 263786 300698 264022 300934
rect 263786 265018 264022 265254
rect 263786 264698 264022 264934
rect 263786 229018 264022 229254
rect 263786 228698 264022 228934
rect 270986 380218 271222 380454
rect 270986 379898 271222 380134
rect 270986 344218 271222 344454
rect 270986 343898 271222 344134
rect 270986 308218 271222 308454
rect 270986 307898 271222 308134
rect 270986 272218 271222 272454
rect 270986 271898 271222 272134
rect 270986 236218 271222 236454
rect 270986 235898 271222 236134
rect 263786 193018 264022 193254
rect 263786 192698 264022 192934
rect 263786 157018 264022 157254
rect 263786 156698 264022 156934
rect 263786 121018 264022 121254
rect 263786 120698 264022 120934
rect 263786 85018 264022 85254
rect 263786 84698 264022 84934
rect 263786 49018 264022 49254
rect 263786 48698 264022 48934
rect 263786 13018 264022 13254
rect 263786 12698 264022 12934
rect 245786 -7162 246022 -6926
rect 245786 -7482 246022 -7246
rect 270986 200218 271222 200454
rect 270986 199898 271222 200134
rect 270986 164218 271222 164454
rect 270986 163898 271222 164134
rect 270986 128218 271222 128454
rect 270986 127898 271222 128134
rect 270986 92218 271222 92454
rect 270986 91898 271222 92134
rect 270986 56218 271222 56454
rect 270986 55898 271222 56134
rect 270986 20218 271222 20454
rect 270986 19898 271222 20134
rect 270986 -1522 271222 -1286
rect 270986 -1842 271222 -1606
rect 274586 671818 274822 672054
rect 274586 671498 274822 671734
rect 274586 635818 274822 636054
rect 274586 635498 274822 635734
rect 274586 599818 274822 600054
rect 274586 599498 274822 599734
rect 274586 563818 274822 564054
rect 274586 563498 274822 563734
rect 274586 527818 274822 528054
rect 274586 527498 274822 527734
rect 274586 491818 274822 492054
rect 274586 491498 274822 491734
rect 274586 455818 274822 456054
rect 274586 455498 274822 455734
rect 274586 419818 274822 420054
rect 274586 419498 274822 419734
rect 274586 383818 274822 384054
rect 274586 383498 274822 383734
rect 274586 347818 274822 348054
rect 274586 347498 274822 347734
rect 274586 311818 274822 312054
rect 274586 311498 274822 311734
rect 274586 275818 274822 276054
rect 274586 275498 274822 275734
rect 274586 239818 274822 240054
rect 274586 239498 274822 239734
rect 274586 203818 274822 204054
rect 274586 203498 274822 203734
rect 274586 167818 274822 168054
rect 274586 167498 274822 167734
rect 274586 131818 274822 132054
rect 274586 131498 274822 131734
rect 274586 95818 274822 96054
rect 274586 95498 274822 95734
rect 274586 59818 274822 60054
rect 274586 59498 274822 59734
rect 274586 23818 274822 24054
rect 274586 23498 274822 23734
rect 274586 -3402 274822 -3166
rect 274586 -3722 274822 -3486
rect 278186 675418 278422 675654
rect 278186 675098 278422 675334
rect 278186 639418 278422 639654
rect 278186 639098 278422 639334
rect 278186 603418 278422 603654
rect 278186 603098 278422 603334
rect 278186 567418 278422 567654
rect 278186 567098 278422 567334
rect 278186 531418 278422 531654
rect 278186 531098 278422 531334
rect 278186 495418 278422 495654
rect 278186 495098 278422 495334
rect 278186 459418 278422 459654
rect 278186 459098 278422 459334
rect 278186 423418 278422 423654
rect 278186 423098 278422 423334
rect 278186 387418 278422 387654
rect 278186 387098 278422 387334
rect 278186 351418 278422 351654
rect 278186 351098 278422 351334
rect 278186 315418 278422 315654
rect 278186 315098 278422 315334
rect 278186 279418 278422 279654
rect 278186 279098 278422 279334
rect 278186 243418 278422 243654
rect 278186 243098 278422 243334
rect 278186 207418 278422 207654
rect 278186 207098 278422 207334
rect 278186 171418 278422 171654
rect 278186 171098 278422 171334
rect 278186 135418 278422 135654
rect 278186 135098 278422 135334
rect 278186 99418 278422 99654
rect 278186 99098 278422 99334
rect 278186 63418 278422 63654
rect 278186 63098 278422 63334
rect 278186 27418 278422 27654
rect 278186 27098 278422 27334
rect 278186 -5282 278422 -5046
rect 278186 -5602 278422 -5366
rect 299786 710242 300022 710478
rect 299786 709922 300022 710158
rect 296186 708362 296422 708598
rect 296186 708042 296422 708278
rect 292586 706482 292822 706718
rect 292586 706162 292822 706398
rect 281786 679018 282022 679254
rect 281786 678698 282022 678934
rect 281786 643018 282022 643254
rect 281786 642698 282022 642934
rect 281786 607018 282022 607254
rect 281786 606698 282022 606934
rect 281786 571018 282022 571254
rect 281786 570698 282022 570934
rect 281786 535018 282022 535254
rect 281786 534698 282022 534934
rect 281786 499018 282022 499254
rect 281786 498698 282022 498934
rect 281786 463018 282022 463254
rect 281786 462698 282022 462934
rect 281786 427018 282022 427254
rect 281786 426698 282022 426934
rect 281786 391018 282022 391254
rect 281786 390698 282022 390934
rect 288986 704602 289222 704838
rect 288986 704282 289222 704518
rect 288986 686218 289222 686454
rect 288986 685898 289222 686134
rect 288986 650218 289222 650454
rect 288986 649898 289222 650134
rect 288986 614218 289222 614454
rect 288986 613898 289222 614134
rect 288986 578218 289222 578454
rect 288986 577898 289222 578134
rect 288986 542218 289222 542454
rect 288986 541898 289222 542134
rect 288986 506218 289222 506454
rect 288986 505898 289222 506134
rect 288986 470218 289222 470454
rect 288986 469898 289222 470134
rect 288986 434218 289222 434454
rect 288986 433898 289222 434134
rect 288986 398218 289222 398454
rect 288986 397898 289222 398134
rect 281786 355018 282022 355254
rect 281786 354698 282022 354934
rect 281786 319018 282022 319254
rect 281786 318698 282022 318934
rect 281786 283018 282022 283254
rect 281786 282698 282022 282934
rect 281786 247018 282022 247254
rect 281786 246698 282022 246934
rect 281786 211018 282022 211254
rect 281786 210698 282022 210934
rect 281786 175018 282022 175254
rect 281786 174698 282022 174934
rect 281786 139018 282022 139254
rect 281786 138698 282022 138934
rect 281786 103018 282022 103254
rect 281786 102698 282022 102934
rect 281786 67018 282022 67254
rect 281786 66698 282022 66934
rect 281786 31018 282022 31254
rect 281786 30698 282022 30934
rect 263786 -6222 264022 -5986
rect 263786 -6542 264022 -6306
rect 288986 362218 289222 362454
rect 288986 361898 289222 362134
rect 288986 326218 289222 326454
rect 288986 325898 289222 326134
rect 288986 290218 289222 290454
rect 288986 289898 289222 290134
rect 288986 254218 289222 254454
rect 288986 253898 289222 254134
rect 288986 218218 289222 218454
rect 288986 217898 289222 218134
rect 288986 182218 289222 182454
rect 288986 181898 289222 182134
rect 288986 146218 289222 146454
rect 288986 145898 289222 146134
rect 288986 110218 289222 110454
rect 288986 109898 289222 110134
rect 288986 74218 289222 74454
rect 288986 73898 289222 74134
rect 288986 38218 289222 38454
rect 288986 37898 289222 38134
rect 288986 2218 289222 2454
rect 288986 1898 289222 2134
rect 288986 -582 289222 -346
rect 288986 -902 289222 -666
rect 292586 689818 292822 690054
rect 292586 689498 292822 689734
rect 292586 653818 292822 654054
rect 292586 653498 292822 653734
rect 292586 617818 292822 618054
rect 292586 617498 292822 617734
rect 292586 581818 292822 582054
rect 292586 581498 292822 581734
rect 292586 545818 292822 546054
rect 292586 545498 292822 545734
rect 292586 509818 292822 510054
rect 292586 509498 292822 509734
rect 292586 473818 292822 474054
rect 292586 473498 292822 473734
rect 292586 437818 292822 438054
rect 292586 437498 292822 437734
rect 292586 401818 292822 402054
rect 292586 401498 292822 401734
rect 292586 365818 292822 366054
rect 292586 365498 292822 365734
rect 292586 329818 292822 330054
rect 292586 329498 292822 329734
rect 292586 293818 292822 294054
rect 292586 293498 292822 293734
rect 292586 257818 292822 258054
rect 292586 257498 292822 257734
rect 292586 221818 292822 222054
rect 292586 221498 292822 221734
rect 292586 185818 292822 186054
rect 292586 185498 292822 185734
rect 292586 149818 292822 150054
rect 292586 149498 292822 149734
rect 292586 113818 292822 114054
rect 292586 113498 292822 113734
rect 292586 77818 292822 78054
rect 292586 77498 292822 77734
rect 292586 41818 292822 42054
rect 292586 41498 292822 41734
rect 292586 5818 292822 6054
rect 292586 5498 292822 5734
rect 292586 -2462 292822 -2226
rect 292586 -2782 292822 -2546
rect 296186 693418 296422 693654
rect 296186 693098 296422 693334
rect 296186 657418 296422 657654
rect 296186 657098 296422 657334
rect 296186 621418 296422 621654
rect 296186 621098 296422 621334
rect 296186 585418 296422 585654
rect 296186 585098 296422 585334
rect 296186 549418 296422 549654
rect 296186 549098 296422 549334
rect 296186 513418 296422 513654
rect 296186 513098 296422 513334
rect 296186 477418 296422 477654
rect 296186 477098 296422 477334
rect 296186 441418 296422 441654
rect 296186 441098 296422 441334
rect 296186 405418 296422 405654
rect 296186 405098 296422 405334
rect 296186 369418 296422 369654
rect 296186 369098 296422 369334
rect 296186 333418 296422 333654
rect 296186 333098 296422 333334
rect 317786 711182 318022 711418
rect 317786 710862 318022 711098
rect 314186 709302 314422 709538
rect 314186 708982 314422 709218
rect 310586 707422 310822 707658
rect 310586 707102 310822 707338
rect 299786 697018 300022 697254
rect 299786 696698 300022 696934
rect 299786 661018 300022 661254
rect 299786 660698 300022 660934
rect 299786 625018 300022 625254
rect 299786 624698 300022 624934
rect 299786 589018 300022 589254
rect 299786 588698 300022 588934
rect 299786 553018 300022 553254
rect 299786 552698 300022 552934
rect 299786 517018 300022 517254
rect 299786 516698 300022 516934
rect 299786 481018 300022 481254
rect 299786 480698 300022 480934
rect 299786 445018 300022 445254
rect 299786 444698 300022 444934
rect 299786 409018 300022 409254
rect 299786 408698 300022 408934
rect 299786 373018 300022 373254
rect 299786 372698 300022 372934
rect 299786 337018 300022 337254
rect 299786 336698 300022 336934
rect 299786 301018 300022 301254
rect 299786 300698 300022 300934
rect 296186 297418 296422 297654
rect 296186 297098 296422 297334
rect 296186 261418 296422 261654
rect 296186 261098 296422 261334
rect 296186 225418 296422 225654
rect 296186 225098 296422 225334
rect 296186 189418 296422 189654
rect 296186 189098 296422 189334
rect 296186 153418 296422 153654
rect 296186 153098 296422 153334
rect 296186 117418 296422 117654
rect 296186 117098 296422 117334
rect 296186 81418 296422 81654
rect 296186 81098 296422 81334
rect 296186 45418 296422 45654
rect 296186 45098 296422 45334
rect 296186 9418 296422 9654
rect 296186 9098 296422 9334
rect 296186 -4342 296422 -4106
rect 296186 -4662 296422 -4426
rect 299786 265018 300022 265254
rect 299786 264698 300022 264934
rect 299786 229018 300022 229254
rect 299786 228698 300022 228934
rect 299786 193018 300022 193254
rect 299786 192698 300022 192934
rect 299786 157018 300022 157254
rect 299786 156698 300022 156934
rect 299786 121018 300022 121254
rect 299786 120698 300022 120934
rect 299786 85018 300022 85254
rect 299786 84698 300022 84934
rect 299786 49018 300022 49254
rect 299786 48698 300022 48934
rect 299786 13018 300022 13254
rect 299786 12698 300022 12934
rect 281786 -7162 282022 -6926
rect 281786 -7482 282022 -7246
rect 306986 705542 307222 705778
rect 306986 705222 307222 705458
rect 306986 668218 307222 668454
rect 306986 667898 307222 668134
rect 306986 632218 307222 632454
rect 306986 631898 307222 632134
rect 306986 596218 307222 596454
rect 306986 595898 307222 596134
rect 306986 560218 307222 560454
rect 306986 559898 307222 560134
rect 306986 524218 307222 524454
rect 306986 523898 307222 524134
rect 306986 488218 307222 488454
rect 306986 487898 307222 488134
rect 306986 452218 307222 452454
rect 306986 451898 307222 452134
rect 306986 416218 307222 416454
rect 306986 415898 307222 416134
rect 306986 380218 307222 380454
rect 306986 379898 307222 380134
rect 306986 344218 307222 344454
rect 306986 343898 307222 344134
rect 306986 308218 307222 308454
rect 306986 307898 307222 308134
rect 306986 272218 307222 272454
rect 306986 271898 307222 272134
rect 306986 236218 307222 236454
rect 306986 235898 307222 236134
rect 306986 200218 307222 200454
rect 306986 199898 307222 200134
rect 306986 164218 307222 164454
rect 306986 163898 307222 164134
rect 306986 128218 307222 128454
rect 306986 127898 307222 128134
rect 306986 92218 307222 92454
rect 306986 91898 307222 92134
rect 306986 56218 307222 56454
rect 306986 55898 307222 56134
rect 306986 20218 307222 20454
rect 306986 19898 307222 20134
rect 306986 -1522 307222 -1286
rect 306986 -1842 307222 -1606
rect 310586 671818 310822 672054
rect 310586 671498 310822 671734
rect 310586 635818 310822 636054
rect 310586 635498 310822 635734
rect 310586 599818 310822 600054
rect 310586 599498 310822 599734
rect 310586 563818 310822 564054
rect 310586 563498 310822 563734
rect 310586 527818 310822 528054
rect 310586 527498 310822 527734
rect 310586 491818 310822 492054
rect 310586 491498 310822 491734
rect 310586 455818 310822 456054
rect 310586 455498 310822 455734
rect 310586 419818 310822 420054
rect 310586 419498 310822 419734
rect 310586 383818 310822 384054
rect 310586 383498 310822 383734
rect 310586 347818 310822 348054
rect 310586 347498 310822 347734
rect 310586 311818 310822 312054
rect 310586 311498 310822 311734
rect 310586 275818 310822 276054
rect 310586 275498 310822 275734
rect 310586 239818 310822 240054
rect 310586 239498 310822 239734
rect 310586 203818 310822 204054
rect 310586 203498 310822 203734
rect 310586 167818 310822 168054
rect 310586 167498 310822 167734
rect 310586 131818 310822 132054
rect 310586 131498 310822 131734
rect 310586 95818 310822 96054
rect 310586 95498 310822 95734
rect 310586 59818 310822 60054
rect 310586 59498 310822 59734
rect 310586 23818 310822 24054
rect 310586 23498 310822 23734
rect 310586 -3402 310822 -3166
rect 310586 -3722 310822 -3486
rect 314186 675418 314422 675654
rect 314186 675098 314422 675334
rect 314186 639418 314422 639654
rect 314186 639098 314422 639334
rect 314186 603418 314422 603654
rect 314186 603098 314422 603334
rect 314186 567418 314422 567654
rect 314186 567098 314422 567334
rect 314186 531418 314422 531654
rect 314186 531098 314422 531334
rect 314186 495418 314422 495654
rect 314186 495098 314422 495334
rect 314186 459418 314422 459654
rect 314186 459098 314422 459334
rect 314186 423418 314422 423654
rect 314186 423098 314422 423334
rect 314186 387418 314422 387654
rect 314186 387098 314422 387334
rect 314186 351418 314422 351654
rect 314186 351098 314422 351334
rect 314186 315418 314422 315654
rect 314186 315098 314422 315334
rect 314186 279418 314422 279654
rect 314186 279098 314422 279334
rect 314186 243418 314422 243654
rect 314186 243098 314422 243334
rect 314186 207418 314422 207654
rect 314186 207098 314422 207334
rect 314186 171418 314422 171654
rect 314186 171098 314422 171334
rect 314186 135418 314422 135654
rect 314186 135098 314422 135334
rect 314186 99418 314422 99654
rect 314186 99098 314422 99334
rect 314186 63418 314422 63654
rect 314186 63098 314422 63334
rect 314186 27418 314422 27654
rect 314186 27098 314422 27334
rect 314186 -5282 314422 -5046
rect 314186 -5602 314422 -5366
rect 335786 710242 336022 710478
rect 335786 709922 336022 710158
rect 332186 708362 332422 708598
rect 332186 708042 332422 708278
rect 328586 706482 328822 706718
rect 328586 706162 328822 706398
rect 317786 679018 318022 679254
rect 317786 678698 318022 678934
rect 317786 643018 318022 643254
rect 317786 642698 318022 642934
rect 317786 607018 318022 607254
rect 317786 606698 318022 606934
rect 317786 571018 318022 571254
rect 317786 570698 318022 570934
rect 317786 535018 318022 535254
rect 317786 534698 318022 534934
rect 317786 499018 318022 499254
rect 317786 498698 318022 498934
rect 317786 463018 318022 463254
rect 317786 462698 318022 462934
rect 317786 427018 318022 427254
rect 317786 426698 318022 426934
rect 317786 391018 318022 391254
rect 317786 390698 318022 390934
rect 317786 355018 318022 355254
rect 317786 354698 318022 354934
rect 317786 319018 318022 319254
rect 317786 318698 318022 318934
rect 317786 283018 318022 283254
rect 317786 282698 318022 282934
rect 317786 247018 318022 247254
rect 317786 246698 318022 246934
rect 317786 211018 318022 211254
rect 317786 210698 318022 210934
rect 317786 175018 318022 175254
rect 317786 174698 318022 174934
rect 317786 139018 318022 139254
rect 317786 138698 318022 138934
rect 317786 103018 318022 103254
rect 317786 102698 318022 102934
rect 317786 67018 318022 67254
rect 317786 66698 318022 66934
rect 317786 31018 318022 31254
rect 317786 30698 318022 30934
rect 299786 -6222 300022 -5986
rect 299786 -6542 300022 -6306
rect 324986 704602 325222 704838
rect 324986 704282 325222 704518
rect 324986 686218 325222 686454
rect 324986 685898 325222 686134
rect 324986 650218 325222 650454
rect 324986 649898 325222 650134
rect 324986 614218 325222 614454
rect 324986 613898 325222 614134
rect 324986 578218 325222 578454
rect 324986 577898 325222 578134
rect 324986 542218 325222 542454
rect 324986 541898 325222 542134
rect 324986 506218 325222 506454
rect 324986 505898 325222 506134
rect 324986 470218 325222 470454
rect 324986 469898 325222 470134
rect 324986 434218 325222 434454
rect 324986 433898 325222 434134
rect 324986 398218 325222 398454
rect 324986 397898 325222 398134
rect 324986 362218 325222 362454
rect 324986 361898 325222 362134
rect 324986 326218 325222 326454
rect 324986 325898 325222 326134
rect 324986 290218 325222 290454
rect 324986 289898 325222 290134
rect 324986 254218 325222 254454
rect 324986 253898 325222 254134
rect 324986 218218 325222 218454
rect 324986 217898 325222 218134
rect 324986 182218 325222 182454
rect 324986 181898 325222 182134
rect 324986 146218 325222 146454
rect 324986 145898 325222 146134
rect 324986 110218 325222 110454
rect 324986 109898 325222 110134
rect 324986 74218 325222 74454
rect 324986 73898 325222 74134
rect 324986 38218 325222 38454
rect 324986 37898 325222 38134
rect 324986 2218 325222 2454
rect 324986 1898 325222 2134
rect 324986 -582 325222 -346
rect 324986 -902 325222 -666
rect 328586 689818 328822 690054
rect 328586 689498 328822 689734
rect 328586 653818 328822 654054
rect 328586 653498 328822 653734
rect 328586 617818 328822 618054
rect 328586 617498 328822 617734
rect 328586 581818 328822 582054
rect 328586 581498 328822 581734
rect 328586 545818 328822 546054
rect 328586 545498 328822 545734
rect 328586 509818 328822 510054
rect 328586 509498 328822 509734
rect 328586 473818 328822 474054
rect 328586 473498 328822 473734
rect 328586 437818 328822 438054
rect 328586 437498 328822 437734
rect 328586 401818 328822 402054
rect 328586 401498 328822 401734
rect 328586 365818 328822 366054
rect 328586 365498 328822 365734
rect 328586 329818 328822 330054
rect 328586 329498 328822 329734
rect 328586 293818 328822 294054
rect 328586 293498 328822 293734
rect 328586 257818 328822 258054
rect 328586 257498 328822 257734
rect 328586 221818 328822 222054
rect 328586 221498 328822 221734
rect 328586 185818 328822 186054
rect 328586 185498 328822 185734
rect 328586 149818 328822 150054
rect 328586 149498 328822 149734
rect 328586 113818 328822 114054
rect 328586 113498 328822 113734
rect 328586 77818 328822 78054
rect 328586 77498 328822 77734
rect 328586 41818 328822 42054
rect 328586 41498 328822 41734
rect 328586 5818 328822 6054
rect 328586 5498 328822 5734
rect 328586 -2462 328822 -2226
rect 328586 -2782 328822 -2546
rect 332186 693418 332422 693654
rect 332186 693098 332422 693334
rect 332186 657418 332422 657654
rect 332186 657098 332422 657334
rect 332186 621418 332422 621654
rect 332186 621098 332422 621334
rect 332186 585418 332422 585654
rect 332186 585098 332422 585334
rect 332186 549418 332422 549654
rect 332186 549098 332422 549334
rect 332186 513418 332422 513654
rect 332186 513098 332422 513334
rect 332186 477418 332422 477654
rect 332186 477098 332422 477334
rect 332186 441418 332422 441654
rect 332186 441098 332422 441334
rect 332186 405418 332422 405654
rect 332186 405098 332422 405334
rect 332186 369418 332422 369654
rect 332186 369098 332422 369334
rect 332186 333418 332422 333654
rect 332186 333098 332422 333334
rect 332186 297418 332422 297654
rect 332186 297098 332422 297334
rect 332186 261418 332422 261654
rect 332186 261098 332422 261334
rect 332186 225418 332422 225654
rect 332186 225098 332422 225334
rect 332186 189418 332422 189654
rect 332186 189098 332422 189334
rect 332186 153418 332422 153654
rect 332186 153098 332422 153334
rect 332186 117418 332422 117654
rect 332186 117098 332422 117334
rect 332186 81418 332422 81654
rect 332186 81098 332422 81334
rect 332186 45418 332422 45654
rect 332186 45098 332422 45334
rect 332186 9418 332422 9654
rect 332186 9098 332422 9334
rect 332186 -4342 332422 -4106
rect 332186 -4662 332422 -4426
rect 353786 711182 354022 711418
rect 353786 710862 354022 711098
rect 350186 709302 350422 709538
rect 350186 708982 350422 709218
rect 346586 707422 346822 707658
rect 346586 707102 346822 707338
rect 335786 697018 336022 697254
rect 335786 696698 336022 696934
rect 335786 661018 336022 661254
rect 335786 660698 336022 660934
rect 335786 625018 336022 625254
rect 335786 624698 336022 624934
rect 335786 589018 336022 589254
rect 335786 588698 336022 588934
rect 335786 553018 336022 553254
rect 335786 552698 336022 552934
rect 335786 517018 336022 517254
rect 335786 516698 336022 516934
rect 335786 481018 336022 481254
rect 335786 480698 336022 480934
rect 335786 445018 336022 445254
rect 335786 444698 336022 444934
rect 335786 409018 336022 409254
rect 335786 408698 336022 408934
rect 335786 373018 336022 373254
rect 335786 372698 336022 372934
rect 335786 337018 336022 337254
rect 335786 336698 336022 336934
rect 335786 301018 336022 301254
rect 335786 300698 336022 300934
rect 335786 265018 336022 265254
rect 335786 264698 336022 264934
rect 335786 229018 336022 229254
rect 335786 228698 336022 228934
rect 335786 193018 336022 193254
rect 335786 192698 336022 192934
rect 335786 157018 336022 157254
rect 335786 156698 336022 156934
rect 335786 121018 336022 121254
rect 335786 120698 336022 120934
rect 335786 85018 336022 85254
rect 335786 84698 336022 84934
rect 335786 49018 336022 49254
rect 335786 48698 336022 48934
rect 335786 13018 336022 13254
rect 335786 12698 336022 12934
rect 317786 -7162 318022 -6926
rect 317786 -7482 318022 -7246
rect 342986 705542 343222 705778
rect 342986 705222 343222 705458
rect 342986 668218 343222 668454
rect 342986 667898 343222 668134
rect 342986 632218 343222 632454
rect 342986 631898 343222 632134
rect 342986 596218 343222 596454
rect 342986 595898 343222 596134
rect 342986 560218 343222 560454
rect 342986 559898 343222 560134
rect 342986 524218 343222 524454
rect 342986 523898 343222 524134
rect 342986 488218 343222 488454
rect 342986 487898 343222 488134
rect 342986 452218 343222 452454
rect 342986 451898 343222 452134
rect 342986 416218 343222 416454
rect 342986 415898 343222 416134
rect 342986 380218 343222 380454
rect 342986 379898 343222 380134
rect 342986 344218 343222 344454
rect 342986 343898 343222 344134
rect 342986 308218 343222 308454
rect 342986 307898 343222 308134
rect 342986 272218 343222 272454
rect 342986 271898 343222 272134
rect 342986 236218 343222 236454
rect 342986 235898 343222 236134
rect 342986 200218 343222 200454
rect 342986 199898 343222 200134
rect 342986 164218 343222 164454
rect 342986 163898 343222 164134
rect 342986 128218 343222 128454
rect 342986 127898 343222 128134
rect 342986 92218 343222 92454
rect 342986 91898 343222 92134
rect 342986 56218 343222 56454
rect 342986 55898 343222 56134
rect 342986 20218 343222 20454
rect 342986 19898 343222 20134
rect 342986 -1522 343222 -1286
rect 342986 -1842 343222 -1606
rect 346586 671818 346822 672054
rect 346586 671498 346822 671734
rect 346586 635818 346822 636054
rect 346586 635498 346822 635734
rect 346586 599818 346822 600054
rect 346586 599498 346822 599734
rect 346586 563818 346822 564054
rect 346586 563498 346822 563734
rect 346586 527818 346822 528054
rect 346586 527498 346822 527734
rect 346586 491818 346822 492054
rect 346586 491498 346822 491734
rect 346586 455818 346822 456054
rect 346586 455498 346822 455734
rect 346586 419818 346822 420054
rect 346586 419498 346822 419734
rect 346586 383818 346822 384054
rect 346586 383498 346822 383734
rect 346586 347818 346822 348054
rect 346586 347498 346822 347734
rect 346586 311818 346822 312054
rect 346586 311498 346822 311734
rect 346586 275818 346822 276054
rect 346586 275498 346822 275734
rect 346586 239818 346822 240054
rect 346586 239498 346822 239734
rect 346586 203818 346822 204054
rect 346586 203498 346822 203734
rect 346586 167818 346822 168054
rect 346586 167498 346822 167734
rect 346586 131818 346822 132054
rect 346586 131498 346822 131734
rect 346586 95818 346822 96054
rect 346586 95498 346822 95734
rect 346586 59818 346822 60054
rect 346586 59498 346822 59734
rect 346586 23818 346822 24054
rect 346586 23498 346822 23734
rect 346586 -3402 346822 -3166
rect 346586 -3722 346822 -3486
rect 350186 675418 350422 675654
rect 350186 675098 350422 675334
rect 350186 639418 350422 639654
rect 350186 639098 350422 639334
rect 350186 603418 350422 603654
rect 350186 603098 350422 603334
rect 350186 567418 350422 567654
rect 350186 567098 350422 567334
rect 350186 531418 350422 531654
rect 350186 531098 350422 531334
rect 350186 495418 350422 495654
rect 350186 495098 350422 495334
rect 350186 459418 350422 459654
rect 350186 459098 350422 459334
rect 350186 423418 350422 423654
rect 350186 423098 350422 423334
rect 350186 387418 350422 387654
rect 350186 387098 350422 387334
rect 350186 351418 350422 351654
rect 350186 351098 350422 351334
rect 350186 315418 350422 315654
rect 350186 315098 350422 315334
rect 350186 279418 350422 279654
rect 350186 279098 350422 279334
rect 350186 243418 350422 243654
rect 350186 243098 350422 243334
rect 350186 207418 350422 207654
rect 350186 207098 350422 207334
rect 350186 171418 350422 171654
rect 350186 171098 350422 171334
rect 350186 135418 350422 135654
rect 350186 135098 350422 135334
rect 350186 99418 350422 99654
rect 350186 99098 350422 99334
rect 350186 63418 350422 63654
rect 350186 63098 350422 63334
rect 350186 27418 350422 27654
rect 350186 27098 350422 27334
rect 350186 -5282 350422 -5046
rect 350186 -5602 350422 -5366
rect 371786 710242 372022 710478
rect 371786 709922 372022 710158
rect 368186 708362 368422 708598
rect 368186 708042 368422 708278
rect 364586 706482 364822 706718
rect 364586 706162 364822 706398
rect 353786 679018 354022 679254
rect 353786 678698 354022 678934
rect 353786 643018 354022 643254
rect 353786 642698 354022 642934
rect 353786 607018 354022 607254
rect 353786 606698 354022 606934
rect 353786 571018 354022 571254
rect 353786 570698 354022 570934
rect 353786 535018 354022 535254
rect 353786 534698 354022 534934
rect 353786 499018 354022 499254
rect 353786 498698 354022 498934
rect 353786 463018 354022 463254
rect 353786 462698 354022 462934
rect 353786 427018 354022 427254
rect 353786 426698 354022 426934
rect 353786 391018 354022 391254
rect 353786 390698 354022 390934
rect 353786 355018 354022 355254
rect 353786 354698 354022 354934
rect 353786 319018 354022 319254
rect 353786 318698 354022 318934
rect 353786 283018 354022 283254
rect 353786 282698 354022 282934
rect 353786 247018 354022 247254
rect 353786 246698 354022 246934
rect 353786 211018 354022 211254
rect 353786 210698 354022 210934
rect 353786 175018 354022 175254
rect 353786 174698 354022 174934
rect 353786 139018 354022 139254
rect 353786 138698 354022 138934
rect 353786 103018 354022 103254
rect 353786 102698 354022 102934
rect 353786 67018 354022 67254
rect 353786 66698 354022 66934
rect 353786 31018 354022 31254
rect 353786 30698 354022 30934
rect 335786 -6222 336022 -5986
rect 335786 -6542 336022 -6306
rect 360986 704602 361222 704838
rect 360986 704282 361222 704518
rect 360986 686218 361222 686454
rect 360986 685898 361222 686134
rect 360986 650218 361222 650454
rect 360986 649898 361222 650134
rect 360986 614218 361222 614454
rect 360986 613898 361222 614134
rect 360986 578218 361222 578454
rect 360986 577898 361222 578134
rect 360986 542218 361222 542454
rect 360986 541898 361222 542134
rect 360986 506218 361222 506454
rect 360986 505898 361222 506134
rect 360986 470218 361222 470454
rect 360986 469898 361222 470134
rect 360986 434218 361222 434454
rect 360986 433898 361222 434134
rect 360986 398218 361222 398454
rect 360986 397898 361222 398134
rect 360986 362218 361222 362454
rect 360986 361898 361222 362134
rect 360986 326218 361222 326454
rect 360986 325898 361222 326134
rect 360986 290218 361222 290454
rect 360986 289898 361222 290134
rect 360986 254218 361222 254454
rect 360986 253898 361222 254134
rect 360986 218218 361222 218454
rect 360986 217898 361222 218134
rect 360986 182218 361222 182454
rect 360986 181898 361222 182134
rect 360986 146218 361222 146454
rect 360986 145898 361222 146134
rect 360986 110218 361222 110454
rect 360986 109898 361222 110134
rect 360986 74218 361222 74454
rect 360986 73898 361222 74134
rect 360986 38218 361222 38454
rect 360986 37898 361222 38134
rect 360986 2218 361222 2454
rect 360986 1898 361222 2134
rect 360986 -582 361222 -346
rect 360986 -902 361222 -666
rect 364586 689818 364822 690054
rect 364586 689498 364822 689734
rect 364586 653818 364822 654054
rect 364586 653498 364822 653734
rect 364586 617818 364822 618054
rect 364586 617498 364822 617734
rect 364586 581818 364822 582054
rect 364586 581498 364822 581734
rect 364586 545818 364822 546054
rect 364586 545498 364822 545734
rect 364586 509818 364822 510054
rect 364586 509498 364822 509734
rect 364586 473818 364822 474054
rect 364586 473498 364822 473734
rect 364586 437818 364822 438054
rect 364586 437498 364822 437734
rect 364586 401818 364822 402054
rect 364586 401498 364822 401734
rect 364586 365818 364822 366054
rect 364586 365498 364822 365734
rect 364586 329818 364822 330054
rect 364586 329498 364822 329734
rect 364586 293818 364822 294054
rect 364586 293498 364822 293734
rect 364586 257818 364822 258054
rect 364586 257498 364822 257734
rect 364586 221818 364822 222054
rect 364586 221498 364822 221734
rect 364586 185818 364822 186054
rect 364586 185498 364822 185734
rect 364586 149818 364822 150054
rect 364586 149498 364822 149734
rect 364586 113818 364822 114054
rect 364586 113498 364822 113734
rect 364586 77818 364822 78054
rect 364586 77498 364822 77734
rect 364586 41818 364822 42054
rect 364586 41498 364822 41734
rect 364586 5818 364822 6054
rect 364586 5498 364822 5734
rect 364586 -2462 364822 -2226
rect 364586 -2782 364822 -2546
rect 368186 693418 368422 693654
rect 368186 693098 368422 693334
rect 368186 657418 368422 657654
rect 368186 657098 368422 657334
rect 368186 621418 368422 621654
rect 368186 621098 368422 621334
rect 368186 585418 368422 585654
rect 368186 585098 368422 585334
rect 368186 549418 368422 549654
rect 368186 549098 368422 549334
rect 368186 513418 368422 513654
rect 368186 513098 368422 513334
rect 368186 477418 368422 477654
rect 368186 477098 368422 477334
rect 368186 441418 368422 441654
rect 368186 441098 368422 441334
rect 368186 405418 368422 405654
rect 368186 405098 368422 405334
rect 368186 369418 368422 369654
rect 368186 369098 368422 369334
rect 368186 333418 368422 333654
rect 368186 333098 368422 333334
rect 368186 297418 368422 297654
rect 368186 297098 368422 297334
rect 368186 261418 368422 261654
rect 368186 261098 368422 261334
rect 368186 225418 368422 225654
rect 368186 225098 368422 225334
rect 368186 189418 368422 189654
rect 368186 189098 368422 189334
rect 368186 153418 368422 153654
rect 368186 153098 368422 153334
rect 368186 117418 368422 117654
rect 368186 117098 368422 117334
rect 368186 81418 368422 81654
rect 368186 81098 368422 81334
rect 368186 45418 368422 45654
rect 368186 45098 368422 45334
rect 368186 9418 368422 9654
rect 368186 9098 368422 9334
rect 368186 -4342 368422 -4106
rect 368186 -4662 368422 -4426
rect 389786 711182 390022 711418
rect 389786 710862 390022 711098
rect 386186 709302 386422 709538
rect 386186 708982 386422 709218
rect 382586 707422 382822 707658
rect 382586 707102 382822 707338
rect 371786 697018 372022 697254
rect 371786 696698 372022 696934
rect 371786 661018 372022 661254
rect 371786 660698 372022 660934
rect 371786 625018 372022 625254
rect 371786 624698 372022 624934
rect 371786 589018 372022 589254
rect 371786 588698 372022 588934
rect 371786 553018 372022 553254
rect 371786 552698 372022 552934
rect 371786 517018 372022 517254
rect 371786 516698 372022 516934
rect 371786 481018 372022 481254
rect 371786 480698 372022 480934
rect 371786 445018 372022 445254
rect 371786 444698 372022 444934
rect 371786 409018 372022 409254
rect 371786 408698 372022 408934
rect 371786 373018 372022 373254
rect 371786 372698 372022 372934
rect 371786 337018 372022 337254
rect 371786 336698 372022 336934
rect 371786 301018 372022 301254
rect 371786 300698 372022 300934
rect 371786 265018 372022 265254
rect 371786 264698 372022 264934
rect 371786 229018 372022 229254
rect 371786 228698 372022 228934
rect 371786 193018 372022 193254
rect 371786 192698 372022 192934
rect 371786 157018 372022 157254
rect 371786 156698 372022 156934
rect 371786 121018 372022 121254
rect 371786 120698 372022 120934
rect 371786 85018 372022 85254
rect 371786 84698 372022 84934
rect 371786 49018 372022 49254
rect 371786 48698 372022 48934
rect 371786 13018 372022 13254
rect 371786 12698 372022 12934
rect 353786 -7162 354022 -6926
rect 353786 -7482 354022 -7246
rect 378986 705542 379222 705778
rect 378986 705222 379222 705458
rect 378986 668218 379222 668454
rect 378986 667898 379222 668134
rect 378986 632218 379222 632454
rect 378986 631898 379222 632134
rect 378986 596218 379222 596454
rect 378986 595898 379222 596134
rect 382586 671818 382822 672054
rect 382586 671498 382822 671734
rect 382586 635818 382822 636054
rect 382586 635498 382822 635734
rect 382586 599818 382822 600054
rect 382586 599498 382822 599734
rect 378986 560218 379222 560454
rect 378986 559898 379222 560134
rect 378986 524218 379222 524454
rect 378986 523898 379222 524134
rect 378986 488218 379222 488454
rect 378986 487898 379222 488134
rect 378986 452218 379222 452454
rect 378986 451898 379222 452134
rect 378986 416218 379222 416454
rect 378986 415898 379222 416134
rect 382586 563818 382822 564054
rect 382586 563498 382822 563734
rect 382586 527818 382822 528054
rect 382586 527498 382822 527734
rect 382586 491818 382822 492054
rect 382586 491498 382822 491734
rect 382586 455818 382822 456054
rect 382586 455498 382822 455734
rect 382586 419818 382822 420054
rect 382586 419498 382822 419734
rect 378986 380218 379222 380454
rect 378986 379898 379222 380134
rect 378986 344218 379222 344454
rect 378986 343898 379222 344134
rect 378986 308218 379222 308454
rect 378986 307898 379222 308134
rect 378986 272218 379222 272454
rect 378986 271898 379222 272134
rect 378986 236218 379222 236454
rect 378986 235898 379222 236134
rect 378986 200218 379222 200454
rect 378986 199898 379222 200134
rect 378986 164218 379222 164454
rect 378986 163898 379222 164134
rect 378986 128218 379222 128454
rect 378986 127898 379222 128134
rect 378986 92218 379222 92454
rect 378986 91898 379222 92134
rect 378986 56218 379222 56454
rect 378986 55898 379222 56134
rect 378986 20218 379222 20454
rect 378986 19898 379222 20134
rect 378986 -1522 379222 -1286
rect 378986 -1842 379222 -1606
rect 382586 383818 382822 384054
rect 382586 383498 382822 383734
rect 382586 347818 382822 348054
rect 382586 347498 382822 347734
rect 382586 311818 382822 312054
rect 382586 311498 382822 311734
rect 382586 275818 382822 276054
rect 382586 275498 382822 275734
rect 382586 239818 382822 240054
rect 382586 239498 382822 239734
rect 382586 203818 382822 204054
rect 382586 203498 382822 203734
rect 382586 167818 382822 168054
rect 382586 167498 382822 167734
rect 382586 131818 382822 132054
rect 382586 131498 382822 131734
rect 382586 95818 382822 96054
rect 382586 95498 382822 95734
rect 382586 59818 382822 60054
rect 382586 59498 382822 59734
rect 382586 23818 382822 24054
rect 382586 23498 382822 23734
rect 382586 -3402 382822 -3166
rect 382586 -3722 382822 -3486
rect 386186 675418 386422 675654
rect 386186 675098 386422 675334
rect 386186 639418 386422 639654
rect 386186 639098 386422 639334
rect 386186 603418 386422 603654
rect 386186 603098 386422 603334
rect 386186 567418 386422 567654
rect 386186 567098 386422 567334
rect 386186 531418 386422 531654
rect 386186 531098 386422 531334
rect 386186 495418 386422 495654
rect 386186 495098 386422 495334
rect 386186 459418 386422 459654
rect 386186 459098 386422 459334
rect 386186 423418 386422 423654
rect 386186 423098 386422 423334
rect 386186 387418 386422 387654
rect 386186 387098 386422 387334
rect 386186 351418 386422 351654
rect 386186 351098 386422 351334
rect 386186 315418 386422 315654
rect 386186 315098 386422 315334
rect 386186 279418 386422 279654
rect 386186 279098 386422 279334
rect 386186 243418 386422 243654
rect 386186 243098 386422 243334
rect 386186 207418 386422 207654
rect 386186 207098 386422 207334
rect 386186 171418 386422 171654
rect 386186 171098 386422 171334
rect 386186 135418 386422 135654
rect 386186 135098 386422 135334
rect 386186 99418 386422 99654
rect 386186 99098 386422 99334
rect 386186 63418 386422 63654
rect 386186 63098 386422 63334
rect 386186 27418 386422 27654
rect 386186 27098 386422 27334
rect 386186 -5282 386422 -5046
rect 386186 -5602 386422 -5366
rect 407786 710242 408022 710478
rect 407786 709922 408022 710158
rect 404186 708362 404422 708598
rect 404186 708042 404422 708278
rect 400586 706482 400822 706718
rect 400586 706162 400822 706398
rect 389786 679018 390022 679254
rect 389786 678698 390022 678934
rect 389786 643018 390022 643254
rect 389786 642698 390022 642934
rect 389786 607018 390022 607254
rect 389786 606698 390022 606934
rect 389786 571018 390022 571254
rect 389786 570698 390022 570934
rect 389786 535018 390022 535254
rect 389786 534698 390022 534934
rect 389786 499018 390022 499254
rect 389786 498698 390022 498934
rect 389786 463018 390022 463254
rect 389786 462698 390022 462934
rect 389786 427018 390022 427254
rect 389786 426698 390022 426934
rect 389786 391018 390022 391254
rect 389786 390698 390022 390934
rect 389786 355018 390022 355254
rect 389786 354698 390022 354934
rect 389786 319018 390022 319254
rect 389786 318698 390022 318934
rect 396986 704602 397222 704838
rect 396986 704282 397222 704518
rect 396986 686218 397222 686454
rect 396986 685898 397222 686134
rect 396986 650218 397222 650454
rect 396986 649898 397222 650134
rect 396986 614218 397222 614454
rect 396986 613898 397222 614134
rect 396986 578218 397222 578454
rect 396986 577898 397222 578134
rect 396986 542218 397222 542454
rect 396986 541898 397222 542134
rect 396986 506218 397222 506454
rect 396986 505898 397222 506134
rect 396986 470218 397222 470454
rect 396986 469898 397222 470134
rect 396986 434218 397222 434454
rect 396986 433898 397222 434134
rect 396986 398218 397222 398454
rect 396986 397898 397222 398134
rect 396986 362218 397222 362454
rect 396986 361898 397222 362134
rect 396986 326218 397222 326454
rect 396986 325898 397222 326134
rect 396986 290218 397222 290454
rect 396986 289898 397222 290134
rect 389786 283018 390022 283254
rect 389786 282698 390022 282934
rect 389786 247018 390022 247254
rect 389786 246698 390022 246934
rect 389786 211018 390022 211254
rect 389786 210698 390022 210934
rect 389786 175018 390022 175254
rect 389786 174698 390022 174934
rect 389786 139018 390022 139254
rect 389786 138698 390022 138934
rect 389786 103018 390022 103254
rect 389786 102698 390022 102934
rect 389786 67018 390022 67254
rect 389786 66698 390022 66934
rect 389786 31018 390022 31254
rect 389786 30698 390022 30934
rect 371786 -6222 372022 -5986
rect 371786 -6542 372022 -6306
rect 396986 254218 397222 254454
rect 396986 253898 397222 254134
rect 396986 218218 397222 218454
rect 396986 217898 397222 218134
rect 396986 182218 397222 182454
rect 396986 181898 397222 182134
rect 396986 146218 397222 146454
rect 396986 145898 397222 146134
rect 396986 110218 397222 110454
rect 396986 109898 397222 110134
rect 396986 74218 397222 74454
rect 396986 73898 397222 74134
rect 396986 38218 397222 38454
rect 396986 37898 397222 38134
rect 396986 2218 397222 2454
rect 396986 1898 397222 2134
rect 396986 -582 397222 -346
rect 396986 -902 397222 -666
rect 400586 689818 400822 690054
rect 400586 689498 400822 689734
rect 400586 653818 400822 654054
rect 400586 653498 400822 653734
rect 400586 617818 400822 618054
rect 400586 617498 400822 617734
rect 400586 581818 400822 582054
rect 400586 581498 400822 581734
rect 400586 545818 400822 546054
rect 400586 545498 400822 545734
rect 400586 509818 400822 510054
rect 400586 509498 400822 509734
rect 400586 473818 400822 474054
rect 400586 473498 400822 473734
rect 400586 437818 400822 438054
rect 400586 437498 400822 437734
rect 400586 401818 400822 402054
rect 400586 401498 400822 401734
rect 400586 365818 400822 366054
rect 400586 365498 400822 365734
rect 400586 329818 400822 330054
rect 400586 329498 400822 329734
rect 400586 293818 400822 294054
rect 400586 293498 400822 293734
rect 400586 257818 400822 258054
rect 400586 257498 400822 257734
rect 400586 221818 400822 222054
rect 400586 221498 400822 221734
rect 400586 185818 400822 186054
rect 400586 185498 400822 185734
rect 400586 149818 400822 150054
rect 400586 149498 400822 149734
rect 400586 113818 400822 114054
rect 400586 113498 400822 113734
rect 400586 77818 400822 78054
rect 400586 77498 400822 77734
rect 400586 41818 400822 42054
rect 400586 41498 400822 41734
rect 400586 5818 400822 6054
rect 400586 5498 400822 5734
rect 400586 -2462 400822 -2226
rect 400586 -2782 400822 -2546
rect 404186 693418 404422 693654
rect 404186 693098 404422 693334
rect 404186 657418 404422 657654
rect 404186 657098 404422 657334
rect 404186 621418 404422 621654
rect 404186 621098 404422 621334
rect 404186 585418 404422 585654
rect 404186 585098 404422 585334
rect 404186 549418 404422 549654
rect 404186 549098 404422 549334
rect 404186 513418 404422 513654
rect 404186 513098 404422 513334
rect 404186 477418 404422 477654
rect 404186 477098 404422 477334
rect 404186 441418 404422 441654
rect 404186 441098 404422 441334
rect 404186 405418 404422 405654
rect 404186 405098 404422 405334
rect 404186 369418 404422 369654
rect 404186 369098 404422 369334
rect 404186 333418 404422 333654
rect 404186 333098 404422 333334
rect 404186 297418 404422 297654
rect 404186 297098 404422 297334
rect 404186 261418 404422 261654
rect 404186 261098 404422 261334
rect 404186 225418 404422 225654
rect 404186 225098 404422 225334
rect 404186 189418 404422 189654
rect 404186 189098 404422 189334
rect 404186 153418 404422 153654
rect 404186 153098 404422 153334
rect 404186 117418 404422 117654
rect 404186 117098 404422 117334
rect 404186 81418 404422 81654
rect 404186 81098 404422 81334
rect 404186 45418 404422 45654
rect 404186 45098 404422 45334
rect 404186 9418 404422 9654
rect 404186 9098 404422 9334
rect 404186 -4342 404422 -4106
rect 404186 -4662 404422 -4426
rect 425786 711182 426022 711418
rect 425786 710862 426022 711098
rect 422186 709302 422422 709538
rect 422186 708982 422422 709218
rect 418586 707422 418822 707658
rect 418586 707102 418822 707338
rect 407786 697018 408022 697254
rect 407786 696698 408022 696934
rect 407786 661018 408022 661254
rect 407786 660698 408022 660934
rect 407786 625018 408022 625254
rect 407786 624698 408022 624934
rect 407786 589018 408022 589254
rect 407786 588698 408022 588934
rect 407786 553018 408022 553254
rect 407786 552698 408022 552934
rect 407786 517018 408022 517254
rect 407786 516698 408022 516934
rect 407786 481018 408022 481254
rect 407786 480698 408022 480934
rect 407786 445018 408022 445254
rect 407786 444698 408022 444934
rect 407786 409018 408022 409254
rect 407786 408698 408022 408934
rect 407786 373018 408022 373254
rect 407786 372698 408022 372934
rect 407786 337018 408022 337254
rect 407786 336698 408022 336934
rect 407786 301018 408022 301254
rect 407786 300698 408022 300934
rect 407786 265018 408022 265254
rect 407786 264698 408022 264934
rect 407786 229018 408022 229254
rect 407786 228698 408022 228934
rect 407786 193018 408022 193254
rect 407786 192698 408022 192934
rect 407786 157018 408022 157254
rect 407786 156698 408022 156934
rect 407786 121018 408022 121254
rect 407786 120698 408022 120934
rect 407786 85018 408022 85254
rect 407786 84698 408022 84934
rect 407786 49018 408022 49254
rect 407786 48698 408022 48934
rect 407786 13018 408022 13254
rect 407786 12698 408022 12934
rect 389786 -7162 390022 -6926
rect 389786 -7482 390022 -7246
rect 414986 705542 415222 705778
rect 414986 705222 415222 705458
rect 414986 668218 415222 668454
rect 414986 667898 415222 668134
rect 414986 632218 415222 632454
rect 414986 631898 415222 632134
rect 414986 596218 415222 596454
rect 414986 595898 415222 596134
rect 414986 560218 415222 560454
rect 414986 559898 415222 560134
rect 414986 524218 415222 524454
rect 414986 523898 415222 524134
rect 414986 488218 415222 488454
rect 414986 487898 415222 488134
rect 414986 452218 415222 452454
rect 414986 451898 415222 452134
rect 414986 416218 415222 416454
rect 414986 415898 415222 416134
rect 414986 380218 415222 380454
rect 414986 379898 415222 380134
rect 414986 344218 415222 344454
rect 414986 343898 415222 344134
rect 414986 308218 415222 308454
rect 414986 307898 415222 308134
rect 414986 272218 415222 272454
rect 414986 271898 415222 272134
rect 414986 236218 415222 236454
rect 414986 235898 415222 236134
rect 414986 200218 415222 200454
rect 414986 199898 415222 200134
rect 414986 164218 415222 164454
rect 414986 163898 415222 164134
rect 414986 128218 415222 128454
rect 414986 127898 415222 128134
rect 414986 92218 415222 92454
rect 414986 91898 415222 92134
rect 414986 56218 415222 56454
rect 414986 55898 415222 56134
rect 414986 20218 415222 20454
rect 414986 19898 415222 20134
rect 414986 -1522 415222 -1286
rect 414986 -1842 415222 -1606
rect 418586 671818 418822 672054
rect 418586 671498 418822 671734
rect 418586 635818 418822 636054
rect 418586 635498 418822 635734
rect 418586 599818 418822 600054
rect 418586 599498 418822 599734
rect 418586 563818 418822 564054
rect 418586 563498 418822 563734
rect 418586 527818 418822 528054
rect 418586 527498 418822 527734
rect 418586 491818 418822 492054
rect 418586 491498 418822 491734
rect 418586 455818 418822 456054
rect 418586 455498 418822 455734
rect 418586 419818 418822 420054
rect 418586 419498 418822 419734
rect 418586 383818 418822 384054
rect 418586 383498 418822 383734
rect 418586 347818 418822 348054
rect 418586 347498 418822 347734
rect 418586 311818 418822 312054
rect 418586 311498 418822 311734
rect 418586 275818 418822 276054
rect 418586 275498 418822 275734
rect 418586 239818 418822 240054
rect 418586 239498 418822 239734
rect 418586 203818 418822 204054
rect 418586 203498 418822 203734
rect 418586 167818 418822 168054
rect 418586 167498 418822 167734
rect 418586 131818 418822 132054
rect 418586 131498 418822 131734
rect 418586 95818 418822 96054
rect 418586 95498 418822 95734
rect 422186 675418 422422 675654
rect 422186 675098 422422 675334
rect 422186 639418 422422 639654
rect 422186 639098 422422 639334
rect 422186 603418 422422 603654
rect 422186 603098 422422 603334
rect 422186 567418 422422 567654
rect 422186 567098 422422 567334
rect 422186 531418 422422 531654
rect 422186 531098 422422 531334
rect 422186 495418 422422 495654
rect 422186 495098 422422 495334
rect 422186 459418 422422 459654
rect 422186 459098 422422 459334
rect 422186 423418 422422 423654
rect 422186 423098 422422 423334
rect 422186 387418 422422 387654
rect 422186 387098 422422 387334
rect 422186 351418 422422 351654
rect 422186 351098 422422 351334
rect 422186 315418 422422 315654
rect 422186 315098 422422 315334
rect 422186 279418 422422 279654
rect 422186 279098 422422 279334
rect 422186 243418 422422 243654
rect 422186 243098 422422 243334
rect 422186 207418 422422 207654
rect 422186 207098 422422 207334
rect 422186 171418 422422 171654
rect 422186 171098 422422 171334
rect 422186 135418 422422 135654
rect 422186 135098 422422 135334
rect 422186 99418 422422 99654
rect 422186 99098 422422 99334
rect 422186 63418 422422 63654
rect 422186 63098 422422 63334
rect 418586 59818 418822 60054
rect 418586 59498 418822 59734
rect 418586 23818 418822 24054
rect 418586 23498 418822 23734
rect 418586 -3402 418822 -3166
rect 418586 -3722 418822 -3486
rect 422186 27418 422422 27654
rect 422186 27098 422422 27334
rect 422186 -5282 422422 -5046
rect 422186 -5602 422422 -5366
rect 443786 710242 444022 710478
rect 443786 709922 444022 710158
rect 440186 708362 440422 708598
rect 440186 708042 440422 708278
rect 436586 706482 436822 706718
rect 436586 706162 436822 706398
rect 425786 679018 426022 679254
rect 425786 678698 426022 678934
rect 425786 643018 426022 643254
rect 425786 642698 426022 642934
rect 425786 607018 426022 607254
rect 425786 606698 426022 606934
rect 425786 571018 426022 571254
rect 425786 570698 426022 570934
rect 425786 535018 426022 535254
rect 425786 534698 426022 534934
rect 425786 499018 426022 499254
rect 425786 498698 426022 498934
rect 425786 463018 426022 463254
rect 425786 462698 426022 462934
rect 425786 427018 426022 427254
rect 425786 426698 426022 426934
rect 425786 391018 426022 391254
rect 425786 390698 426022 390934
rect 425786 355018 426022 355254
rect 425786 354698 426022 354934
rect 425786 319018 426022 319254
rect 425786 318698 426022 318934
rect 425786 283018 426022 283254
rect 425786 282698 426022 282934
rect 425786 247018 426022 247254
rect 425786 246698 426022 246934
rect 425786 211018 426022 211254
rect 425786 210698 426022 210934
rect 425786 175018 426022 175254
rect 425786 174698 426022 174934
rect 425786 139018 426022 139254
rect 425786 138698 426022 138934
rect 425786 103018 426022 103254
rect 425786 102698 426022 102934
rect 425786 67018 426022 67254
rect 425786 66698 426022 66934
rect 425786 31018 426022 31254
rect 425786 30698 426022 30934
rect 407786 -6222 408022 -5986
rect 407786 -6542 408022 -6306
rect 432986 704602 433222 704838
rect 432986 704282 433222 704518
rect 432986 686218 433222 686454
rect 432986 685898 433222 686134
rect 432986 650218 433222 650454
rect 432986 649898 433222 650134
rect 432986 614218 433222 614454
rect 432986 613898 433222 614134
rect 432986 578218 433222 578454
rect 432986 577898 433222 578134
rect 432986 542218 433222 542454
rect 432986 541898 433222 542134
rect 432986 506218 433222 506454
rect 432986 505898 433222 506134
rect 432986 470218 433222 470454
rect 432986 469898 433222 470134
rect 432986 434218 433222 434454
rect 432986 433898 433222 434134
rect 432986 398218 433222 398454
rect 432986 397898 433222 398134
rect 432986 362218 433222 362454
rect 432986 361898 433222 362134
rect 432986 326218 433222 326454
rect 432986 325898 433222 326134
rect 432986 290218 433222 290454
rect 432986 289898 433222 290134
rect 432986 254218 433222 254454
rect 432986 253898 433222 254134
rect 432986 218218 433222 218454
rect 432986 217898 433222 218134
rect 432986 182218 433222 182454
rect 432986 181898 433222 182134
rect 432986 146218 433222 146454
rect 432986 145898 433222 146134
rect 432986 110218 433222 110454
rect 432986 109898 433222 110134
rect 432986 74218 433222 74454
rect 432986 73898 433222 74134
rect 432986 38218 433222 38454
rect 432986 37898 433222 38134
rect 432986 2218 433222 2454
rect 432986 1898 433222 2134
rect 432986 -582 433222 -346
rect 432986 -902 433222 -666
rect 436586 689818 436822 690054
rect 436586 689498 436822 689734
rect 436586 653818 436822 654054
rect 436586 653498 436822 653734
rect 436586 617818 436822 618054
rect 436586 617498 436822 617734
rect 436586 581818 436822 582054
rect 436586 581498 436822 581734
rect 436586 545818 436822 546054
rect 436586 545498 436822 545734
rect 436586 509818 436822 510054
rect 436586 509498 436822 509734
rect 436586 473818 436822 474054
rect 436586 473498 436822 473734
rect 436586 437818 436822 438054
rect 436586 437498 436822 437734
rect 436586 401818 436822 402054
rect 436586 401498 436822 401734
rect 436586 365818 436822 366054
rect 436586 365498 436822 365734
rect 436586 329818 436822 330054
rect 436586 329498 436822 329734
rect 436586 293818 436822 294054
rect 436586 293498 436822 293734
rect 436586 257818 436822 258054
rect 436586 257498 436822 257734
rect 436586 221818 436822 222054
rect 436586 221498 436822 221734
rect 436586 185818 436822 186054
rect 436586 185498 436822 185734
rect 436586 149818 436822 150054
rect 436586 149498 436822 149734
rect 436586 113818 436822 114054
rect 436586 113498 436822 113734
rect 436586 77818 436822 78054
rect 436586 77498 436822 77734
rect 436586 41818 436822 42054
rect 436586 41498 436822 41734
rect 436586 5818 436822 6054
rect 436586 5498 436822 5734
rect 436586 -2462 436822 -2226
rect 436586 -2782 436822 -2546
rect 440186 693418 440422 693654
rect 440186 693098 440422 693334
rect 440186 657418 440422 657654
rect 440186 657098 440422 657334
rect 440186 621418 440422 621654
rect 440186 621098 440422 621334
rect 440186 585418 440422 585654
rect 440186 585098 440422 585334
rect 440186 549418 440422 549654
rect 440186 549098 440422 549334
rect 440186 513418 440422 513654
rect 440186 513098 440422 513334
rect 440186 477418 440422 477654
rect 440186 477098 440422 477334
rect 440186 441418 440422 441654
rect 440186 441098 440422 441334
rect 440186 405418 440422 405654
rect 440186 405098 440422 405334
rect 440186 369418 440422 369654
rect 440186 369098 440422 369334
rect 440186 333418 440422 333654
rect 440186 333098 440422 333334
rect 440186 297418 440422 297654
rect 440186 297098 440422 297334
rect 440186 261418 440422 261654
rect 440186 261098 440422 261334
rect 440186 225418 440422 225654
rect 440186 225098 440422 225334
rect 440186 189418 440422 189654
rect 440186 189098 440422 189334
rect 440186 153418 440422 153654
rect 440186 153098 440422 153334
rect 440186 117418 440422 117654
rect 440186 117098 440422 117334
rect 440186 81418 440422 81654
rect 440186 81098 440422 81334
rect 440186 45418 440422 45654
rect 440186 45098 440422 45334
rect 440186 9418 440422 9654
rect 440186 9098 440422 9334
rect 440186 -4342 440422 -4106
rect 440186 -4662 440422 -4426
rect 461786 711182 462022 711418
rect 461786 710862 462022 711098
rect 458186 709302 458422 709538
rect 458186 708982 458422 709218
rect 454586 707422 454822 707658
rect 454586 707102 454822 707338
rect 443786 697018 444022 697254
rect 443786 696698 444022 696934
rect 443786 661018 444022 661254
rect 443786 660698 444022 660934
rect 443786 625018 444022 625254
rect 443786 624698 444022 624934
rect 443786 589018 444022 589254
rect 443786 588698 444022 588934
rect 443786 553018 444022 553254
rect 443786 552698 444022 552934
rect 443786 517018 444022 517254
rect 443786 516698 444022 516934
rect 443786 481018 444022 481254
rect 443786 480698 444022 480934
rect 443786 445018 444022 445254
rect 443786 444698 444022 444934
rect 443786 409018 444022 409254
rect 443786 408698 444022 408934
rect 443786 373018 444022 373254
rect 443786 372698 444022 372934
rect 443786 337018 444022 337254
rect 443786 336698 444022 336934
rect 443786 301018 444022 301254
rect 443786 300698 444022 300934
rect 443786 265018 444022 265254
rect 443786 264698 444022 264934
rect 443786 229018 444022 229254
rect 443786 228698 444022 228934
rect 443786 193018 444022 193254
rect 443786 192698 444022 192934
rect 443786 157018 444022 157254
rect 443786 156698 444022 156934
rect 443786 121018 444022 121254
rect 443786 120698 444022 120934
rect 443786 85018 444022 85254
rect 443786 84698 444022 84934
rect 443786 49018 444022 49254
rect 443786 48698 444022 48934
rect 443786 13018 444022 13254
rect 443786 12698 444022 12934
rect 425786 -7162 426022 -6926
rect 425786 -7482 426022 -7246
rect 450986 705542 451222 705778
rect 450986 705222 451222 705458
rect 450986 668218 451222 668454
rect 450986 667898 451222 668134
rect 450986 632218 451222 632454
rect 450986 631898 451222 632134
rect 450986 596218 451222 596454
rect 450986 595898 451222 596134
rect 450986 560218 451222 560454
rect 450986 559898 451222 560134
rect 450986 524218 451222 524454
rect 450986 523898 451222 524134
rect 450986 488218 451222 488454
rect 450986 487898 451222 488134
rect 450986 452218 451222 452454
rect 450986 451898 451222 452134
rect 450986 416218 451222 416454
rect 450986 415898 451222 416134
rect 450986 380218 451222 380454
rect 450986 379898 451222 380134
rect 450986 344218 451222 344454
rect 450986 343898 451222 344134
rect 450986 308218 451222 308454
rect 450986 307898 451222 308134
rect 450986 272218 451222 272454
rect 450986 271898 451222 272134
rect 450986 236218 451222 236454
rect 450986 235898 451222 236134
rect 450986 200218 451222 200454
rect 450986 199898 451222 200134
rect 450986 164218 451222 164454
rect 450986 163898 451222 164134
rect 450986 128218 451222 128454
rect 450986 127898 451222 128134
rect 450986 92218 451222 92454
rect 450986 91898 451222 92134
rect 450986 56218 451222 56454
rect 450986 55898 451222 56134
rect 450986 20218 451222 20454
rect 450986 19898 451222 20134
rect 450986 -1522 451222 -1286
rect 450986 -1842 451222 -1606
rect 454586 671818 454822 672054
rect 454586 671498 454822 671734
rect 454586 635818 454822 636054
rect 454586 635498 454822 635734
rect 454586 599818 454822 600054
rect 454586 599498 454822 599734
rect 454586 563818 454822 564054
rect 454586 563498 454822 563734
rect 454586 527818 454822 528054
rect 454586 527498 454822 527734
rect 454586 491818 454822 492054
rect 454586 491498 454822 491734
rect 454586 455818 454822 456054
rect 454586 455498 454822 455734
rect 454586 419818 454822 420054
rect 454586 419498 454822 419734
rect 454586 383818 454822 384054
rect 454586 383498 454822 383734
rect 454586 347818 454822 348054
rect 454586 347498 454822 347734
rect 454586 311818 454822 312054
rect 454586 311498 454822 311734
rect 454586 275818 454822 276054
rect 454586 275498 454822 275734
rect 454586 239818 454822 240054
rect 454586 239498 454822 239734
rect 454586 203818 454822 204054
rect 454586 203498 454822 203734
rect 454586 167818 454822 168054
rect 454586 167498 454822 167734
rect 454586 131818 454822 132054
rect 454586 131498 454822 131734
rect 454586 95818 454822 96054
rect 454586 95498 454822 95734
rect 454586 59818 454822 60054
rect 454586 59498 454822 59734
rect 454586 23818 454822 24054
rect 454586 23498 454822 23734
rect 454586 -3402 454822 -3166
rect 454586 -3722 454822 -3486
rect 458186 675418 458422 675654
rect 458186 675098 458422 675334
rect 458186 639418 458422 639654
rect 458186 639098 458422 639334
rect 458186 603418 458422 603654
rect 458186 603098 458422 603334
rect 458186 567418 458422 567654
rect 458186 567098 458422 567334
rect 458186 531418 458422 531654
rect 458186 531098 458422 531334
rect 458186 495418 458422 495654
rect 458186 495098 458422 495334
rect 458186 459418 458422 459654
rect 458186 459098 458422 459334
rect 458186 423418 458422 423654
rect 458186 423098 458422 423334
rect 458186 387418 458422 387654
rect 458186 387098 458422 387334
rect 458186 351418 458422 351654
rect 458186 351098 458422 351334
rect 458186 315418 458422 315654
rect 458186 315098 458422 315334
rect 458186 279418 458422 279654
rect 458186 279098 458422 279334
rect 458186 243418 458422 243654
rect 458186 243098 458422 243334
rect 458186 207418 458422 207654
rect 458186 207098 458422 207334
rect 458186 171418 458422 171654
rect 458186 171098 458422 171334
rect 458186 135418 458422 135654
rect 458186 135098 458422 135334
rect 458186 99418 458422 99654
rect 458186 99098 458422 99334
rect 458186 63418 458422 63654
rect 458186 63098 458422 63334
rect 458186 27418 458422 27654
rect 458186 27098 458422 27334
rect 458186 -5282 458422 -5046
rect 458186 -5602 458422 -5366
rect 479786 710242 480022 710478
rect 479786 709922 480022 710158
rect 476186 708362 476422 708598
rect 476186 708042 476422 708278
rect 472586 706482 472822 706718
rect 472586 706162 472822 706398
rect 461786 679018 462022 679254
rect 461786 678698 462022 678934
rect 461786 643018 462022 643254
rect 461786 642698 462022 642934
rect 461786 607018 462022 607254
rect 461786 606698 462022 606934
rect 461786 571018 462022 571254
rect 461786 570698 462022 570934
rect 461786 535018 462022 535254
rect 461786 534698 462022 534934
rect 461786 499018 462022 499254
rect 461786 498698 462022 498934
rect 461786 463018 462022 463254
rect 461786 462698 462022 462934
rect 461786 427018 462022 427254
rect 461786 426698 462022 426934
rect 461786 391018 462022 391254
rect 461786 390698 462022 390934
rect 461786 355018 462022 355254
rect 461786 354698 462022 354934
rect 461786 319018 462022 319254
rect 461786 318698 462022 318934
rect 461786 283018 462022 283254
rect 461786 282698 462022 282934
rect 461786 247018 462022 247254
rect 461786 246698 462022 246934
rect 461786 211018 462022 211254
rect 461786 210698 462022 210934
rect 461786 175018 462022 175254
rect 461786 174698 462022 174934
rect 461786 139018 462022 139254
rect 461786 138698 462022 138934
rect 461786 103018 462022 103254
rect 461786 102698 462022 102934
rect 461786 67018 462022 67254
rect 461786 66698 462022 66934
rect 461786 31018 462022 31254
rect 461786 30698 462022 30934
rect 443786 -6222 444022 -5986
rect 443786 -6542 444022 -6306
rect 468986 704602 469222 704838
rect 468986 704282 469222 704518
rect 468986 686218 469222 686454
rect 468986 685898 469222 686134
rect 468986 650218 469222 650454
rect 468986 649898 469222 650134
rect 468986 614218 469222 614454
rect 468986 613898 469222 614134
rect 468986 578218 469222 578454
rect 468986 577898 469222 578134
rect 468986 542218 469222 542454
rect 468986 541898 469222 542134
rect 468986 506218 469222 506454
rect 468986 505898 469222 506134
rect 468986 470218 469222 470454
rect 468986 469898 469222 470134
rect 468986 434218 469222 434454
rect 468986 433898 469222 434134
rect 468986 398218 469222 398454
rect 468986 397898 469222 398134
rect 468986 362218 469222 362454
rect 468986 361898 469222 362134
rect 468986 326218 469222 326454
rect 468986 325898 469222 326134
rect 468986 290218 469222 290454
rect 468986 289898 469222 290134
rect 468986 254218 469222 254454
rect 468986 253898 469222 254134
rect 468986 218218 469222 218454
rect 468986 217898 469222 218134
rect 468986 182218 469222 182454
rect 468986 181898 469222 182134
rect 468986 146218 469222 146454
rect 468986 145898 469222 146134
rect 468986 110218 469222 110454
rect 468986 109898 469222 110134
rect 468986 74218 469222 74454
rect 468986 73898 469222 74134
rect 468986 38218 469222 38454
rect 468986 37898 469222 38134
rect 468986 2218 469222 2454
rect 468986 1898 469222 2134
rect 468986 -582 469222 -346
rect 468986 -902 469222 -666
rect 472586 689818 472822 690054
rect 472586 689498 472822 689734
rect 472586 653818 472822 654054
rect 472586 653498 472822 653734
rect 472586 617818 472822 618054
rect 472586 617498 472822 617734
rect 472586 581818 472822 582054
rect 472586 581498 472822 581734
rect 472586 545818 472822 546054
rect 472586 545498 472822 545734
rect 472586 509818 472822 510054
rect 472586 509498 472822 509734
rect 472586 473818 472822 474054
rect 472586 473498 472822 473734
rect 472586 437818 472822 438054
rect 472586 437498 472822 437734
rect 472586 401818 472822 402054
rect 472586 401498 472822 401734
rect 472586 365818 472822 366054
rect 472586 365498 472822 365734
rect 472586 329818 472822 330054
rect 472586 329498 472822 329734
rect 472586 293818 472822 294054
rect 472586 293498 472822 293734
rect 472586 257818 472822 258054
rect 472586 257498 472822 257734
rect 472586 221818 472822 222054
rect 472586 221498 472822 221734
rect 472586 185818 472822 186054
rect 472586 185498 472822 185734
rect 472586 149818 472822 150054
rect 472586 149498 472822 149734
rect 472586 113818 472822 114054
rect 472586 113498 472822 113734
rect 472586 77818 472822 78054
rect 472586 77498 472822 77734
rect 472586 41818 472822 42054
rect 472586 41498 472822 41734
rect 472586 5818 472822 6054
rect 472586 5498 472822 5734
rect 472586 -2462 472822 -2226
rect 472586 -2782 472822 -2546
rect 476186 693418 476422 693654
rect 476186 693098 476422 693334
rect 476186 657418 476422 657654
rect 476186 657098 476422 657334
rect 476186 621418 476422 621654
rect 476186 621098 476422 621334
rect 476186 585418 476422 585654
rect 476186 585098 476422 585334
rect 476186 549418 476422 549654
rect 476186 549098 476422 549334
rect 476186 513418 476422 513654
rect 476186 513098 476422 513334
rect 476186 477418 476422 477654
rect 476186 477098 476422 477334
rect 476186 441418 476422 441654
rect 476186 441098 476422 441334
rect 476186 405418 476422 405654
rect 476186 405098 476422 405334
rect 476186 369418 476422 369654
rect 476186 369098 476422 369334
rect 476186 333418 476422 333654
rect 476186 333098 476422 333334
rect 476186 297418 476422 297654
rect 476186 297098 476422 297334
rect 476186 261418 476422 261654
rect 476186 261098 476422 261334
rect 476186 225418 476422 225654
rect 476186 225098 476422 225334
rect 476186 189418 476422 189654
rect 476186 189098 476422 189334
rect 476186 153418 476422 153654
rect 476186 153098 476422 153334
rect 476186 117418 476422 117654
rect 476186 117098 476422 117334
rect 476186 81418 476422 81654
rect 476186 81098 476422 81334
rect 476186 45418 476422 45654
rect 476186 45098 476422 45334
rect 476186 9418 476422 9654
rect 476186 9098 476422 9334
rect 476186 -4342 476422 -4106
rect 476186 -4662 476422 -4426
rect 497786 711182 498022 711418
rect 497786 710862 498022 711098
rect 494186 709302 494422 709538
rect 494186 708982 494422 709218
rect 490586 707422 490822 707658
rect 490586 707102 490822 707338
rect 479786 697018 480022 697254
rect 479786 696698 480022 696934
rect 479786 661018 480022 661254
rect 479786 660698 480022 660934
rect 479786 625018 480022 625254
rect 479786 624698 480022 624934
rect 479786 589018 480022 589254
rect 479786 588698 480022 588934
rect 479786 553018 480022 553254
rect 479786 552698 480022 552934
rect 479786 517018 480022 517254
rect 479786 516698 480022 516934
rect 479786 481018 480022 481254
rect 479786 480698 480022 480934
rect 479786 445018 480022 445254
rect 479786 444698 480022 444934
rect 479786 409018 480022 409254
rect 479786 408698 480022 408934
rect 479786 373018 480022 373254
rect 479786 372698 480022 372934
rect 479786 337018 480022 337254
rect 479786 336698 480022 336934
rect 479786 301018 480022 301254
rect 479786 300698 480022 300934
rect 479786 265018 480022 265254
rect 479786 264698 480022 264934
rect 479786 229018 480022 229254
rect 479786 228698 480022 228934
rect 479786 193018 480022 193254
rect 479786 192698 480022 192934
rect 479786 157018 480022 157254
rect 479786 156698 480022 156934
rect 479786 121018 480022 121254
rect 479786 120698 480022 120934
rect 479786 85018 480022 85254
rect 479786 84698 480022 84934
rect 479786 49018 480022 49254
rect 479786 48698 480022 48934
rect 479786 13018 480022 13254
rect 479786 12698 480022 12934
rect 461786 -7162 462022 -6926
rect 461786 -7482 462022 -7246
rect 486986 705542 487222 705778
rect 486986 705222 487222 705458
rect 486986 668218 487222 668454
rect 486986 667898 487222 668134
rect 486986 632218 487222 632454
rect 486986 631898 487222 632134
rect 486986 596218 487222 596454
rect 486986 595898 487222 596134
rect 486986 560218 487222 560454
rect 486986 559898 487222 560134
rect 486986 524218 487222 524454
rect 486986 523898 487222 524134
rect 486986 488218 487222 488454
rect 486986 487898 487222 488134
rect 486986 452218 487222 452454
rect 486986 451898 487222 452134
rect 486986 416218 487222 416454
rect 486986 415898 487222 416134
rect 486986 380218 487222 380454
rect 486986 379898 487222 380134
rect 486986 344218 487222 344454
rect 486986 343898 487222 344134
rect 486986 308218 487222 308454
rect 486986 307898 487222 308134
rect 486986 272218 487222 272454
rect 486986 271898 487222 272134
rect 486986 236218 487222 236454
rect 486986 235898 487222 236134
rect 486986 200218 487222 200454
rect 486986 199898 487222 200134
rect 486986 164218 487222 164454
rect 486986 163898 487222 164134
rect 486986 128218 487222 128454
rect 486986 127898 487222 128134
rect 486986 92218 487222 92454
rect 486986 91898 487222 92134
rect 486986 56218 487222 56454
rect 486986 55898 487222 56134
rect 486986 20218 487222 20454
rect 486986 19898 487222 20134
rect 486986 -1522 487222 -1286
rect 486986 -1842 487222 -1606
rect 490586 671818 490822 672054
rect 490586 671498 490822 671734
rect 490586 635818 490822 636054
rect 490586 635498 490822 635734
rect 490586 599818 490822 600054
rect 490586 599498 490822 599734
rect 490586 563818 490822 564054
rect 490586 563498 490822 563734
rect 490586 527818 490822 528054
rect 490586 527498 490822 527734
rect 490586 491818 490822 492054
rect 490586 491498 490822 491734
rect 490586 455818 490822 456054
rect 490586 455498 490822 455734
rect 490586 419818 490822 420054
rect 490586 419498 490822 419734
rect 490586 383818 490822 384054
rect 490586 383498 490822 383734
rect 490586 347818 490822 348054
rect 490586 347498 490822 347734
rect 490586 311818 490822 312054
rect 490586 311498 490822 311734
rect 490586 275818 490822 276054
rect 490586 275498 490822 275734
rect 490586 239818 490822 240054
rect 490586 239498 490822 239734
rect 490586 203818 490822 204054
rect 490586 203498 490822 203734
rect 490586 167818 490822 168054
rect 490586 167498 490822 167734
rect 490586 131818 490822 132054
rect 490586 131498 490822 131734
rect 490586 95818 490822 96054
rect 490586 95498 490822 95734
rect 490586 59818 490822 60054
rect 490586 59498 490822 59734
rect 490586 23818 490822 24054
rect 490586 23498 490822 23734
rect 490586 -3402 490822 -3166
rect 490586 -3722 490822 -3486
rect 494186 675418 494422 675654
rect 494186 675098 494422 675334
rect 494186 639418 494422 639654
rect 494186 639098 494422 639334
rect 494186 603418 494422 603654
rect 494186 603098 494422 603334
rect 494186 567418 494422 567654
rect 494186 567098 494422 567334
rect 494186 531418 494422 531654
rect 494186 531098 494422 531334
rect 494186 495418 494422 495654
rect 494186 495098 494422 495334
rect 494186 459418 494422 459654
rect 494186 459098 494422 459334
rect 494186 423418 494422 423654
rect 494186 423098 494422 423334
rect 494186 387418 494422 387654
rect 494186 387098 494422 387334
rect 494186 351418 494422 351654
rect 494186 351098 494422 351334
rect 494186 315418 494422 315654
rect 494186 315098 494422 315334
rect 494186 279418 494422 279654
rect 494186 279098 494422 279334
rect 494186 243418 494422 243654
rect 494186 243098 494422 243334
rect 494186 207418 494422 207654
rect 494186 207098 494422 207334
rect 494186 171418 494422 171654
rect 494186 171098 494422 171334
rect 494186 135418 494422 135654
rect 494186 135098 494422 135334
rect 494186 99418 494422 99654
rect 494186 99098 494422 99334
rect 494186 63418 494422 63654
rect 494186 63098 494422 63334
rect 494186 27418 494422 27654
rect 494186 27098 494422 27334
rect 494186 -5282 494422 -5046
rect 494186 -5602 494422 -5366
rect 515786 710242 516022 710478
rect 515786 709922 516022 710158
rect 512186 708362 512422 708598
rect 512186 708042 512422 708278
rect 508586 706482 508822 706718
rect 508586 706162 508822 706398
rect 497786 679018 498022 679254
rect 497786 678698 498022 678934
rect 497786 643018 498022 643254
rect 497786 642698 498022 642934
rect 497786 607018 498022 607254
rect 497786 606698 498022 606934
rect 497786 571018 498022 571254
rect 497786 570698 498022 570934
rect 497786 535018 498022 535254
rect 497786 534698 498022 534934
rect 497786 499018 498022 499254
rect 497786 498698 498022 498934
rect 497786 463018 498022 463254
rect 497786 462698 498022 462934
rect 497786 427018 498022 427254
rect 497786 426698 498022 426934
rect 497786 391018 498022 391254
rect 497786 390698 498022 390934
rect 497786 355018 498022 355254
rect 497786 354698 498022 354934
rect 497786 319018 498022 319254
rect 497786 318698 498022 318934
rect 497786 283018 498022 283254
rect 497786 282698 498022 282934
rect 497786 247018 498022 247254
rect 497786 246698 498022 246934
rect 497786 211018 498022 211254
rect 497786 210698 498022 210934
rect 497786 175018 498022 175254
rect 497786 174698 498022 174934
rect 497786 139018 498022 139254
rect 497786 138698 498022 138934
rect 497786 103018 498022 103254
rect 497786 102698 498022 102934
rect 497786 67018 498022 67254
rect 497786 66698 498022 66934
rect 497786 31018 498022 31254
rect 497786 30698 498022 30934
rect 479786 -6222 480022 -5986
rect 479786 -6542 480022 -6306
rect 504986 704602 505222 704838
rect 504986 704282 505222 704518
rect 504986 686218 505222 686454
rect 504986 685898 505222 686134
rect 504986 650218 505222 650454
rect 504986 649898 505222 650134
rect 504986 614218 505222 614454
rect 504986 613898 505222 614134
rect 504986 578218 505222 578454
rect 504986 577898 505222 578134
rect 504986 542218 505222 542454
rect 504986 541898 505222 542134
rect 504986 506218 505222 506454
rect 504986 505898 505222 506134
rect 504986 470218 505222 470454
rect 504986 469898 505222 470134
rect 504986 434218 505222 434454
rect 504986 433898 505222 434134
rect 504986 398218 505222 398454
rect 504986 397898 505222 398134
rect 504986 362218 505222 362454
rect 504986 361898 505222 362134
rect 504986 326218 505222 326454
rect 504986 325898 505222 326134
rect 504986 290218 505222 290454
rect 504986 289898 505222 290134
rect 504986 254218 505222 254454
rect 504986 253898 505222 254134
rect 504986 218218 505222 218454
rect 504986 217898 505222 218134
rect 504986 182218 505222 182454
rect 504986 181898 505222 182134
rect 504986 146218 505222 146454
rect 504986 145898 505222 146134
rect 504986 110218 505222 110454
rect 504986 109898 505222 110134
rect 504986 74218 505222 74454
rect 504986 73898 505222 74134
rect 504986 38218 505222 38454
rect 504986 37898 505222 38134
rect 504986 2218 505222 2454
rect 504986 1898 505222 2134
rect 504986 -582 505222 -346
rect 504986 -902 505222 -666
rect 508586 689818 508822 690054
rect 508586 689498 508822 689734
rect 508586 653818 508822 654054
rect 508586 653498 508822 653734
rect 508586 617818 508822 618054
rect 508586 617498 508822 617734
rect 508586 581818 508822 582054
rect 508586 581498 508822 581734
rect 508586 545818 508822 546054
rect 508586 545498 508822 545734
rect 508586 509818 508822 510054
rect 508586 509498 508822 509734
rect 508586 473818 508822 474054
rect 508586 473498 508822 473734
rect 508586 437818 508822 438054
rect 508586 437498 508822 437734
rect 508586 401818 508822 402054
rect 508586 401498 508822 401734
rect 508586 365818 508822 366054
rect 508586 365498 508822 365734
rect 508586 329818 508822 330054
rect 508586 329498 508822 329734
rect 508586 293818 508822 294054
rect 508586 293498 508822 293734
rect 508586 257818 508822 258054
rect 508586 257498 508822 257734
rect 508586 221818 508822 222054
rect 508586 221498 508822 221734
rect 508586 185818 508822 186054
rect 508586 185498 508822 185734
rect 508586 149818 508822 150054
rect 508586 149498 508822 149734
rect 508586 113818 508822 114054
rect 508586 113498 508822 113734
rect 508586 77818 508822 78054
rect 508586 77498 508822 77734
rect 508586 41818 508822 42054
rect 508586 41498 508822 41734
rect 508586 5818 508822 6054
rect 508586 5498 508822 5734
rect 508586 -2462 508822 -2226
rect 508586 -2782 508822 -2546
rect 512186 693418 512422 693654
rect 512186 693098 512422 693334
rect 512186 657418 512422 657654
rect 512186 657098 512422 657334
rect 512186 621418 512422 621654
rect 512186 621098 512422 621334
rect 512186 585418 512422 585654
rect 512186 585098 512422 585334
rect 512186 549418 512422 549654
rect 512186 549098 512422 549334
rect 512186 513418 512422 513654
rect 512186 513098 512422 513334
rect 512186 477418 512422 477654
rect 512186 477098 512422 477334
rect 512186 441418 512422 441654
rect 512186 441098 512422 441334
rect 512186 405418 512422 405654
rect 512186 405098 512422 405334
rect 512186 369418 512422 369654
rect 512186 369098 512422 369334
rect 512186 333418 512422 333654
rect 512186 333098 512422 333334
rect 512186 297418 512422 297654
rect 512186 297098 512422 297334
rect 512186 261418 512422 261654
rect 512186 261098 512422 261334
rect 512186 225418 512422 225654
rect 512186 225098 512422 225334
rect 512186 189418 512422 189654
rect 512186 189098 512422 189334
rect 512186 153418 512422 153654
rect 512186 153098 512422 153334
rect 512186 117418 512422 117654
rect 512186 117098 512422 117334
rect 512186 81418 512422 81654
rect 512186 81098 512422 81334
rect 512186 45418 512422 45654
rect 512186 45098 512422 45334
rect 512186 9418 512422 9654
rect 512186 9098 512422 9334
rect 512186 -4342 512422 -4106
rect 512186 -4662 512422 -4426
rect 533786 711182 534022 711418
rect 533786 710862 534022 711098
rect 530186 709302 530422 709538
rect 530186 708982 530422 709218
rect 526586 707422 526822 707658
rect 526586 707102 526822 707338
rect 515786 697018 516022 697254
rect 515786 696698 516022 696934
rect 515786 661018 516022 661254
rect 515786 660698 516022 660934
rect 515786 625018 516022 625254
rect 515786 624698 516022 624934
rect 515786 589018 516022 589254
rect 515786 588698 516022 588934
rect 515786 553018 516022 553254
rect 515786 552698 516022 552934
rect 515786 517018 516022 517254
rect 515786 516698 516022 516934
rect 515786 481018 516022 481254
rect 515786 480698 516022 480934
rect 515786 445018 516022 445254
rect 515786 444698 516022 444934
rect 515786 409018 516022 409254
rect 515786 408698 516022 408934
rect 515786 373018 516022 373254
rect 515786 372698 516022 372934
rect 515786 337018 516022 337254
rect 515786 336698 516022 336934
rect 515786 301018 516022 301254
rect 515786 300698 516022 300934
rect 515786 265018 516022 265254
rect 515786 264698 516022 264934
rect 515786 229018 516022 229254
rect 515786 228698 516022 228934
rect 515786 193018 516022 193254
rect 515786 192698 516022 192934
rect 515786 157018 516022 157254
rect 515786 156698 516022 156934
rect 515786 121018 516022 121254
rect 515786 120698 516022 120934
rect 515786 85018 516022 85254
rect 515786 84698 516022 84934
rect 515786 49018 516022 49254
rect 515786 48698 516022 48934
rect 515786 13018 516022 13254
rect 515786 12698 516022 12934
rect 497786 -7162 498022 -6926
rect 497786 -7482 498022 -7246
rect 522986 705542 523222 705778
rect 522986 705222 523222 705458
rect 522986 668218 523222 668454
rect 522986 667898 523222 668134
rect 522986 632218 523222 632454
rect 522986 631898 523222 632134
rect 522986 596218 523222 596454
rect 522986 595898 523222 596134
rect 522986 560218 523222 560454
rect 522986 559898 523222 560134
rect 522986 524218 523222 524454
rect 522986 523898 523222 524134
rect 522986 488218 523222 488454
rect 522986 487898 523222 488134
rect 522986 452218 523222 452454
rect 522986 451898 523222 452134
rect 522986 416218 523222 416454
rect 522986 415898 523222 416134
rect 522986 380218 523222 380454
rect 522986 379898 523222 380134
rect 522986 344218 523222 344454
rect 522986 343898 523222 344134
rect 522986 308218 523222 308454
rect 522986 307898 523222 308134
rect 522986 272218 523222 272454
rect 522986 271898 523222 272134
rect 522986 236218 523222 236454
rect 522986 235898 523222 236134
rect 522986 200218 523222 200454
rect 522986 199898 523222 200134
rect 522986 164218 523222 164454
rect 522986 163898 523222 164134
rect 522986 128218 523222 128454
rect 522986 127898 523222 128134
rect 522986 92218 523222 92454
rect 522986 91898 523222 92134
rect 522986 56218 523222 56454
rect 522986 55898 523222 56134
rect 522986 20218 523222 20454
rect 522986 19898 523222 20134
rect 522986 -1522 523222 -1286
rect 522986 -1842 523222 -1606
rect 526586 671818 526822 672054
rect 526586 671498 526822 671734
rect 526586 635818 526822 636054
rect 526586 635498 526822 635734
rect 526586 599818 526822 600054
rect 526586 599498 526822 599734
rect 526586 563818 526822 564054
rect 526586 563498 526822 563734
rect 526586 527818 526822 528054
rect 526586 527498 526822 527734
rect 526586 491818 526822 492054
rect 526586 491498 526822 491734
rect 526586 455818 526822 456054
rect 526586 455498 526822 455734
rect 526586 419818 526822 420054
rect 526586 419498 526822 419734
rect 526586 383818 526822 384054
rect 526586 383498 526822 383734
rect 526586 347818 526822 348054
rect 526586 347498 526822 347734
rect 526586 311818 526822 312054
rect 526586 311498 526822 311734
rect 526586 275818 526822 276054
rect 526586 275498 526822 275734
rect 526586 239818 526822 240054
rect 526586 239498 526822 239734
rect 526586 203818 526822 204054
rect 526586 203498 526822 203734
rect 526586 167818 526822 168054
rect 526586 167498 526822 167734
rect 526586 131818 526822 132054
rect 526586 131498 526822 131734
rect 526586 95818 526822 96054
rect 526586 95498 526822 95734
rect 526586 59818 526822 60054
rect 526586 59498 526822 59734
rect 526586 23818 526822 24054
rect 526586 23498 526822 23734
rect 526586 -3402 526822 -3166
rect 526586 -3722 526822 -3486
rect 530186 675418 530422 675654
rect 530186 675098 530422 675334
rect 530186 639418 530422 639654
rect 530186 639098 530422 639334
rect 530186 603418 530422 603654
rect 530186 603098 530422 603334
rect 530186 567418 530422 567654
rect 530186 567098 530422 567334
rect 530186 531418 530422 531654
rect 530186 531098 530422 531334
rect 530186 495418 530422 495654
rect 530186 495098 530422 495334
rect 530186 459418 530422 459654
rect 530186 459098 530422 459334
rect 530186 423418 530422 423654
rect 530186 423098 530422 423334
rect 530186 387418 530422 387654
rect 530186 387098 530422 387334
rect 530186 351418 530422 351654
rect 530186 351098 530422 351334
rect 530186 315418 530422 315654
rect 530186 315098 530422 315334
rect 530186 279418 530422 279654
rect 530186 279098 530422 279334
rect 530186 243418 530422 243654
rect 530186 243098 530422 243334
rect 530186 207418 530422 207654
rect 530186 207098 530422 207334
rect 530186 171418 530422 171654
rect 530186 171098 530422 171334
rect 530186 135418 530422 135654
rect 530186 135098 530422 135334
rect 530186 99418 530422 99654
rect 530186 99098 530422 99334
rect 530186 63418 530422 63654
rect 530186 63098 530422 63334
rect 530186 27418 530422 27654
rect 530186 27098 530422 27334
rect 530186 -5282 530422 -5046
rect 530186 -5602 530422 -5366
rect 551786 710242 552022 710478
rect 551786 709922 552022 710158
rect 548186 708362 548422 708598
rect 548186 708042 548422 708278
rect 544586 706482 544822 706718
rect 544586 706162 544822 706398
rect 533786 679018 534022 679254
rect 533786 678698 534022 678934
rect 533786 643018 534022 643254
rect 533786 642698 534022 642934
rect 533786 607018 534022 607254
rect 533786 606698 534022 606934
rect 533786 571018 534022 571254
rect 533786 570698 534022 570934
rect 533786 535018 534022 535254
rect 533786 534698 534022 534934
rect 533786 499018 534022 499254
rect 533786 498698 534022 498934
rect 533786 463018 534022 463254
rect 533786 462698 534022 462934
rect 533786 427018 534022 427254
rect 533786 426698 534022 426934
rect 533786 391018 534022 391254
rect 533786 390698 534022 390934
rect 533786 355018 534022 355254
rect 533786 354698 534022 354934
rect 533786 319018 534022 319254
rect 533786 318698 534022 318934
rect 533786 283018 534022 283254
rect 533786 282698 534022 282934
rect 533786 247018 534022 247254
rect 533786 246698 534022 246934
rect 533786 211018 534022 211254
rect 533786 210698 534022 210934
rect 533786 175018 534022 175254
rect 533786 174698 534022 174934
rect 533786 139018 534022 139254
rect 533786 138698 534022 138934
rect 533786 103018 534022 103254
rect 533786 102698 534022 102934
rect 533786 67018 534022 67254
rect 533786 66698 534022 66934
rect 533786 31018 534022 31254
rect 533786 30698 534022 30934
rect 515786 -6222 516022 -5986
rect 515786 -6542 516022 -6306
rect 540986 704602 541222 704838
rect 540986 704282 541222 704518
rect 540986 686218 541222 686454
rect 540986 685898 541222 686134
rect 540986 650218 541222 650454
rect 540986 649898 541222 650134
rect 540986 614218 541222 614454
rect 540986 613898 541222 614134
rect 540986 578218 541222 578454
rect 540986 577898 541222 578134
rect 540986 542218 541222 542454
rect 540986 541898 541222 542134
rect 540986 506218 541222 506454
rect 540986 505898 541222 506134
rect 540986 470218 541222 470454
rect 540986 469898 541222 470134
rect 540986 434218 541222 434454
rect 540986 433898 541222 434134
rect 540986 398218 541222 398454
rect 540986 397898 541222 398134
rect 540986 362218 541222 362454
rect 540986 361898 541222 362134
rect 540986 326218 541222 326454
rect 540986 325898 541222 326134
rect 540986 290218 541222 290454
rect 540986 289898 541222 290134
rect 540986 254218 541222 254454
rect 540986 253898 541222 254134
rect 540986 218218 541222 218454
rect 540986 217898 541222 218134
rect 540986 182218 541222 182454
rect 540986 181898 541222 182134
rect 540986 146218 541222 146454
rect 540986 145898 541222 146134
rect 540986 110218 541222 110454
rect 540986 109898 541222 110134
rect 540986 74218 541222 74454
rect 540986 73898 541222 74134
rect 540986 38218 541222 38454
rect 540986 37898 541222 38134
rect 540986 2218 541222 2454
rect 540986 1898 541222 2134
rect 540986 -582 541222 -346
rect 540986 -902 541222 -666
rect 544586 689818 544822 690054
rect 544586 689498 544822 689734
rect 544586 653818 544822 654054
rect 544586 653498 544822 653734
rect 544586 617818 544822 618054
rect 544586 617498 544822 617734
rect 544586 581818 544822 582054
rect 544586 581498 544822 581734
rect 544586 545818 544822 546054
rect 544586 545498 544822 545734
rect 544586 509818 544822 510054
rect 544586 509498 544822 509734
rect 544586 473818 544822 474054
rect 544586 473498 544822 473734
rect 544586 437818 544822 438054
rect 544586 437498 544822 437734
rect 544586 401818 544822 402054
rect 544586 401498 544822 401734
rect 544586 365818 544822 366054
rect 544586 365498 544822 365734
rect 544586 329818 544822 330054
rect 544586 329498 544822 329734
rect 544586 293818 544822 294054
rect 544586 293498 544822 293734
rect 544586 257818 544822 258054
rect 544586 257498 544822 257734
rect 544586 221818 544822 222054
rect 544586 221498 544822 221734
rect 544586 185818 544822 186054
rect 544586 185498 544822 185734
rect 544586 149818 544822 150054
rect 544586 149498 544822 149734
rect 544586 113818 544822 114054
rect 544586 113498 544822 113734
rect 544586 77818 544822 78054
rect 544586 77498 544822 77734
rect 544586 41818 544822 42054
rect 544586 41498 544822 41734
rect 544586 5818 544822 6054
rect 544586 5498 544822 5734
rect 544586 -2462 544822 -2226
rect 544586 -2782 544822 -2546
rect 548186 693418 548422 693654
rect 548186 693098 548422 693334
rect 548186 657418 548422 657654
rect 548186 657098 548422 657334
rect 548186 621418 548422 621654
rect 548186 621098 548422 621334
rect 548186 585418 548422 585654
rect 548186 585098 548422 585334
rect 548186 549418 548422 549654
rect 548186 549098 548422 549334
rect 548186 513418 548422 513654
rect 548186 513098 548422 513334
rect 548186 477418 548422 477654
rect 548186 477098 548422 477334
rect 548186 441418 548422 441654
rect 548186 441098 548422 441334
rect 548186 405418 548422 405654
rect 548186 405098 548422 405334
rect 548186 369418 548422 369654
rect 548186 369098 548422 369334
rect 548186 333418 548422 333654
rect 548186 333098 548422 333334
rect 548186 297418 548422 297654
rect 548186 297098 548422 297334
rect 548186 261418 548422 261654
rect 548186 261098 548422 261334
rect 548186 225418 548422 225654
rect 548186 225098 548422 225334
rect 548186 189418 548422 189654
rect 548186 189098 548422 189334
rect 548186 153418 548422 153654
rect 548186 153098 548422 153334
rect 548186 117418 548422 117654
rect 548186 117098 548422 117334
rect 548186 81418 548422 81654
rect 548186 81098 548422 81334
rect 548186 45418 548422 45654
rect 548186 45098 548422 45334
rect 548186 9418 548422 9654
rect 548186 9098 548422 9334
rect 548186 -4342 548422 -4106
rect 548186 -4662 548422 -4426
rect 569786 711182 570022 711418
rect 569786 710862 570022 711098
rect 566186 709302 566422 709538
rect 566186 708982 566422 709218
rect 562586 707422 562822 707658
rect 562586 707102 562822 707338
rect 551786 697018 552022 697254
rect 551786 696698 552022 696934
rect 551786 661018 552022 661254
rect 551786 660698 552022 660934
rect 551786 625018 552022 625254
rect 551786 624698 552022 624934
rect 551786 589018 552022 589254
rect 551786 588698 552022 588934
rect 551786 553018 552022 553254
rect 551786 552698 552022 552934
rect 551786 517018 552022 517254
rect 551786 516698 552022 516934
rect 551786 481018 552022 481254
rect 551786 480698 552022 480934
rect 551786 445018 552022 445254
rect 551786 444698 552022 444934
rect 551786 409018 552022 409254
rect 551786 408698 552022 408934
rect 551786 373018 552022 373254
rect 551786 372698 552022 372934
rect 551786 337018 552022 337254
rect 551786 336698 552022 336934
rect 551786 301018 552022 301254
rect 551786 300698 552022 300934
rect 551786 265018 552022 265254
rect 551786 264698 552022 264934
rect 551786 229018 552022 229254
rect 551786 228698 552022 228934
rect 551786 193018 552022 193254
rect 551786 192698 552022 192934
rect 551786 157018 552022 157254
rect 551786 156698 552022 156934
rect 551786 121018 552022 121254
rect 551786 120698 552022 120934
rect 551786 85018 552022 85254
rect 551786 84698 552022 84934
rect 551786 49018 552022 49254
rect 551786 48698 552022 48934
rect 551786 13018 552022 13254
rect 551786 12698 552022 12934
rect 533786 -7162 534022 -6926
rect 533786 -7482 534022 -7246
rect 558986 705542 559222 705778
rect 558986 705222 559222 705458
rect 558986 668218 559222 668454
rect 558986 667898 559222 668134
rect 558986 632218 559222 632454
rect 558986 631898 559222 632134
rect 558986 596218 559222 596454
rect 558986 595898 559222 596134
rect 558986 560218 559222 560454
rect 558986 559898 559222 560134
rect 558986 524218 559222 524454
rect 558986 523898 559222 524134
rect 558986 488218 559222 488454
rect 558986 487898 559222 488134
rect 558986 452218 559222 452454
rect 558986 451898 559222 452134
rect 558986 416218 559222 416454
rect 558986 415898 559222 416134
rect 558986 380218 559222 380454
rect 558986 379898 559222 380134
rect 558986 344218 559222 344454
rect 558986 343898 559222 344134
rect 558986 308218 559222 308454
rect 558986 307898 559222 308134
rect 558986 272218 559222 272454
rect 558986 271898 559222 272134
rect 558986 236218 559222 236454
rect 558986 235898 559222 236134
rect 558986 200218 559222 200454
rect 558986 199898 559222 200134
rect 558986 164218 559222 164454
rect 558986 163898 559222 164134
rect 558986 128218 559222 128454
rect 558986 127898 559222 128134
rect 558986 92218 559222 92454
rect 558986 91898 559222 92134
rect 558986 56218 559222 56454
rect 558986 55898 559222 56134
rect 558986 20218 559222 20454
rect 558986 19898 559222 20134
rect 558986 -1522 559222 -1286
rect 558986 -1842 559222 -1606
rect 562586 671818 562822 672054
rect 562586 671498 562822 671734
rect 562586 635818 562822 636054
rect 562586 635498 562822 635734
rect 562586 599818 562822 600054
rect 562586 599498 562822 599734
rect 562586 563818 562822 564054
rect 562586 563498 562822 563734
rect 562586 527818 562822 528054
rect 562586 527498 562822 527734
rect 562586 491818 562822 492054
rect 562586 491498 562822 491734
rect 562586 455818 562822 456054
rect 562586 455498 562822 455734
rect 562586 419818 562822 420054
rect 562586 419498 562822 419734
rect 562586 383818 562822 384054
rect 562586 383498 562822 383734
rect 562586 347818 562822 348054
rect 562586 347498 562822 347734
rect 562586 311818 562822 312054
rect 562586 311498 562822 311734
rect 562586 275818 562822 276054
rect 562586 275498 562822 275734
rect 562586 239818 562822 240054
rect 562586 239498 562822 239734
rect 562586 203818 562822 204054
rect 562586 203498 562822 203734
rect 562586 167818 562822 168054
rect 562586 167498 562822 167734
rect 562586 131818 562822 132054
rect 562586 131498 562822 131734
rect 562586 95818 562822 96054
rect 562586 95498 562822 95734
rect 562586 59818 562822 60054
rect 562586 59498 562822 59734
rect 562586 23818 562822 24054
rect 562586 23498 562822 23734
rect 562586 -3402 562822 -3166
rect 562586 -3722 562822 -3486
rect 566186 675418 566422 675654
rect 566186 675098 566422 675334
rect 566186 639418 566422 639654
rect 566186 639098 566422 639334
rect 566186 603418 566422 603654
rect 566186 603098 566422 603334
rect 566186 567418 566422 567654
rect 566186 567098 566422 567334
rect 566186 531418 566422 531654
rect 566186 531098 566422 531334
rect 566186 495418 566422 495654
rect 566186 495098 566422 495334
rect 566186 459418 566422 459654
rect 566186 459098 566422 459334
rect 566186 423418 566422 423654
rect 566186 423098 566422 423334
rect 566186 387418 566422 387654
rect 566186 387098 566422 387334
rect 566186 351418 566422 351654
rect 566186 351098 566422 351334
rect 566186 315418 566422 315654
rect 566186 315098 566422 315334
rect 566186 279418 566422 279654
rect 566186 279098 566422 279334
rect 566186 243418 566422 243654
rect 566186 243098 566422 243334
rect 566186 207418 566422 207654
rect 566186 207098 566422 207334
rect 566186 171418 566422 171654
rect 566186 171098 566422 171334
rect 566186 135418 566422 135654
rect 566186 135098 566422 135334
rect 566186 99418 566422 99654
rect 566186 99098 566422 99334
rect 566186 63418 566422 63654
rect 566186 63098 566422 63334
rect 566186 27418 566422 27654
rect 566186 27098 566422 27334
rect 566186 -5282 566422 -5046
rect 566186 -5602 566422 -5366
rect 592082 711182 592318 711418
rect 592082 710862 592318 711098
rect 591142 710242 591378 710478
rect 591142 709922 591378 710158
rect 590202 709302 590438 709538
rect 590202 708982 590438 709218
rect 589262 708362 589498 708598
rect 589262 708042 589498 708278
rect 588322 707422 588558 707658
rect 588322 707102 588558 707338
rect 580586 706482 580822 706718
rect 580586 706162 580822 706398
rect 569786 679018 570022 679254
rect 569786 678698 570022 678934
rect 569786 643018 570022 643254
rect 569786 642698 570022 642934
rect 569786 607018 570022 607254
rect 569786 606698 570022 606934
rect 569786 571018 570022 571254
rect 569786 570698 570022 570934
rect 569786 535018 570022 535254
rect 569786 534698 570022 534934
rect 569786 499018 570022 499254
rect 569786 498698 570022 498934
rect 569786 463018 570022 463254
rect 569786 462698 570022 462934
rect 569786 427018 570022 427254
rect 569786 426698 570022 426934
rect 569786 391018 570022 391254
rect 569786 390698 570022 390934
rect 569786 355018 570022 355254
rect 569786 354698 570022 354934
rect 569786 319018 570022 319254
rect 569786 318698 570022 318934
rect 569786 283018 570022 283254
rect 569786 282698 570022 282934
rect 569786 247018 570022 247254
rect 569786 246698 570022 246934
rect 569786 211018 570022 211254
rect 569786 210698 570022 210934
rect 569786 175018 570022 175254
rect 569786 174698 570022 174934
rect 569786 139018 570022 139254
rect 569786 138698 570022 138934
rect 569786 103018 570022 103254
rect 569786 102698 570022 102934
rect 569786 67018 570022 67254
rect 569786 66698 570022 66934
rect 569786 31018 570022 31254
rect 569786 30698 570022 30934
rect 551786 -6222 552022 -5986
rect 551786 -6542 552022 -6306
rect 576986 704602 577222 704838
rect 576986 704282 577222 704518
rect 576986 686218 577222 686454
rect 576986 685898 577222 686134
rect 576986 650218 577222 650454
rect 576986 649898 577222 650134
rect 576986 614218 577222 614454
rect 576986 613898 577222 614134
rect 576986 578218 577222 578454
rect 576986 577898 577222 578134
rect 576986 542218 577222 542454
rect 576986 541898 577222 542134
rect 576986 506218 577222 506454
rect 576986 505898 577222 506134
rect 576986 470218 577222 470454
rect 576986 469898 577222 470134
rect 576986 434218 577222 434454
rect 576986 433898 577222 434134
rect 576986 398218 577222 398454
rect 576986 397898 577222 398134
rect 576986 362218 577222 362454
rect 576986 361898 577222 362134
rect 576986 326218 577222 326454
rect 576986 325898 577222 326134
rect 576986 290218 577222 290454
rect 576986 289898 577222 290134
rect 576986 254218 577222 254454
rect 576986 253898 577222 254134
rect 576986 218218 577222 218454
rect 576986 217898 577222 218134
rect 576986 182218 577222 182454
rect 576986 181898 577222 182134
rect 576986 146218 577222 146454
rect 576986 145898 577222 146134
rect 576986 110218 577222 110454
rect 576986 109898 577222 110134
rect 576986 74218 577222 74454
rect 576986 73898 577222 74134
rect 576986 38218 577222 38454
rect 576986 37898 577222 38134
rect 576986 2218 577222 2454
rect 576986 1898 577222 2134
rect 576986 -582 577222 -346
rect 576986 -902 577222 -666
rect 587382 706482 587618 706718
rect 587382 706162 587618 706398
rect 586442 705542 586678 705778
rect 586442 705222 586678 705458
rect 580586 689818 580822 690054
rect 580586 689498 580822 689734
rect 580586 653818 580822 654054
rect 580586 653498 580822 653734
rect 580586 617818 580822 618054
rect 580586 617498 580822 617734
rect 580586 581818 580822 582054
rect 580586 581498 580822 581734
rect 580586 545818 580822 546054
rect 580586 545498 580822 545734
rect 580586 509818 580822 510054
rect 580586 509498 580822 509734
rect 580586 473818 580822 474054
rect 580586 473498 580822 473734
rect 580586 437818 580822 438054
rect 580586 437498 580822 437734
rect 580586 401818 580822 402054
rect 580586 401498 580822 401734
rect 580586 365818 580822 366054
rect 580586 365498 580822 365734
rect 580586 329818 580822 330054
rect 580586 329498 580822 329734
rect 580586 293818 580822 294054
rect 580586 293498 580822 293734
rect 580586 257818 580822 258054
rect 580586 257498 580822 257734
rect 580586 221818 580822 222054
rect 580586 221498 580822 221734
rect 580586 185818 580822 186054
rect 580586 185498 580822 185734
rect 580586 149818 580822 150054
rect 580586 149498 580822 149734
rect 580586 113818 580822 114054
rect 580586 113498 580822 113734
rect 580586 77818 580822 78054
rect 580586 77498 580822 77734
rect 580586 41818 580822 42054
rect 580586 41498 580822 41734
rect 580586 5818 580822 6054
rect 580586 5498 580822 5734
rect 585502 704602 585738 704838
rect 585502 704282 585738 704518
rect 585502 686218 585738 686454
rect 585502 685898 585738 686134
rect 585502 650218 585738 650454
rect 585502 649898 585738 650134
rect 585502 614218 585738 614454
rect 585502 613898 585738 614134
rect 585502 578218 585738 578454
rect 585502 577898 585738 578134
rect 585502 542218 585738 542454
rect 585502 541898 585738 542134
rect 585502 506218 585738 506454
rect 585502 505898 585738 506134
rect 585502 470218 585738 470454
rect 585502 469898 585738 470134
rect 585502 434218 585738 434454
rect 585502 433898 585738 434134
rect 585502 398218 585738 398454
rect 585502 397898 585738 398134
rect 585502 362218 585738 362454
rect 585502 361898 585738 362134
rect 585502 326218 585738 326454
rect 585502 325898 585738 326134
rect 585502 290218 585738 290454
rect 585502 289898 585738 290134
rect 585502 254218 585738 254454
rect 585502 253898 585738 254134
rect 585502 218218 585738 218454
rect 585502 217898 585738 218134
rect 585502 182218 585738 182454
rect 585502 181898 585738 182134
rect 585502 146218 585738 146454
rect 585502 145898 585738 146134
rect 585502 110218 585738 110454
rect 585502 109898 585738 110134
rect 585502 74218 585738 74454
rect 585502 73898 585738 74134
rect 585502 38218 585738 38454
rect 585502 37898 585738 38134
rect 585502 2218 585738 2454
rect 585502 1898 585738 2134
rect 585502 -582 585738 -346
rect 585502 -902 585738 -666
rect 586442 668218 586678 668454
rect 586442 667898 586678 668134
rect 586442 632218 586678 632454
rect 586442 631898 586678 632134
rect 586442 596218 586678 596454
rect 586442 595898 586678 596134
rect 586442 560218 586678 560454
rect 586442 559898 586678 560134
rect 586442 524218 586678 524454
rect 586442 523898 586678 524134
rect 586442 488218 586678 488454
rect 586442 487898 586678 488134
rect 586442 452218 586678 452454
rect 586442 451898 586678 452134
rect 586442 416218 586678 416454
rect 586442 415898 586678 416134
rect 586442 380218 586678 380454
rect 586442 379898 586678 380134
rect 586442 344218 586678 344454
rect 586442 343898 586678 344134
rect 586442 308218 586678 308454
rect 586442 307898 586678 308134
rect 586442 272218 586678 272454
rect 586442 271898 586678 272134
rect 586442 236218 586678 236454
rect 586442 235898 586678 236134
rect 586442 200218 586678 200454
rect 586442 199898 586678 200134
rect 586442 164218 586678 164454
rect 586442 163898 586678 164134
rect 586442 128218 586678 128454
rect 586442 127898 586678 128134
rect 586442 92218 586678 92454
rect 586442 91898 586678 92134
rect 586442 56218 586678 56454
rect 586442 55898 586678 56134
rect 586442 20218 586678 20454
rect 586442 19898 586678 20134
rect 586442 -1522 586678 -1286
rect 586442 -1842 586678 -1606
rect 587382 689818 587618 690054
rect 587382 689498 587618 689734
rect 587382 653818 587618 654054
rect 587382 653498 587618 653734
rect 587382 617818 587618 618054
rect 587382 617498 587618 617734
rect 587382 581818 587618 582054
rect 587382 581498 587618 581734
rect 587382 545818 587618 546054
rect 587382 545498 587618 545734
rect 587382 509818 587618 510054
rect 587382 509498 587618 509734
rect 587382 473818 587618 474054
rect 587382 473498 587618 473734
rect 587382 437818 587618 438054
rect 587382 437498 587618 437734
rect 587382 401818 587618 402054
rect 587382 401498 587618 401734
rect 587382 365818 587618 366054
rect 587382 365498 587618 365734
rect 587382 329818 587618 330054
rect 587382 329498 587618 329734
rect 587382 293818 587618 294054
rect 587382 293498 587618 293734
rect 587382 257818 587618 258054
rect 587382 257498 587618 257734
rect 587382 221818 587618 222054
rect 587382 221498 587618 221734
rect 587382 185818 587618 186054
rect 587382 185498 587618 185734
rect 587382 149818 587618 150054
rect 587382 149498 587618 149734
rect 587382 113818 587618 114054
rect 587382 113498 587618 113734
rect 587382 77818 587618 78054
rect 587382 77498 587618 77734
rect 587382 41818 587618 42054
rect 587382 41498 587618 41734
rect 587382 5818 587618 6054
rect 587382 5498 587618 5734
rect 580586 -2462 580822 -2226
rect 580586 -2782 580822 -2546
rect 587382 -2462 587618 -2226
rect 587382 -2782 587618 -2546
rect 588322 671818 588558 672054
rect 588322 671498 588558 671734
rect 588322 635818 588558 636054
rect 588322 635498 588558 635734
rect 588322 599818 588558 600054
rect 588322 599498 588558 599734
rect 588322 563818 588558 564054
rect 588322 563498 588558 563734
rect 588322 527818 588558 528054
rect 588322 527498 588558 527734
rect 588322 491818 588558 492054
rect 588322 491498 588558 491734
rect 588322 455818 588558 456054
rect 588322 455498 588558 455734
rect 588322 419818 588558 420054
rect 588322 419498 588558 419734
rect 588322 383818 588558 384054
rect 588322 383498 588558 383734
rect 588322 347818 588558 348054
rect 588322 347498 588558 347734
rect 588322 311818 588558 312054
rect 588322 311498 588558 311734
rect 588322 275818 588558 276054
rect 588322 275498 588558 275734
rect 588322 239818 588558 240054
rect 588322 239498 588558 239734
rect 588322 203818 588558 204054
rect 588322 203498 588558 203734
rect 588322 167818 588558 168054
rect 588322 167498 588558 167734
rect 588322 131818 588558 132054
rect 588322 131498 588558 131734
rect 588322 95818 588558 96054
rect 588322 95498 588558 95734
rect 588322 59818 588558 60054
rect 588322 59498 588558 59734
rect 588322 23818 588558 24054
rect 588322 23498 588558 23734
rect 588322 -3402 588558 -3166
rect 588322 -3722 588558 -3486
rect 589262 693418 589498 693654
rect 589262 693098 589498 693334
rect 589262 657418 589498 657654
rect 589262 657098 589498 657334
rect 589262 621418 589498 621654
rect 589262 621098 589498 621334
rect 589262 585418 589498 585654
rect 589262 585098 589498 585334
rect 589262 549418 589498 549654
rect 589262 549098 589498 549334
rect 589262 513418 589498 513654
rect 589262 513098 589498 513334
rect 589262 477418 589498 477654
rect 589262 477098 589498 477334
rect 589262 441418 589498 441654
rect 589262 441098 589498 441334
rect 589262 405418 589498 405654
rect 589262 405098 589498 405334
rect 589262 369418 589498 369654
rect 589262 369098 589498 369334
rect 589262 333418 589498 333654
rect 589262 333098 589498 333334
rect 589262 297418 589498 297654
rect 589262 297098 589498 297334
rect 589262 261418 589498 261654
rect 589262 261098 589498 261334
rect 589262 225418 589498 225654
rect 589262 225098 589498 225334
rect 589262 189418 589498 189654
rect 589262 189098 589498 189334
rect 589262 153418 589498 153654
rect 589262 153098 589498 153334
rect 589262 117418 589498 117654
rect 589262 117098 589498 117334
rect 589262 81418 589498 81654
rect 589262 81098 589498 81334
rect 589262 45418 589498 45654
rect 589262 45098 589498 45334
rect 589262 9418 589498 9654
rect 589262 9098 589498 9334
rect 589262 -4342 589498 -4106
rect 589262 -4662 589498 -4426
rect 590202 675418 590438 675654
rect 590202 675098 590438 675334
rect 590202 639418 590438 639654
rect 590202 639098 590438 639334
rect 590202 603418 590438 603654
rect 590202 603098 590438 603334
rect 590202 567418 590438 567654
rect 590202 567098 590438 567334
rect 590202 531418 590438 531654
rect 590202 531098 590438 531334
rect 590202 495418 590438 495654
rect 590202 495098 590438 495334
rect 590202 459418 590438 459654
rect 590202 459098 590438 459334
rect 590202 423418 590438 423654
rect 590202 423098 590438 423334
rect 590202 387418 590438 387654
rect 590202 387098 590438 387334
rect 590202 351418 590438 351654
rect 590202 351098 590438 351334
rect 590202 315418 590438 315654
rect 590202 315098 590438 315334
rect 590202 279418 590438 279654
rect 590202 279098 590438 279334
rect 590202 243418 590438 243654
rect 590202 243098 590438 243334
rect 590202 207418 590438 207654
rect 590202 207098 590438 207334
rect 590202 171418 590438 171654
rect 590202 171098 590438 171334
rect 590202 135418 590438 135654
rect 590202 135098 590438 135334
rect 590202 99418 590438 99654
rect 590202 99098 590438 99334
rect 590202 63418 590438 63654
rect 590202 63098 590438 63334
rect 590202 27418 590438 27654
rect 590202 27098 590438 27334
rect 590202 -5282 590438 -5046
rect 590202 -5602 590438 -5366
rect 591142 697018 591378 697254
rect 591142 696698 591378 696934
rect 591142 661018 591378 661254
rect 591142 660698 591378 660934
rect 591142 625018 591378 625254
rect 591142 624698 591378 624934
rect 591142 589018 591378 589254
rect 591142 588698 591378 588934
rect 591142 553018 591378 553254
rect 591142 552698 591378 552934
rect 591142 517018 591378 517254
rect 591142 516698 591378 516934
rect 591142 481018 591378 481254
rect 591142 480698 591378 480934
rect 591142 445018 591378 445254
rect 591142 444698 591378 444934
rect 591142 409018 591378 409254
rect 591142 408698 591378 408934
rect 591142 373018 591378 373254
rect 591142 372698 591378 372934
rect 591142 337018 591378 337254
rect 591142 336698 591378 336934
rect 591142 301018 591378 301254
rect 591142 300698 591378 300934
rect 591142 265018 591378 265254
rect 591142 264698 591378 264934
rect 591142 229018 591378 229254
rect 591142 228698 591378 228934
rect 591142 193018 591378 193254
rect 591142 192698 591378 192934
rect 591142 157018 591378 157254
rect 591142 156698 591378 156934
rect 591142 121018 591378 121254
rect 591142 120698 591378 120934
rect 591142 85018 591378 85254
rect 591142 84698 591378 84934
rect 591142 49018 591378 49254
rect 591142 48698 591378 48934
rect 591142 13018 591378 13254
rect 591142 12698 591378 12934
rect 591142 -6222 591378 -5986
rect 591142 -6542 591378 -6306
rect 592082 679018 592318 679254
rect 592082 678698 592318 678934
rect 592082 643018 592318 643254
rect 592082 642698 592318 642934
rect 592082 607018 592318 607254
rect 592082 606698 592318 606934
rect 592082 571018 592318 571254
rect 592082 570698 592318 570934
rect 592082 535018 592318 535254
rect 592082 534698 592318 534934
rect 592082 499018 592318 499254
rect 592082 498698 592318 498934
rect 592082 463018 592318 463254
rect 592082 462698 592318 462934
rect 592082 427018 592318 427254
rect 592082 426698 592318 426934
rect 592082 391018 592318 391254
rect 592082 390698 592318 390934
rect 592082 355018 592318 355254
rect 592082 354698 592318 354934
rect 592082 319018 592318 319254
rect 592082 318698 592318 318934
rect 592082 283018 592318 283254
rect 592082 282698 592318 282934
rect 592082 247018 592318 247254
rect 592082 246698 592318 246934
rect 592082 211018 592318 211254
rect 592082 210698 592318 210934
rect 592082 175018 592318 175254
rect 592082 174698 592318 174934
rect 592082 139018 592318 139254
rect 592082 138698 592318 138934
rect 592082 103018 592318 103254
rect 592082 102698 592318 102934
rect 592082 67018 592318 67254
rect 592082 66698 592318 66934
rect 592082 31018 592318 31254
rect 592082 30698 592318 30934
rect 569786 -7162 570022 -6926
rect 569786 -7482 570022 -7246
rect 592082 -7162 592318 -6926
rect 592082 -7482 592318 -7246
<< metal5 >>
rect -8576 711440 -7976 711442
rect 29604 711440 30204 711442
rect 65604 711440 66204 711442
rect 101604 711440 102204 711442
rect 137604 711440 138204 711442
rect 173604 711440 174204 711442
rect 209604 711440 210204 711442
rect 245604 711440 246204 711442
rect 281604 711440 282204 711442
rect 317604 711440 318204 711442
rect 353604 711440 354204 711442
rect 389604 711440 390204 711442
rect 425604 711440 426204 711442
rect 461604 711440 462204 711442
rect 497604 711440 498204 711442
rect 533604 711440 534204 711442
rect 569604 711440 570204 711442
rect 591900 711440 592500 711442
rect -8576 711418 592500 711440
rect -8576 711182 -8394 711418
rect -8158 711182 29786 711418
rect 30022 711182 65786 711418
rect 66022 711182 101786 711418
rect 102022 711182 137786 711418
rect 138022 711182 173786 711418
rect 174022 711182 209786 711418
rect 210022 711182 245786 711418
rect 246022 711182 281786 711418
rect 282022 711182 317786 711418
rect 318022 711182 353786 711418
rect 354022 711182 389786 711418
rect 390022 711182 425786 711418
rect 426022 711182 461786 711418
rect 462022 711182 497786 711418
rect 498022 711182 533786 711418
rect 534022 711182 569786 711418
rect 570022 711182 592082 711418
rect 592318 711182 592500 711418
rect -8576 711098 592500 711182
rect -8576 710862 -8394 711098
rect -8158 710862 29786 711098
rect 30022 710862 65786 711098
rect 66022 710862 101786 711098
rect 102022 710862 137786 711098
rect 138022 710862 173786 711098
rect 174022 710862 209786 711098
rect 210022 710862 245786 711098
rect 246022 710862 281786 711098
rect 282022 710862 317786 711098
rect 318022 710862 353786 711098
rect 354022 710862 389786 711098
rect 390022 710862 425786 711098
rect 426022 710862 461786 711098
rect 462022 710862 497786 711098
rect 498022 710862 533786 711098
rect 534022 710862 569786 711098
rect 570022 710862 592082 711098
rect 592318 710862 592500 711098
rect -8576 710840 592500 710862
rect -8576 710838 -7976 710840
rect 29604 710838 30204 710840
rect 65604 710838 66204 710840
rect 101604 710838 102204 710840
rect 137604 710838 138204 710840
rect 173604 710838 174204 710840
rect 209604 710838 210204 710840
rect 245604 710838 246204 710840
rect 281604 710838 282204 710840
rect 317604 710838 318204 710840
rect 353604 710838 354204 710840
rect 389604 710838 390204 710840
rect 425604 710838 426204 710840
rect 461604 710838 462204 710840
rect 497604 710838 498204 710840
rect 533604 710838 534204 710840
rect 569604 710838 570204 710840
rect 591900 710838 592500 710840
rect -7636 710500 -7036 710502
rect 11604 710500 12204 710502
rect 47604 710500 48204 710502
rect 83604 710500 84204 710502
rect 119604 710500 120204 710502
rect 155604 710500 156204 710502
rect 191604 710500 192204 710502
rect 227604 710500 228204 710502
rect 263604 710500 264204 710502
rect 299604 710500 300204 710502
rect 335604 710500 336204 710502
rect 371604 710500 372204 710502
rect 407604 710500 408204 710502
rect 443604 710500 444204 710502
rect 479604 710500 480204 710502
rect 515604 710500 516204 710502
rect 551604 710500 552204 710502
rect 590960 710500 591560 710502
rect -7636 710478 591560 710500
rect -7636 710242 -7454 710478
rect -7218 710242 11786 710478
rect 12022 710242 47786 710478
rect 48022 710242 83786 710478
rect 84022 710242 119786 710478
rect 120022 710242 155786 710478
rect 156022 710242 191786 710478
rect 192022 710242 227786 710478
rect 228022 710242 263786 710478
rect 264022 710242 299786 710478
rect 300022 710242 335786 710478
rect 336022 710242 371786 710478
rect 372022 710242 407786 710478
rect 408022 710242 443786 710478
rect 444022 710242 479786 710478
rect 480022 710242 515786 710478
rect 516022 710242 551786 710478
rect 552022 710242 591142 710478
rect 591378 710242 591560 710478
rect -7636 710158 591560 710242
rect -7636 709922 -7454 710158
rect -7218 709922 11786 710158
rect 12022 709922 47786 710158
rect 48022 709922 83786 710158
rect 84022 709922 119786 710158
rect 120022 709922 155786 710158
rect 156022 709922 191786 710158
rect 192022 709922 227786 710158
rect 228022 709922 263786 710158
rect 264022 709922 299786 710158
rect 300022 709922 335786 710158
rect 336022 709922 371786 710158
rect 372022 709922 407786 710158
rect 408022 709922 443786 710158
rect 444022 709922 479786 710158
rect 480022 709922 515786 710158
rect 516022 709922 551786 710158
rect 552022 709922 591142 710158
rect 591378 709922 591560 710158
rect -7636 709900 591560 709922
rect -7636 709898 -7036 709900
rect 11604 709898 12204 709900
rect 47604 709898 48204 709900
rect 83604 709898 84204 709900
rect 119604 709898 120204 709900
rect 155604 709898 156204 709900
rect 191604 709898 192204 709900
rect 227604 709898 228204 709900
rect 263604 709898 264204 709900
rect 299604 709898 300204 709900
rect 335604 709898 336204 709900
rect 371604 709898 372204 709900
rect 407604 709898 408204 709900
rect 443604 709898 444204 709900
rect 479604 709898 480204 709900
rect 515604 709898 516204 709900
rect 551604 709898 552204 709900
rect 590960 709898 591560 709900
rect -6696 709560 -6096 709562
rect 26004 709560 26604 709562
rect 62004 709560 62604 709562
rect 98004 709560 98604 709562
rect 134004 709560 134604 709562
rect 170004 709560 170604 709562
rect 206004 709560 206604 709562
rect 242004 709560 242604 709562
rect 278004 709560 278604 709562
rect 314004 709560 314604 709562
rect 350004 709560 350604 709562
rect 386004 709560 386604 709562
rect 422004 709560 422604 709562
rect 458004 709560 458604 709562
rect 494004 709560 494604 709562
rect 530004 709560 530604 709562
rect 566004 709560 566604 709562
rect 590020 709560 590620 709562
rect -6696 709538 590620 709560
rect -6696 709302 -6514 709538
rect -6278 709302 26186 709538
rect 26422 709302 62186 709538
rect 62422 709302 98186 709538
rect 98422 709302 134186 709538
rect 134422 709302 170186 709538
rect 170422 709302 206186 709538
rect 206422 709302 242186 709538
rect 242422 709302 278186 709538
rect 278422 709302 314186 709538
rect 314422 709302 350186 709538
rect 350422 709302 386186 709538
rect 386422 709302 422186 709538
rect 422422 709302 458186 709538
rect 458422 709302 494186 709538
rect 494422 709302 530186 709538
rect 530422 709302 566186 709538
rect 566422 709302 590202 709538
rect 590438 709302 590620 709538
rect -6696 709218 590620 709302
rect -6696 708982 -6514 709218
rect -6278 708982 26186 709218
rect 26422 708982 62186 709218
rect 62422 708982 98186 709218
rect 98422 708982 134186 709218
rect 134422 708982 170186 709218
rect 170422 708982 206186 709218
rect 206422 708982 242186 709218
rect 242422 708982 278186 709218
rect 278422 708982 314186 709218
rect 314422 708982 350186 709218
rect 350422 708982 386186 709218
rect 386422 708982 422186 709218
rect 422422 708982 458186 709218
rect 458422 708982 494186 709218
rect 494422 708982 530186 709218
rect 530422 708982 566186 709218
rect 566422 708982 590202 709218
rect 590438 708982 590620 709218
rect -6696 708960 590620 708982
rect -6696 708958 -6096 708960
rect 26004 708958 26604 708960
rect 62004 708958 62604 708960
rect 98004 708958 98604 708960
rect 134004 708958 134604 708960
rect 170004 708958 170604 708960
rect 206004 708958 206604 708960
rect 242004 708958 242604 708960
rect 278004 708958 278604 708960
rect 314004 708958 314604 708960
rect 350004 708958 350604 708960
rect 386004 708958 386604 708960
rect 422004 708958 422604 708960
rect 458004 708958 458604 708960
rect 494004 708958 494604 708960
rect 530004 708958 530604 708960
rect 566004 708958 566604 708960
rect 590020 708958 590620 708960
rect -5756 708620 -5156 708622
rect 8004 708620 8604 708622
rect 44004 708620 44604 708622
rect 80004 708620 80604 708622
rect 116004 708620 116604 708622
rect 152004 708620 152604 708622
rect 188004 708620 188604 708622
rect 224004 708620 224604 708622
rect 260004 708620 260604 708622
rect 296004 708620 296604 708622
rect 332004 708620 332604 708622
rect 368004 708620 368604 708622
rect 404004 708620 404604 708622
rect 440004 708620 440604 708622
rect 476004 708620 476604 708622
rect 512004 708620 512604 708622
rect 548004 708620 548604 708622
rect 589080 708620 589680 708622
rect -5756 708598 589680 708620
rect -5756 708362 -5574 708598
rect -5338 708362 8186 708598
rect 8422 708362 44186 708598
rect 44422 708362 80186 708598
rect 80422 708362 116186 708598
rect 116422 708362 152186 708598
rect 152422 708362 188186 708598
rect 188422 708362 224186 708598
rect 224422 708362 260186 708598
rect 260422 708362 296186 708598
rect 296422 708362 332186 708598
rect 332422 708362 368186 708598
rect 368422 708362 404186 708598
rect 404422 708362 440186 708598
rect 440422 708362 476186 708598
rect 476422 708362 512186 708598
rect 512422 708362 548186 708598
rect 548422 708362 589262 708598
rect 589498 708362 589680 708598
rect -5756 708278 589680 708362
rect -5756 708042 -5574 708278
rect -5338 708042 8186 708278
rect 8422 708042 44186 708278
rect 44422 708042 80186 708278
rect 80422 708042 116186 708278
rect 116422 708042 152186 708278
rect 152422 708042 188186 708278
rect 188422 708042 224186 708278
rect 224422 708042 260186 708278
rect 260422 708042 296186 708278
rect 296422 708042 332186 708278
rect 332422 708042 368186 708278
rect 368422 708042 404186 708278
rect 404422 708042 440186 708278
rect 440422 708042 476186 708278
rect 476422 708042 512186 708278
rect 512422 708042 548186 708278
rect 548422 708042 589262 708278
rect 589498 708042 589680 708278
rect -5756 708020 589680 708042
rect -5756 708018 -5156 708020
rect 8004 708018 8604 708020
rect 44004 708018 44604 708020
rect 80004 708018 80604 708020
rect 116004 708018 116604 708020
rect 152004 708018 152604 708020
rect 188004 708018 188604 708020
rect 224004 708018 224604 708020
rect 260004 708018 260604 708020
rect 296004 708018 296604 708020
rect 332004 708018 332604 708020
rect 368004 708018 368604 708020
rect 404004 708018 404604 708020
rect 440004 708018 440604 708020
rect 476004 708018 476604 708020
rect 512004 708018 512604 708020
rect 548004 708018 548604 708020
rect 589080 708018 589680 708020
rect -4816 707680 -4216 707682
rect 22404 707680 23004 707682
rect 58404 707680 59004 707682
rect 94404 707680 95004 707682
rect 130404 707680 131004 707682
rect 166404 707680 167004 707682
rect 202404 707680 203004 707682
rect 238404 707680 239004 707682
rect 274404 707680 275004 707682
rect 310404 707680 311004 707682
rect 346404 707680 347004 707682
rect 382404 707680 383004 707682
rect 418404 707680 419004 707682
rect 454404 707680 455004 707682
rect 490404 707680 491004 707682
rect 526404 707680 527004 707682
rect 562404 707680 563004 707682
rect 588140 707680 588740 707682
rect -4816 707658 588740 707680
rect -4816 707422 -4634 707658
rect -4398 707422 22586 707658
rect 22822 707422 58586 707658
rect 58822 707422 94586 707658
rect 94822 707422 130586 707658
rect 130822 707422 166586 707658
rect 166822 707422 202586 707658
rect 202822 707422 238586 707658
rect 238822 707422 274586 707658
rect 274822 707422 310586 707658
rect 310822 707422 346586 707658
rect 346822 707422 382586 707658
rect 382822 707422 418586 707658
rect 418822 707422 454586 707658
rect 454822 707422 490586 707658
rect 490822 707422 526586 707658
rect 526822 707422 562586 707658
rect 562822 707422 588322 707658
rect 588558 707422 588740 707658
rect -4816 707338 588740 707422
rect -4816 707102 -4634 707338
rect -4398 707102 22586 707338
rect 22822 707102 58586 707338
rect 58822 707102 94586 707338
rect 94822 707102 130586 707338
rect 130822 707102 166586 707338
rect 166822 707102 202586 707338
rect 202822 707102 238586 707338
rect 238822 707102 274586 707338
rect 274822 707102 310586 707338
rect 310822 707102 346586 707338
rect 346822 707102 382586 707338
rect 382822 707102 418586 707338
rect 418822 707102 454586 707338
rect 454822 707102 490586 707338
rect 490822 707102 526586 707338
rect 526822 707102 562586 707338
rect 562822 707102 588322 707338
rect 588558 707102 588740 707338
rect -4816 707080 588740 707102
rect -4816 707078 -4216 707080
rect 22404 707078 23004 707080
rect 58404 707078 59004 707080
rect 94404 707078 95004 707080
rect 130404 707078 131004 707080
rect 166404 707078 167004 707080
rect 202404 707078 203004 707080
rect 238404 707078 239004 707080
rect 274404 707078 275004 707080
rect 310404 707078 311004 707080
rect 346404 707078 347004 707080
rect 382404 707078 383004 707080
rect 418404 707078 419004 707080
rect 454404 707078 455004 707080
rect 490404 707078 491004 707080
rect 526404 707078 527004 707080
rect 562404 707078 563004 707080
rect 588140 707078 588740 707080
rect -3876 706740 -3276 706742
rect 4404 706740 5004 706742
rect 40404 706740 41004 706742
rect 76404 706740 77004 706742
rect 112404 706740 113004 706742
rect 148404 706740 149004 706742
rect 184404 706740 185004 706742
rect 220404 706740 221004 706742
rect 256404 706740 257004 706742
rect 292404 706740 293004 706742
rect 328404 706740 329004 706742
rect 364404 706740 365004 706742
rect 400404 706740 401004 706742
rect 436404 706740 437004 706742
rect 472404 706740 473004 706742
rect 508404 706740 509004 706742
rect 544404 706740 545004 706742
rect 580404 706740 581004 706742
rect 587200 706740 587800 706742
rect -3876 706718 587800 706740
rect -3876 706482 -3694 706718
rect -3458 706482 4586 706718
rect 4822 706482 40586 706718
rect 40822 706482 76586 706718
rect 76822 706482 112586 706718
rect 112822 706482 148586 706718
rect 148822 706482 184586 706718
rect 184822 706482 220586 706718
rect 220822 706482 256586 706718
rect 256822 706482 292586 706718
rect 292822 706482 328586 706718
rect 328822 706482 364586 706718
rect 364822 706482 400586 706718
rect 400822 706482 436586 706718
rect 436822 706482 472586 706718
rect 472822 706482 508586 706718
rect 508822 706482 544586 706718
rect 544822 706482 580586 706718
rect 580822 706482 587382 706718
rect 587618 706482 587800 706718
rect -3876 706398 587800 706482
rect -3876 706162 -3694 706398
rect -3458 706162 4586 706398
rect 4822 706162 40586 706398
rect 40822 706162 76586 706398
rect 76822 706162 112586 706398
rect 112822 706162 148586 706398
rect 148822 706162 184586 706398
rect 184822 706162 220586 706398
rect 220822 706162 256586 706398
rect 256822 706162 292586 706398
rect 292822 706162 328586 706398
rect 328822 706162 364586 706398
rect 364822 706162 400586 706398
rect 400822 706162 436586 706398
rect 436822 706162 472586 706398
rect 472822 706162 508586 706398
rect 508822 706162 544586 706398
rect 544822 706162 580586 706398
rect 580822 706162 587382 706398
rect 587618 706162 587800 706398
rect -3876 706140 587800 706162
rect -3876 706138 -3276 706140
rect 4404 706138 5004 706140
rect 40404 706138 41004 706140
rect 76404 706138 77004 706140
rect 112404 706138 113004 706140
rect 148404 706138 149004 706140
rect 184404 706138 185004 706140
rect 220404 706138 221004 706140
rect 256404 706138 257004 706140
rect 292404 706138 293004 706140
rect 328404 706138 329004 706140
rect 364404 706138 365004 706140
rect 400404 706138 401004 706140
rect 436404 706138 437004 706140
rect 472404 706138 473004 706140
rect 508404 706138 509004 706140
rect 544404 706138 545004 706140
rect 580404 706138 581004 706140
rect 587200 706138 587800 706140
rect -2936 705800 -2336 705802
rect 18804 705800 19404 705802
rect 54804 705800 55404 705802
rect 90804 705800 91404 705802
rect 126804 705800 127404 705802
rect 162804 705800 163404 705802
rect 198804 705800 199404 705802
rect 234804 705800 235404 705802
rect 270804 705800 271404 705802
rect 306804 705800 307404 705802
rect 342804 705800 343404 705802
rect 378804 705800 379404 705802
rect 414804 705800 415404 705802
rect 450804 705800 451404 705802
rect 486804 705800 487404 705802
rect 522804 705800 523404 705802
rect 558804 705800 559404 705802
rect 586260 705800 586860 705802
rect -2936 705778 586860 705800
rect -2936 705542 -2754 705778
rect -2518 705542 18986 705778
rect 19222 705542 54986 705778
rect 55222 705542 90986 705778
rect 91222 705542 126986 705778
rect 127222 705542 162986 705778
rect 163222 705542 198986 705778
rect 199222 705542 234986 705778
rect 235222 705542 270986 705778
rect 271222 705542 306986 705778
rect 307222 705542 342986 705778
rect 343222 705542 378986 705778
rect 379222 705542 414986 705778
rect 415222 705542 450986 705778
rect 451222 705542 486986 705778
rect 487222 705542 522986 705778
rect 523222 705542 558986 705778
rect 559222 705542 586442 705778
rect 586678 705542 586860 705778
rect -2936 705458 586860 705542
rect -2936 705222 -2754 705458
rect -2518 705222 18986 705458
rect 19222 705222 54986 705458
rect 55222 705222 90986 705458
rect 91222 705222 126986 705458
rect 127222 705222 162986 705458
rect 163222 705222 198986 705458
rect 199222 705222 234986 705458
rect 235222 705222 270986 705458
rect 271222 705222 306986 705458
rect 307222 705222 342986 705458
rect 343222 705222 378986 705458
rect 379222 705222 414986 705458
rect 415222 705222 450986 705458
rect 451222 705222 486986 705458
rect 487222 705222 522986 705458
rect 523222 705222 558986 705458
rect 559222 705222 586442 705458
rect 586678 705222 586860 705458
rect -2936 705200 586860 705222
rect -2936 705198 -2336 705200
rect 18804 705198 19404 705200
rect 54804 705198 55404 705200
rect 90804 705198 91404 705200
rect 126804 705198 127404 705200
rect 162804 705198 163404 705200
rect 198804 705198 199404 705200
rect 234804 705198 235404 705200
rect 270804 705198 271404 705200
rect 306804 705198 307404 705200
rect 342804 705198 343404 705200
rect 378804 705198 379404 705200
rect 414804 705198 415404 705200
rect 450804 705198 451404 705200
rect 486804 705198 487404 705200
rect 522804 705198 523404 705200
rect 558804 705198 559404 705200
rect 586260 705198 586860 705200
rect -1996 704860 -1396 704862
rect 804 704860 1404 704862
rect 36804 704860 37404 704862
rect 72804 704860 73404 704862
rect 108804 704860 109404 704862
rect 144804 704860 145404 704862
rect 180804 704860 181404 704862
rect 216804 704860 217404 704862
rect 252804 704860 253404 704862
rect 288804 704860 289404 704862
rect 324804 704860 325404 704862
rect 360804 704860 361404 704862
rect 396804 704860 397404 704862
rect 432804 704860 433404 704862
rect 468804 704860 469404 704862
rect 504804 704860 505404 704862
rect 540804 704860 541404 704862
rect 576804 704860 577404 704862
rect 585320 704860 585920 704862
rect -1996 704838 585920 704860
rect -1996 704602 -1814 704838
rect -1578 704602 986 704838
rect 1222 704602 36986 704838
rect 37222 704602 72986 704838
rect 73222 704602 108986 704838
rect 109222 704602 144986 704838
rect 145222 704602 180986 704838
rect 181222 704602 216986 704838
rect 217222 704602 252986 704838
rect 253222 704602 288986 704838
rect 289222 704602 324986 704838
rect 325222 704602 360986 704838
rect 361222 704602 396986 704838
rect 397222 704602 432986 704838
rect 433222 704602 468986 704838
rect 469222 704602 504986 704838
rect 505222 704602 540986 704838
rect 541222 704602 576986 704838
rect 577222 704602 585502 704838
rect 585738 704602 585920 704838
rect -1996 704518 585920 704602
rect -1996 704282 -1814 704518
rect -1578 704282 986 704518
rect 1222 704282 36986 704518
rect 37222 704282 72986 704518
rect 73222 704282 108986 704518
rect 109222 704282 144986 704518
rect 145222 704282 180986 704518
rect 181222 704282 216986 704518
rect 217222 704282 252986 704518
rect 253222 704282 288986 704518
rect 289222 704282 324986 704518
rect 325222 704282 360986 704518
rect 361222 704282 396986 704518
rect 397222 704282 432986 704518
rect 433222 704282 468986 704518
rect 469222 704282 504986 704518
rect 505222 704282 540986 704518
rect 541222 704282 576986 704518
rect 577222 704282 585502 704518
rect 585738 704282 585920 704518
rect -1996 704260 585920 704282
rect -1996 704258 -1396 704260
rect 804 704258 1404 704260
rect 36804 704258 37404 704260
rect 72804 704258 73404 704260
rect 108804 704258 109404 704260
rect 144804 704258 145404 704260
rect 180804 704258 181404 704260
rect 216804 704258 217404 704260
rect 252804 704258 253404 704260
rect 288804 704258 289404 704260
rect 324804 704258 325404 704260
rect 360804 704258 361404 704260
rect 396804 704258 397404 704260
rect 432804 704258 433404 704260
rect 468804 704258 469404 704260
rect 504804 704258 505404 704260
rect 540804 704258 541404 704260
rect 576804 704258 577404 704260
rect 585320 704258 585920 704260
rect -7636 697276 -7036 697278
rect 11604 697276 12204 697278
rect 47604 697276 48204 697278
rect 83604 697276 84204 697278
rect 119604 697276 120204 697278
rect 155604 697276 156204 697278
rect 191604 697276 192204 697278
rect 227604 697276 228204 697278
rect 263604 697276 264204 697278
rect 299604 697276 300204 697278
rect 335604 697276 336204 697278
rect 371604 697276 372204 697278
rect 407604 697276 408204 697278
rect 443604 697276 444204 697278
rect 479604 697276 480204 697278
rect 515604 697276 516204 697278
rect 551604 697276 552204 697278
rect 590960 697276 591560 697278
rect -8576 697254 592500 697276
rect -8576 697018 -7454 697254
rect -7218 697018 11786 697254
rect 12022 697018 47786 697254
rect 48022 697018 83786 697254
rect 84022 697018 119786 697254
rect 120022 697018 155786 697254
rect 156022 697018 191786 697254
rect 192022 697018 227786 697254
rect 228022 697018 263786 697254
rect 264022 697018 299786 697254
rect 300022 697018 335786 697254
rect 336022 697018 371786 697254
rect 372022 697018 407786 697254
rect 408022 697018 443786 697254
rect 444022 697018 479786 697254
rect 480022 697018 515786 697254
rect 516022 697018 551786 697254
rect 552022 697018 591142 697254
rect 591378 697018 592500 697254
rect -8576 696934 592500 697018
rect -8576 696698 -7454 696934
rect -7218 696698 11786 696934
rect 12022 696698 47786 696934
rect 48022 696698 83786 696934
rect 84022 696698 119786 696934
rect 120022 696698 155786 696934
rect 156022 696698 191786 696934
rect 192022 696698 227786 696934
rect 228022 696698 263786 696934
rect 264022 696698 299786 696934
rect 300022 696698 335786 696934
rect 336022 696698 371786 696934
rect 372022 696698 407786 696934
rect 408022 696698 443786 696934
rect 444022 696698 479786 696934
rect 480022 696698 515786 696934
rect 516022 696698 551786 696934
rect 552022 696698 591142 696934
rect 591378 696698 592500 696934
rect -8576 696676 592500 696698
rect -7636 696674 -7036 696676
rect 11604 696674 12204 696676
rect 47604 696674 48204 696676
rect 83604 696674 84204 696676
rect 119604 696674 120204 696676
rect 155604 696674 156204 696676
rect 191604 696674 192204 696676
rect 227604 696674 228204 696676
rect 263604 696674 264204 696676
rect 299604 696674 300204 696676
rect 335604 696674 336204 696676
rect 371604 696674 372204 696676
rect 407604 696674 408204 696676
rect 443604 696674 444204 696676
rect 479604 696674 480204 696676
rect 515604 696674 516204 696676
rect 551604 696674 552204 696676
rect 590960 696674 591560 696676
rect -5756 693676 -5156 693678
rect 8004 693676 8604 693678
rect 44004 693676 44604 693678
rect 80004 693676 80604 693678
rect 116004 693676 116604 693678
rect 152004 693676 152604 693678
rect 188004 693676 188604 693678
rect 224004 693676 224604 693678
rect 260004 693676 260604 693678
rect 296004 693676 296604 693678
rect 332004 693676 332604 693678
rect 368004 693676 368604 693678
rect 404004 693676 404604 693678
rect 440004 693676 440604 693678
rect 476004 693676 476604 693678
rect 512004 693676 512604 693678
rect 548004 693676 548604 693678
rect 589080 693676 589680 693678
rect -6696 693654 590620 693676
rect -6696 693418 -5574 693654
rect -5338 693418 8186 693654
rect 8422 693418 44186 693654
rect 44422 693418 80186 693654
rect 80422 693418 116186 693654
rect 116422 693418 152186 693654
rect 152422 693418 188186 693654
rect 188422 693418 224186 693654
rect 224422 693418 260186 693654
rect 260422 693418 296186 693654
rect 296422 693418 332186 693654
rect 332422 693418 368186 693654
rect 368422 693418 404186 693654
rect 404422 693418 440186 693654
rect 440422 693418 476186 693654
rect 476422 693418 512186 693654
rect 512422 693418 548186 693654
rect 548422 693418 589262 693654
rect 589498 693418 590620 693654
rect -6696 693334 590620 693418
rect -6696 693098 -5574 693334
rect -5338 693098 8186 693334
rect 8422 693098 44186 693334
rect 44422 693098 80186 693334
rect 80422 693098 116186 693334
rect 116422 693098 152186 693334
rect 152422 693098 188186 693334
rect 188422 693098 224186 693334
rect 224422 693098 260186 693334
rect 260422 693098 296186 693334
rect 296422 693098 332186 693334
rect 332422 693098 368186 693334
rect 368422 693098 404186 693334
rect 404422 693098 440186 693334
rect 440422 693098 476186 693334
rect 476422 693098 512186 693334
rect 512422 693098 548186 693334
rect 548422 693098 589262 693334
rect 589498 693098 590620 693334
rect -6696 693076 590620 693098
rect -5756 693074 -5156 693076
rect 8004 693074 8604 693076
rect 44004 693074 44604 693076
rect 80004 693074 80604 693076
rect 116004 693074 116604 693076
rect 152004 693074 152604 693076
rect 188004 693074 188604 693076
rect 224004 693074 224604 693076
rect 260004 693074 260604 693076
rect 296004 693074 296604 693076
rect 332004 693074 332604 693076
rect 368004 693074 368604 693076
rect 404004 693074 404604 693076
rect 440004 693074 440604 693076
rect 476004 693074 476604 693076
rect 512004 693074 512604 693076
rect 548004 693074 548604 693076
rect 589080 693074 589680 693076
rect -3876 690076 -3276 690078
rect 4404 690076 5004 690078
rect 40404 690076 41004 690078
rect 76404 690076 77004 690078
rect 112404 690076 113004 690078
rect 148404 690076 149004 690078
rect 184404 690076 185004 690078
rect 220404 690076 221004 690078
rect 256404 690076 257004 690078
rect 292404 690076 293004 690078
rect 328404 690076 329004 690078
rect 364404 690076 365004 690078
rect 400404 690076 401004 690078
rect 436404 690076 437004 690078
rect 472404 690076 473004 690078
rect 508404 690076 509004 690078
rect 544404 690076 545004 690078
rect 580404 690076 581004 690078
rect 587200 690076 587800 690078
rect -4816 690054 588740 690076
rect -4816 689818 -3694 690054
rect -3458 689818 4586 690054
rect 4822 689818 40586 690054
rect 40822 689818 76586 690054
rect 76822 689818 112586 690054
rect 112822 689818 148586 690054
rect 148822 689818 184586 690054
rect 184822 689818 220586 690054
rect 220822 689818 256586 690054
rect 256822 689818 292586 690054
rect 292822 689818 328586 690054
rect 328822 689818 364586 690054
rect 364822 689818 400586 690054
rect 400822 689818 436586 690054
rect 436822 689818 472586 690054
rect 472822 689818 508586 690054
rect 508822 689818 544586 690054
rect 544822 689818 580586 690054
rect 580822 689818 587382 690054
rect 587618 689818 588740 690054
rect -4816 689734 588740 689818
rect -4816 689498 -3694 689734
rect -3458 689498 4586 689734
rect 4822 689498 40586 689734
rect 40822 689498 76586 689734
rect 76822 689498 112586 689734
rect 112822 689498 148586 689734
rect 148822 689498 184586 689734
rect 184822 689498 220586 689734
rect 220822 689498 256586 689734
rect 256822 689498 292586 689734
rect 292822 689498 328586 689734
rect 328822 689498 364586 689734
rect 364822 689498 400586 689734
rect 400822 689498 436586 689734
rect 436822 689498 472586 689734
rect 472822 689498 508586 689734
rect 508822 689498 544586 689734
rect 544822 689498 580586 689734
rect 580822 689498 587382 689734
rect 587618 689498 588740 689734
rect -4816 689476 588740 689498
rect -3876 689474 -3276 689476
rect 4404 689474 5004 689476
rect 40404 689474 41004 689476
rect 76404 689474 77004 689476
rect 112404 689474 113004 689476
rect 148404 689474 149004 689476
rect 184404 689474 185004 689476
rect 220404 689474 221004 689476
rect 256404 689474 257004 689476
rect 292404 689474 293004 689476
rect 328404 689474 329004 689476
rect 364404 689474 365004 689476
rect 400404 689474 401004 689476
rect 436404 689474 437004 689476
rect 472404 689474 473004 689476
rect 508404 689474 509004 689476
rect 544404 689474 545004 689476
rect 580404 689474 581004 689476
rect 587200 689474 587800 689476
rect -1996 686476 -1396 686478
rect 804 686476 1404 686478
rect 36804 686476 37404 686478
rect 72804 686476 73404 686478
rect 108804 686476 109404 686478
rect 144804 686476 145404 686478
rect 180804 686476 181404 686478
rect 216804 686476 217404 686478
rect 252804 686476 253404 686478
rect 288804 686476 289404 686478
rect 324804 686476 325404 686478
rect 360804 686476 361404 686478
rect 396804 686476 397404 686478
rect 432804 686476 433404 686478
rect 468804 686476 469404 686478
rect 504804 686476 505404 686478
rect 540804 686476 541404 686478
rect 576804 686476 577404 686478
rect 585320 686476 585920 686478
rect -2936 686454 586860 686476
rect -2936 686218 -1814 686454
rect -1578 686218 986 686454
rect 1222 686218 36986 686454
rect 37222 686218 72986 686454
rect 73222 686218 108986 686454
rect 109222 686218 144986 686454
rect 145222 686218 180986 686454
rect 181222 686218 216986 686454
rect 217222 686218 252986 686454
rect 253222 686218 288986 686454
rect 289222 686218 324986 686454
rect 325222 686218 360986 686454
rect 361222 686218 396986 686454
rect 397222 686218 432986 686454
rect 433222 686218 468986 686454
rect 469222 686218 504986 686454
rect 505222 686218 540986 686454
rect 541222 686218 576986 686454
rect 577222 686218 585502 686454
rect 585738 686218 586860 686454
rect -2936 686134 586860 686218
rect -2936 685898 -1814 686134
rect -1578 685898 986 686134
rect 1222 685898 36986 686134
rect 37222 685898 72986 686134
rect 73222 685898 108986 686134
rect 109222 685898 144986 686134
rect 145222 685898 180986 686134
rect 181222 685898 216986 686134
rect 217222 685898 252986 686134
rect 253222 685898 288986 686134
rect 289222 685898 324986 686134
rect 325222 685898 360986 686134
rect 361222 685898 396986 686134
rect 397222 685898 432986 686134
rect 433222 685898 468986 686134
rect 469222 685898 504986 686134
rect 505222 685898 540986 686134
rect 541222 685898 576986 686134
rect 577222 685898 585502 686134
rect 585738 685898 586860 686134
rect -2936 685876 586860 685898
rect -1996 685874 -1396 685876
rect 804 685874 1404 685876
rect 36804 685874 37404 685876
rect 72804 685874 73404 685876
rect 108804 685874 109404 685876
rect 144804 685874 145404 685876
rect 180804 685874 181404 685876
rect 216804 685874 217404 685876
rect 252804 685874 253404 685876
rect 288804 685874 289404 685876
rect 324804 685874 325404 685876
rect 360804 685874 361404 685876
rect 396804 685874 397404 685876
rect 432804 685874 433404 685876
rect 468804 685874 469404 685876
rect 504804 685874 505404 685876
rect 540804 685874 541404 685876
rect 576804 685874 577404 685876
rect 585320 685874 585920 685876
rect -8576 679276 -7976 679278
rect 29604 679276 30204 679278
rect 65604 679276 66204 679278
rect 101604 679276 102204 679278
rect 137604 679276 138204 679278
rect 173604 679276 174204 679278
rect 209604 679276 210204 679278
rect 245604 679276 246204 679278
rect 281604 679276 282204 679278
rect 317604 679276 318204 679278
rect 353604 679276 354204 679278
rect 389604 679276 390204 679278
rect 425604 679276 426204 679278
rect 461604 679276 462204 679278
rect 497604 679276 498204 679278
rect 533604 679276 534204 679278
rect 569604 679276 570204 679278
rect 591900 679276 592500 679278
rect -8576 679254 592500 679276
rect -8576 679018 -8394 679254
rect -8158 679018 29786 679254
rect 30022 679018 65786 679254
rect 66022 679018 101786 679254
rect 102022 679018 137786 679254
rect 138022 679018 173786 679254
rect 174022 679018 209786 679254
rect 210022 679018 245786 679254
rect 246022 679018 281786 679254
rect 282022 679018 317786 679254
rect 318022 679018 353786 679254
rect 354022 679018 389786 679254
rect 390022 679018 425786 679254
rect 426022 679018 461786 679254
rect 462022 679018 497786 679254
rect 498022 679018 533786 679254
rect 534022 679018 569786 679254
rect 570022 679018 592082 679254
rect 592318 679018 592500 679254
rect -8576 678934 592500 679018
rect -8576 678698 -8394 678934
rect -8158 678698 29786 678934
rect 30022 678698 65786 678934
rect 66022 678698 101786 678934
rect 102022 678698 137786 678934
rect 138022 678698 173786 678934
rect 174022 678698 209786 678934
rect 210022 678698 245786 678934
rect 246022 678698 281786 678934
rect 282022 678698 317786 678934
rect 318022 678698 353786 678934
rect 354022 678698 389786 678934
rect 390022 678698 425786 678934
rect 426022 678698 461786 678934
rect 462022 678698 497786 678934
rect 498022 678698 533786 678934
rect 534022 678698 569786 678934
rect 570022 678698 592082 678934
rect 592318 678698 592500 678934
rect -8576 678676 592500 678698
rect -8576 678674 -7976 678676
rect 29604 678674 30204 678676
rect 65604 678674 66204 678676
rect 101604 678674 102204 678676
rect 137604 678674 138204 678676
rect 173604 678674 174204 678676
rect 209604 678674 210204 678676
rect 245604 678674 246204 678676
rect 281604 678674 282204 678676
rect 317604 678674 318204 678676
rect 353604 678674 354204 678676
rect 389604 678674 390204 678676
rect 425604 678674 426204 678676
rect 461604 678674 462204 678676
rect 497604 678674 498204 678676
rect 533604 678674 534204 678676
rect 569604 678674 570204 678676
rect 591900 678674 592500 678676
rect -6696 675676 -6096 675678
rect 26004 675676 26604 675678
rect 62004 675676 62604 675678
rect 98004 675676 98604 675678
rect 134004 675676 134604 675678
rect 170004 675676 170604 675678
rect 206004 675676 206604 675678
rect 242004 675676 242604 675678
rect 278004 675676 278604 675678
rect 314004 675676 314604 675678
rect 350004 675676 350604 675678
rect 386004 675676 386604 675678
rect 422004 675676 422604 675678
rect 458004 675676 458604 675678
rect 494004 675676 494604 675678
rect 530004 675676 530604 675678
rect 566004 675676 566604 675678
rect 590020 675676 590620 675678
rect -6696 675654 590620 675676
rect -6696 675418 -6514 675654
rect -6278 675418 26186 675654
rect 26422 675418 62186 675654
rect 62422 675418 98186 675654
rect 98422 675418 134186 675654
rect 134422 675418 170186 675654
rect 170422 675418 206186 675654
rect 206422 675418 242186 675654
rect 242422 675418 278186 675654
rect 278422 675418 314186 675654
rect 314422 675418 350186 675654
rect 350422 675418 386186 675654
rect 386422 675418 422186 675654
rect 422422 675418 458186 675654
rect 458422 675418 494186 675654
rect 494422 675418 530186 675654
rect 530422 675418 566186 675654
rect 566422 675418 590202 675654
rect 590438 675418 590620 675654
rect -6696 675334 590620 675418
rect -6696 675098 -6514 675334
rect -6278 675098 26186 675334
rect 26422 675098 62186 675334
rect 62422 675098 98186 675334
rect 98422 675098 134186 675334
rect 134422 675098 170186 675334
rect 170422 675098 206186 675334
rect 206422 675098 242186 675334
rect 242422 675098 278186 675334
rect 278422 675098 314186 675334
rect 314422 675098 350186 675334
rect 350422 675098 386186 675334
rect 386422 675098 422186 675334
rect 422422 675098 458186 675334
rect 458422 675098 494186 675334
rect 494422 675098 530186 675334
rect 530422 675098 566186 675334
rect 566422 675098 590202 675334
rect 590438 675098 590620 675334
rect -6696 675076 590620 675098
rect -6696 675074 -6096 675076
rect 26004 675074 26604 675076
rect 62004 675074 62604 675076
rect 98004 675074 98604 675076
rect 134004 675074 134604 675076
rect 170004 675074 170604 675076
rect 206004 675074 206604 675076
rect 242004 675074 242604 675076
rect 278004 675074 278604 675076
rect 314004 675074 314604 675076
rect 350004 675074 350604 675076
rect 386004 675074 386604 675076
rect 422004 675074 422604 675076
rect 458004 675074 458604 675076
rect 494004 675074 494604 675076
rect 530004 675074 530604 675076
rect 566004 675074 566604 675076
rect 590020 675074 590620 675076
rect -4816 672076 -4216 672078
rect 22404 672076 23004 672078
rect 58404 672076 59004 672078
rect 94404 672076 95004 672078
rect 130404 672076 131004 672078
rect 166404 672076 167004 672078
rect 202404 672076 203004 672078
rect 238404 672076 239004 672078
rect 274404 672076 275004 672078
rect 310404 672076 311004 672078
rect 346404 672076 347004 672078
rect 382404 672076 383004 672078
rect 418404 672076 419004 672078
rect 454404 672076 455004 672078
rect 490404 672076 491004 672078
rect 526404 672076 527004 672078
rect 562404 672076 563004 672078
rect 588140 672076 588740 672078
rect -4816 672054 588740 672076
rect -4816 671818 -4634 672054
rect -4398 671818 22586 672054
rect 22822 671818 58586 672054
rect 58822 671818 94586 672054
rect 94822 671818 130586 672054
rect 130822 671818 166586 672054
rect 166822 671818 202586 672054
rect 202822 671818 238586 672054
rect 238822 671818 274586 672054
rect 274822 671818 310586 672054
rect 310822 671818 346586 672054
rect 346822 671818 382586 672054
rect 382822 671818 418586 672054
rect 418822 671818 454586 672054
rect 454822 671818 490586 672054
rect 490822 671818 526586 672054
rect 526822 671818 562586 672054
rect 562822 671818 588322 672054
rect 588558 671818 588740 672054
rect -4816 671734 588740 671818
rect -4816 671498 -4634 671734
rect -4398 671498 22586 671734
rect 22822 671498 58586 671734
rect 58822 671498 94586 671734
rect 94822 671498 130586 671734
rect 130822 671498 166586 671734
rect 166822 671498 202586 671734
rect 202822 671498 238586 671734
rect 238822 671498 274586 671734
rect 274822 671498 310586 671734
rect 310822 671498 346586 671734
rect 346822 671498 382586 671734
rect 382822 671498 418586 671734
rect 418822 671498 454586 671734
rect 454822 671498 490586 671734
rect 490822 671498 526586 671734
rect 526822 671498 562586 671734
rect 562822 671498 588322 671734
rect 588558 671498 588740 671734
rect -4816 671476 588740 671498
rect -4816 671474 -4216 671476
rect 22404 671474 23004 671476
rect 58404 671474 59004 671476
rect 94404 671474 95004 671476
rect 130404 671474 131004 671476
rect 166404 671474 167004 671476
rect 202404 671474 203004 671476
rect 238404 671474 239004 671476
rect 274404 671474 275004 671476
rect 310404 671474 311004 671476
rect 346404 671474 347004 671476
rect 382404 671474 383004 671476
rect 418404 671474 419004 671476
rect 454404 671474 455004 671476
rect 490404 671474 491004 671476
rect 526404 671474 527004 671476
rect 562404 671474 563004 671476
rect 588140 671474 588740 671476
rect -2936 668476 -2336 668478
rect 18804 668476 19404 668478
rect 54804 668476 55404 668478
rect 90804 668476 91404 668478
rect 126804 668476 127404 668478
rect 162804 668476 163404 668478
rect 198804 668476 199404 668478
rect 234804 668476 235404 668478
rect 270804 668476 271404 668478
rect 306804 668476 307404 668478
rect 342804 668476 343404 668478
rect 378804 668476 379404 668478
rect 414804 668476 415404 668478
rect 450804 668476 451404 668478
rect 486804 668476 487404 668478
rect 522804 668476 523404 668478
rect 558804 668476 559404 668478
rect 586260 668476 586860 668478
rect -2936 668454 586860 668476
rect -2936 668218 -2754 668454
rect -2518 668218 18986 668454
rect 19222 668218 54986 668454
rect 55222 668218 90986 668454
rect 91222 668218 126986 668454
rect 127222 668218 162986 668454
rect 163222 668218 198986 668454
rect 199222 668218 234986 668454
rect 235222 668218 270986 668454
rect 271222 668218 306986 668454
rect 307222 668218 342986 668454
rect 343222 668218 378986 668454
rect 379222 668218 414986 668454
rect 415222 668218 450986 668454
rect 451222 668218 486986 668454
rect 487222 668218 522986 668454
rect 523222 668218 558986 668454
rect 559222 668218 586442 668454
rect 586678 668218 586860 668454
rect -2936 668134 586860 668218
rect -2936 667898 -2754 668134
rect -2518 667898 18986 668134
rect 19222 667898 54986 668134
rect 55222 667898 90986 668134
rect 91222 667898 126986 668134
rect 127222 667898 162986 668134
rect 163222 667898 198986 668134
rect 199222 667898 234986 668134
rect 235222 667898 270986 668134
rect 271222 667898 306986 668134
rect 307222 667898 342986 668134
rect 343222 667898 378986 668134
rect 379222 667898 414986 668134
rect 415222 667898 450986 668134
rect 451222 667898 486986 668134
rect 487222 667898 522986 668134
rect 523222 667898 558986 668134
rect 559222 667898 586442 668134
rect 586678 667898 586860 668134
rect -2936 667876 586860 667898
rect -2936 667874 -2336 667876
rect 18804 667874 19404 667876
rect 54804 667874 55404 667876
rect 90804 667874 91404 667876
rect 126804 667874 127404 667876
rect 162804 667874 163404 667876
rect 198804 667874 199404 667876
rect 234804 667874 235404 667876
rect 270804 667874 271404 667876
rect 306804 667874 307404 667876
rect 342804 667874 343404 667876
rect 378804 667874 379404 667876
rect 414804 667874 415404 667876
rect 450804 667874 451404 667876
rect 486804 667874 487404 667876
rect 522804 667874 523404 667876
rect 558804 667874 559404 667876
rect 586260 667874 586860 667876
rect -7636 661276 -7036 661278
rect 11604 661276 12204 661278
rect 47604 661276 48204 661278
rect 83604 661276 84204 661278
rect 119604 661276 120204 661278
rect 155604 661276 156204 661278
rect 191604 661276 192204 661278
rect 227604 661276 228204 661278
rect 263604 661276 264204 661278
rect 299604 661276 300204 661278
rect 335604 661276 336204 661278
rect 371604 661276 372204 661278
rect 407604 661276 408204 661278
rect 443604 661276 444204 661278
rect 479604 661276 480204 661278
rect 515604 661276 516204 661278
rect 551604 661276 552204 661278
rect 590960 661276 591560 661278
rect -8576 661254 592500 661276
rect -8576 661018 -7454 661254
rect -7218 661018 11786 661254
rect 12022 661018 47786 661254
rect 48022 661018 83786 661254
rect 84022 661018 119786 661254
rect 120022 661018 155786 661254
rect 156022 661018 191786 661254
rect 192022 661018 227786 661254
rect 228022 661018 263786 661254
rect 264022 661018 299786 661254
rect 300022 661018 335786 661254
rect 336022 661018 371786 661254
rect 372022 661018 407786 661254
rect 408022 661018 443786 661254
rect 444022 661018 479786 661254
rect 480022 661018 515786 661254
rect 516022 661018 551786 661254
rect 552022 661018 591142 661254
rect 591378 661018 592500 661254
rect -8576 660934 592500 661018
rect -8576 660698 -7454 660934
rect -7218 660698 11786 660934
rect 12022 660698 47786 660934
rect 48022 660698 83786 660934
rect 84022 660698 119786 660934
rect 120022 660698 155786 660934
rect 156022 660698 191786 660934
rect 192022 660698 227786 660934
rect 228022 660698 263786 660934
rect 264022 660698 299786 660934
rect 300022 660698 335786 660934
rect 336022 660698 371786 660934
rect 372022 660698 407786 660934
rect 408022 660698 443786 660934
rect 444022 660698 479786 660934
rect 480022 660698 515786 660934
rect 516022 660698 551786 660934
rect 552022 660698 591142 660934
rect 591378 660698 592500 660934
rect -8576 660676 592500 660698
rect -7636 660674 -7036 660676
rect 11604 660674 12204 660676
rect 47604 660674 48204 660676
rect 83604 660674 84204 660676
rect 119604 660674 120204 660676
rect 155604 660674 156204 660676
rect 191604 660674 192204 660676
rect 227604 660674 228204 660676
rect 263604 660674 264204 660676
rect 299604 660674 300204 660676
rect 335604 660674 336204 660676
rect 371604 660674 372204 660676
rect 407604 660674 408204 660676
rect 443604 660674 444204 660676
rect 479604 660674 480204 660676
rect 515604 660674 516204 660676
rect 551604 660674 552204 660676
rect 590960 660674 591560 660676
rect -5756 657676 -5156 657678
rect 8004 657676 8604 657678
rect 44004 657676 44604 657678
rect 80004 657676 80604 657678
rect 116004 657676 116604 657678
rect 152004 657676 152604 657678
rect 188004 657676 188604 657678
rect 224004 657676 224604 657678
rect 260004 657676 260604 657678
rect 296004 657676 296604 657678
rect 332004 657676 332604 657678
rect 368004 657676 368604 657678
rect 404004 657676 404604 657678
rect 440004 657676 440604 657678
rect 476004 657676 476604 657678
rect 512004 657676 512604 657678
rect 548004 657676 548604 657678
rect 589080 657676 589680 657678
rect -6696 657654 590620 657676
rect -6696 657418 -5574 657654
rect -5338 657418 8186 657654
rect 8422 657418 44186 657654
rect 44422 657418 80186 657654
rect 80422 657418 116186 657654
rect 116422 657418 152186 657654
rect 152422 657418 188186 657654
rect 188422 657418 224186 657654
rect 224422 657418 260186 657654
rect 260422 657418 296186 657654
rect 296422 657418 332186 657654
rect 332422 657418 368186 657654
rect 368422 657418 404186 657654
rect 404422 657418 440186 657654
rect 440422 657418 476186 657654
rect 476422 657418 512186 657654
rect 512422 657418 548186 657654
rect 548422 657418 589262 657654
rect 589498 657418 590620 657654
rect -6696 657334 590620 657418
rect -6696 657098 -5574 657334
rect -5338 657098 8186 657334
rect 8422 657098 44186 657334
rect 44422 657098 80186 657334
rect 80422 657098 116186 657334
rect 116422 657098 152186 657334
rect 152422 657098 188186 657334
rect 188422 657098 224186 657334
rect 224422 657098 260186 657334
rect 260422 657098 296186 657334
rect 296422 657098 332186 657334
rect 332422 657098 368186 657334
rect 368422 657098 404186 657334
rect 404422 657098 440186 657334
rect 440422 657098 476186 657334
rect 476422 657098 512186 657334
rect 512422 657098 548186 657334
rect 548422 657098 589262 657334
rect 589498 657098 590620 657334
rect -6696 657076 590620 657098
rect -5756 657074 -5156 657076
rect 8004 657074 8604 657076
rect 44004 657074 44604 657076
rect 80004 657074 80604 657076
rect 116004 657074 116604 657076
rect 152004 657074 152604 657076
rect 188004 657074 188604 657076
rect 224004 657074 224604 657076
rect 260004 657074 260604 657076
rect 296004 657074 296604 657076
rect 332004 657074 332604 657076
rect 368004 657074 368604 657076
rect 404004 657074 404604 657076
rect 440004 657074 440604 657076
rect 476004 657074 476604 657076
rect 512004 657074 512604 657076
rect 548004 657074 548604 657076
rect 589080 657074 589680 657076
rect -3876 654076 -3276 654078
rect 4404 654076 5004 654078
rect 40404 654076 41004 654078
rect 76404 654076 77004 654078
rect 112404 654076 113004 654078
rect 148404 654076 149004 654078
rect 184404 654076 185004 654078
rect 220404 654076 221004 654078
rect 256404 654076 257004 654078
rect 292404 654076 293004 654078
rect 328404 654076 329004 654078
rect 364404 654076 365004 654078
rect 400404 654076 401004 654078
rect 436404 654076 437004 654078
rect 472404 654076 473004 654078
rect 508404 654076 509004 654078
rect 544404 654076 545004 654078
rect 580404 654076 581004 654078
rect 587200 654076 587800 654078
rect -4816 654054 588740 654076
rect -4816 653818 -3694 654054
rect -3458 653818 4586 654054
rect 4822 653818 40586 654054
rect 40822 653818 76586 654054
rect 76822 653818 112586 654054
rect 112822 653818 148586 654054
rect 148822 653818 184586 654054
rect 184822 653818 220586 654054
rect 220822 653818 256586 654054
rect 256822 653818 292586 654054
rect 292822 653818 328586 654054
rect 328822 653818 364586 654054
rect 364822 653818 400586 654054
rect 400822 653818 436586 654054
rect 436822 653818 472586 654054
rect 472822 653818 508586 654054
rect 508822 653818 544586 654054
rect 544822 653818 580586 654054
rect 580822 653818 587382 654054
rect 587618 653818 588740 654054
rect -4816 653734 588740 653818
rect -4816 653498 -3694 653734
rect -3458 653498 4586 653734
rect 4822 653498 40586 653734
rect 40822 653498 76586 653734
rect 76822 653498 112586 653734
rect 112822 653498 148586 653734
rect 148822 653498 184586 653734
rect 184822 653498 220586 653734
rect 220822 653498 256586 653734
rect 256822 653498 292586 653734
rect 292822 653498 328586 653734
rect 328822 653498 364586 653734
rect 364822 653498 400586 653734
rect 400822 653498 436586 653734
rect 436822 653498 472586 653734
rect 472822 653498 508586 653734
rect 508822 653498 544586 653734
rect 544822 653498 580586 653734
rect 580822 653498 587382 653734
rect 587618 653498 588740 653734
rect -4816 653476 588740 653498
rect -3876 653474 -3276 653476
rect 4404 653474 5004 653476
rect 40404 653474 41004 653476
rect 76404 653474 77004 653476
rect 112404 653474 113004 653476
rect 148404 653474 149004 653476
rect 184404 653474 185004 653476
rect 220404 653474 221004 653476
rect 256404 653474 257004 653476
rect 292404 653474 293004 653476
rect 328404 653474 329004 653476
rect 364404 653474 365004 653476
rect 400404 653474 401004 653476
rect 436404 653474 437004 653476
rect 472404 653474 473004 653476
rect 508404 653474 509004 653476
rect 544404 653474 545004 653476
rect 580404 653474 581004 653476
rect 587200 653474 587800 653476
rect -1996 650476 -1396 650478
rect 804 650476 1404 650478
rect 36804 650476 37404 650478
rect 72804 650476 73404 650478
rect 108804 650476 109404 650478
rect 144804 650476 145404 650478
rect 180804 650476 181404 650478
rect 216804 650476 217404 650478
rect 252804 650476 253404 650478
rect 288804 650476 289404 650478
rect 324804 650476 325404 650478
rect 360804 650476 361404 650478
rect 396804 650476 397404 650478
rect 432804 650476 433404 650478
rect 468804 650476 469404 650478
rect 504804 650476 505404 650478
rect 540804 650476 541404 650478
rect 576804 650476 577404 650478
rect 585320 650476 585920 650478
rect -2936 650454 586860 650476
rect -2936 650218 -1814 650454
rect -1578 650218 986 650454
rect 1222 650218 36986 650454
rect 37222 650218 72986 650454
rect 73222 650218 108986 650454
rect 109222 650218 144986 650454
rect 145222 650218 180986 650454
rect 181222 650218 216986 650454
rect 217222 650218 252986 650454
rect 253222 650218 288986 650454
rect 289222 650218 324986 650454
rect 325222 650218 360986 650454
rect 361222 650218 396986 650454
rect 397222 650218 432986 650454
rect 433222 650218 468986 650454
rect 469222 650218 504986 650454
rect 505222 650218 540986 650454
rect 541222 650218 576986 650454
rect 577222 650218 585502 650454
rect 585738 650218 586860 650454
rect -2936 650134 586860 650218
rect -2936 649898 -1814 650134
rect -1578 649898 986 650134
rect 1222 649898 36986 650134
rect 37222 649898 72986 650134
rect 73222 649898 108986 650134
rect 109222 649898 144986 650134
rect 145222 649898 180986 650134
rect 181222 649898 216986 650134
rect 217222 649898 252986 650134
rect 253222 649898 288986 650134
rect 289222 649898 324986 650134
rect 325222 649898 360986 650134
rect 361222 649898 396986 650134
rect 397222 649898 432986 650134
rect 433222 649898 468986 650134
rect 469222 649898 504986 650134
rect 505222 649898 540986 650134
rect 541222 649898 576986 650134
rect 577222 649898 585502 650134
rect 585738 649898 586860 650134
rect -2936 649876 586860 649898
rect -1996 649874 -1396 649876
rect 804 649874 1404 649876
rect 36804 649874 37404 649876
rect 72804 649874 73404 649876
rect 108804 649874 109404 649876
rect 144804 649874 145404 649876
rect 180804 649874 181404 649876
rect 216804 649874 217404 649876
rect 252804 649874 253404 649876
rect 288804 649874 289404 649876
rect 324804 649874 325404 649876
rect 360804 649874 361404 649876
rect 396804 649874 397404 649876
rect 432804 649874 433404 649876
rect 468804 649874 469404 649876
rect 504804 649874 505404 649876
rect 540804 649874 541404 649876
rect 576804 649874 577404 649876
rect 585320 649874 585920 649876
rect -8576 643276 -7976 643278
rect 29604 643276 30204 643278
rect 65604 643276 66204 643278
rect 101604 643276 102204 643278
rect 137604 643276 138204 643278
rect 173604 643276 174204 643278
rect 209604 643276 210204 643278
rect 245604 643276 246204 643278
rect 281604 643276 282204 643278
rect 317604 643276 318204 643278
rect 353604 643276 354204 643278
rect 389604 643276 390204 643278
rect 425604 643276 426204 643278
rect 461604 643276 462204 643278
rect 497604 643276 498204 643278
rect 533604 643276 534204 643278
rect 569604 643276 570204 643278
rect 591900 643276 592500 643278
rect -8576 643254 592500 643276
rect -8576 643018 -8394 643254
rect -8158 643018 29786 643254
rect 30022 643018 65786 643254
rect 66022 643018 101786 643254
rect 102022 643018 137786 643254
rect 138022 643018 173786 643254
rect 174022 643018 209786 643254
rect 210022 643018 245786 643254
rect 246022 643018 281786 643254
rect 282022 643018 317786 643254
rect 318022 643018 353786 643254
rect 354022 643018 389786 643254
rect 390022 643018 425786 643254
rect 426022 643018 461786 643254
rect 462022 643018 497786 643254
rect 498022 643018 533786 643254
rect 534022 643018 569786 643254
rect 570022 643018 592082 643254
rect 592318 643018 592500 643254
rect -8576 642934 592500 643018
rect -8576 642698 -8394 642934
rect -8158 642698 29786 642934
rect 30022 642698 65786 642934
rect 66022 642698 101786 642934
rect 102022 642698 137786 642934
rect 138022 642698 173786 642934
rect 174022 642698 209786 642934
rect 210022 642698 245786 642934
rect 246022 642698 281786 642934
rect 282022 642698 317786 642934
rect 318022 642698 353786 642934
rect 354022 642698 389786 642934
rect 390022 642698 425786 642934
rect 426022 642698 461786 642934
rect 462022 642698 497786 642934
rect 498022 642698 533786 642934
rect 534022 642698 569786 642934
rect 570022 642698 592082 642934
rect 592318 642698 592500 642934
rect -8576 642676 592500 642698
rect -8576 642674 -7976 642676
rect 29604 642674 30204 642676
rect 65604 642674 66204 642676
rect 101604 642674 102204 642676
rect 137604 642674 138204 642676
rect 173604 642674 174204 642676
rect 209604 642674 210204 642676
rect 245604 642674 246204 642676
rect 281604 642674 282204 642676
rect 317604 642674 318204 642676
rect 353604 642674 354204 642676
rect 389604 642674 390204 642676
rect 425604 642674 426204 642676
rect 461604 642674 462204 642676
rect 497604 642674 498204 642676
rect 533604 642674 534204 642676
rect 569604 642674 570204 642676
rect 591900 642674 592500 642676
rect -6696 639676 -6096 639678
rect 26004 639676 26604 639678
rect 62004 639676 62604 639678
rect 98004 639676 98604 639678
rect 134004 639676 134604 639678
rect 170004 639676 170604 639678
rect 206004 639676 206604 639678
rect 242004 639676 242604 639678
rect 278004 639676 278604 639678
rect 314004 639676 314604 639678
rect 350004 639676 350604 639678
rect 386004 639676 386604 639678
rect 422004 639676 422604 639678
rect 458004 639676 458604 639678
rect 494004 639676 494604 639678
rect 530004 639676 530604 639678
rect 566004 639676 566604 639678
rect 590020 639676 590620 639678
rect -6696 639654 590620 639676
rect -6696 639418 -6514 639654
rect -6278 639418 26186 639654
rect 26422 639418 62186 639654
rect 62422 639418 98186 639654
rect 98422 639418 134186 639654
rect 134422 639418 170186 639654
rect 170422 639418 206186 639654
rect 206422 639418 242186 639654
rect 242422 639418 278186 639654
rect 278422 639418 314186 639654
rect 314422 639418 350186 639654
rect 350422 639418 386186 639654
rect 386422 639418 422186 639654
rect 422422 639418 458186 639654
rect 458422 639418 494186 639654
rect 494422 639418 530186 639654
rect 530422 639418 566186 639654
rect 566422 639418 590202 639654
rect 590438 639418 590620 639654
rect -6696 639334 590620 639418
rect -6696 639098 -6514 639334
rect -6278 639098 26186 639334
rect 26422 639098 62186 639334
rect 62422 639098 98186 639334
rect 98422 639098 134186 639334
rect 134422 639098 170186 639334
rect 170422 639098 206186 639334
rect 206422 639098 242186 639334
rect 242422 639098 278186 639334
rect 278422 639098 314186 639334
rect 314422 639098 350186 639334
rect 350422 639098 386186 639334
rect 386422 639098 422186 639334
rect 422422 639098 458186 639334
rect 458422 639098 494186 639334
rect 494422 639098 530186 639334
rect 530422 639098 566186 639334
rect 566422 639098 590202 639334
rect 590438 639098 590620 639334
rect -6696 639076 590620 639098
rect -6696 639074 -6096 639076
rect 26004 639074 26604 639076
rect 62004 639074 62604 639076
rect 98004 639074 98604 639076
rect 134004 639074 134604 639076
rect 170004 639074 170604 639076
rect 206004 639074 206604 639076
rect 242004 639074 242604 639076
rect 278004 639074 278604 639076
rect 314004 639074 314604 639076
rect 350004 639074 350604 639076
rect 386004 639074 386604 639076
rect 422004 639074 422604 639076
rect 458004 639074 458604 639076
rect 494004 639074 494604 639076
rect 530004 639074 530604 639076
rect 566004 639074 566604 639076
rect 590020 639074 590620 639076
rect -4816 636076 -4216 636078
rect 22404 636076 23004 636078
rect 58404 636076 59004 636078
rect 94404 636076 95004 636078
rect 130404 636076 131004 636078
rect 166404 636076 167004 636078
rect 202404 636076 203004 636078
rect 238404 636076 239004 636078
rect 274404 636076 275004 636078
rect 310404 636076 311004 636078
rect 346404 636076 347004 636078
rect 382404 636076 383004 636078
rect 418404 636076 419004 636078
rect 454404 636076 455004 636078
rect 490404 636076 491004 636078
rect 526404 636076 527004 636078
rect 562404 636076 563004 636078
rect 588140 636076 588740 636078
rect -4816 636054 588740 636076
rect -4816 635818 -4634 636054
rect -4398 635818 22586 636054
rect 22822 635818 58586 636054
rect 58822 635818 94586 636054
rect 94822 635818 130586 636054
rect 130822 635818 166586 636054
rect 166822 635818 202586 636054
rect 202822 635818 238586 636054
rect 238822 635818 274586 636054
rect 274822 635818 310586 636054
rect 310822 635818 346586 636054
rect 346822 635818 382586 636054
rect 382822 635818 418586 636054
rect 418822 635818 454586 636054
rect 454822 635818 490586 636054
rect 490822 635818 526586 636054
rect 526822 635818 562586 636054
rect 562822 635818 588322 636054
rect 588558 635818 588740 636054
rect -4816 635734 588740 635818
rect -4816 635498 -4634 635734
rect -4398 635498 22586 635734
rect 22822 635498 58586 635734
rect 58822 635498 94586 635734
rect 94822 635498 130586 635734
rect 130822 635498 166586 635734
rect 166822 635498 202586 635734
rect 202822 635498 238586 635734
rect 238822 635498 274586 635734
rect 274822 635498 310586 635734
rect 310822 635498 346586 635734
rect 346822 635498 382586 635734
rect 382822 635498 418586 635734
rect 418822 635498 454586 635734
rect 454822 635498 490586 635734
rect 490822 635498 526586 635734
rect 526822 635498 562586 635734
rect 562822 635498 588322 635734
rect 588558 635498 588740 635734
rect -4816 635476 588740 635498
rect -4816 635474 -4216 635476
rect 22404 635474 23004 635476
rect 58404 635474 59004 635476
rect 94404 635474 95004 635476
rect 130404 635474 131004 635476
rect 166404 635474 167004 635476
rect 202404 635474 203004 635476
rect 238404 635474 239004 635476
rect 274404 635474 275004 635476
rect 310404 635474 311004 635476
rect 346404 635474 347004 635476
rect 382404 635474 383004 635476
rect 418404 635474 419004 635476
rect 454404 635474 455004 635476
rect 490404 635474 491004 635476
rect 526404 635474 527004 635476
rect 562404 635474 563004 635476
rect 588140 635474 588740 635476
rect -2936 632476 -2336 632478
rect 18804 632476 19404 632478
rect 54804 632476 55404 632478
rect 90804 632476 91404 632478
rect 126804 632476 127404 632478
rect 162804 632476 163404 632478
rect 198804 632476 199404 632478
rect 234804 632476 235404 632478
rect 270804 632476 271404 632478
rect 306804 632476 307404 632478
rect 342804 632476 343404 632478
rect 378804 632476 379404 632478
rect 414804 632476 415404 632478
rect 450804 632476 451404 632478
rect 486804 632476 487404 632478
rect 522804 632476 523404 632478
rect 558804 632476 559404 632478
rect 586260 632476 586860 632478
rect -2936 632454 586860 632476
rect -2936 632218 -2754 632454
rect -2518 632218 18986 632454
rect 19222 632218 54986 632454
rect 55222 632218 90986 632454
rect 91222 632218 126986 632454
rect 127222 632218 162986 632454
rect 163222 632218 198986 632454
rect 199222 632218 234986 632454
rect 235222 632218 270986 632454
rect 271222 632218 306986 632454
rect 307222 632218 342986 632454
rect 343222 632218 378986 632454
rect 379222 632218 414986 632454
rect 415222 632218 450986 632454
rect 451222 632218 486986 632454
rect 487222 632218 522986 632454
rect 523222 632218 558986 632454
rect 559222 632218 586442 632454
rect 586678 632218 586860 632454
rect -2936 632134 586860 632218
rect -2936 631898 -2754 632134
rect -2518 631898 18986 632134
rect 19222 631898 54986 632134
rect 55222 631898 90986 632134
rect 91222 631898 126986 632134
rect 127222 631898 162986 632134
rect 163222 631898 198986 632134
rect 199222 631898 234986 632134
rect 235222 631898 270986 632134
rect 271222 631898 306986 632134
rect 307222 631898 342986 632134
rect 343222 631898 378986 632134
rect 379222 631898 414986 632134
rect 415222 631898 450986 632134
rect 451222 631898 486986 632134
rect 487222 631898 522986 632134
rect 523222 631898 558986 632134
rect 559222 631898 586442 632134
rect 586678 631898 586860 632134
rect -2936 631876 586860 631898
rect -2936 631874 -2336 631876
rect 18804 631874 19404 631876
rect 54804 631874 55404 631876
rect 90804 631874 91404 631876
rect 126804 631874 127404 631876
rect 162804 631874 163404 631876
rect 198804 631874 199404 631876
rect 234804 631874 235404 631876
rect 270804 631874 271404 631876
rect 306804 631874 307404 631876
rect 342804 631874 343404 631876
rect 378804 631874 379404 631876
rect 414804 631874 415404 631876
rect 450804 631874 451404 631876
rect 486804 631874 487404 631876
rect 522804 631874 523404 631876
rect 558804 631874 559404 631876
rect 586260 631874 586860 631876
rect -7636 625276 -7036 625278
rect 11604 625276 12204 625278
rect 47604 625276 48204 625278
rect 83604 625276 84204 625278
rect 119604 625276 120204 625278
rect 155604 625276 156204 625278
rect 191604 625276 192204 625278
rect 227604 625276 228204 625278
rect 263604 625276 264204 625278
rect 299604 625276 300204 625278
rect 335604 625276 336204 625278
rect 371604 625276 372204 625278
rect 407604 625276 408204 625278
rect 443604 625276 444204 625278
rect 479604 625276 480204 625278
rect 515604 625276 516204 625278
rect 551604 625276 552204 625278
rect 590960 625276 591560 625278
rect -8576 625254 592500 625276
rect -8576 625018 -7454 625254
rect -7218 625018 11786 625254
rect 12022 625018 47786 625254
rect 48022 625018 83786 625254
rect 84022 625018 119786 625254
rect 120022 625018 155786 625254
rect 156022 625018 191786 625254
rect 192022 625018 227786 625254
rect 228022 625018 263786 625254
rect 264022 625018 299786 625254
rect 300022 625018 335786 625254
rect 336022 625018 371786 625254
rect 372022 625018 407786 625254
rect 408022 625018 443786 625254
rect 444022 625018 479786 625254
rect 480022 625018 515786 625254
rect 516022 625018 551786 625254
rect 552022 625018 591142 625254
rect 591378 625018 592500 625254
rect -8576 624934 592500 625018
rect -8576 624698 -7454 624934
rect -7218 624698 11786 624934
rect 12022 624698 47786 624934
rect 48022 624698 83786 624934
rect 84022 624698 119786 624934
rect 120022 624698 155786 624934
rect 156022 624698 191786 624934
rect 192022 624698 227786 624934
rect 228022 624698 263786 624934
rect 264022 624698 299786 624934
rect 300022 624698 335786 624934
rect 336022 624698 371786 624934
rect 372022 624698 407786 624934
rect 408022 624698 443786 624934
rect 444022 624698 479786 624934
rect 480022 624698 515786 624934
rect 516022 624698 551786 624934
rect 552022 624698 591142 624934
rect 591378 624698 592500 624934
rect -8576 624676 592500 624698
rect -7636 624674 -7036 624676
rect 11604 624674 12204 624676
rect 47604 624674 48204 624676
rect 83604 624674 84204 624676
rect 119604 624674 120204 624676
rect 155604 624674 156204 624676
rect 191604 624674 192204 624676
rect 227604 624674 228204 624676
rect 263604 624674 264204 624676
rect 299604 624674 300204 624676
rect 335604 624674 336204 624676
rect 371604 624674 372204 624676
rect 407604 624674 408204 624676
rect 443604 624674 444204 624676
rect 479604 624674 480204 624676
rect 515604 624674 516204 624676
rect 551604 624674 552204 624676
rect 590960 624674 591560 624676
rect -5756 621676 -5156 621678
rect 8004 621676 8604 621678
rect 44004 621676 44604 621678
rect 80004 621676 80604 621678
rect 116004 621676 116604 621678
rect 152004 621676 152604 621678
rect 188004 621676 188604 621678
rect 224004 621676 224604 621678
rect 260004 621676 260604 621678
rect 296004 621676 296604 621678
rect 332004 621676 332604 621678
rect 368004 621676 368604 621678
rect 404004 621676 404604 621678
rect 440004 621676 440604 621678
rect 476004 621676 476604 621678
rect 512004 621676 512604 621678
rect 548004 621676 548604 621678
rect 589080 621676 589680 621678
rect -6696 621654 590620 621676
rect -6696 621418 -5574 621654
rect -5338 621418 8186 621654
rect 8422 621418 44186 621654
rect 44422 621418 80186 621654
rect 80422 621418 116186 621654
rect 116422 621418 152186 621654
rect 152422 621418 188186 621654
rect 188422 621418 224186 621654
rect 224422 621418 260186 621654
rect 260422 621418 296186 621654
rect 296422 621418 332186 621654
rect 332422 621418 368186 621654
rect 368422 621418 404186 621654
rect 404422 621418 440186 621654
rect 440422 621418 476186 621654
rect 476422 621418 512186 621654
rect 512422 621418 548186 621654
rect 548422 621418 589262 621654
rect 589498 621418 590620 621654
rect -6696 621334 590620 621418
rect -6696 621098 -5574 621334
rect -5338 621098 8186 621334
rect 8422 621098 44186 621334
rect 44422 621098 80186 621334
rect 80422 621098 116186 621334
rect 116422 621098 152186 621334
rect 152422 621098 188186 621334
rect 188422 621098 224186 621334
rect 224422 621098 260186 621334
rect 260422 621098 296186 621334
rect 296422 621098 332186 621334
rect 332422 621098 368186 621334
rect 368422 621098 404186 621334
rect 404422 621098 440186 621334
rect 440422 621098 476186 621334
rect 476422 621098 512186 621334
rect 512422 621098 548186 621334
rect 548422 621098 589262 621334
rect 589498 621098 590620 621334
rect -6696 621076 590620 621098
rect -5756 621074 -5156 621076
rect 8004 621074 8604 621076
rect 44004 621074 44604 621076
rect 80004 621074 80604 621076
rect 116004 621074 116604 621076
rect 152004 621074 152604 621076
rect 188004 621074 188604 621076
rect 224004 621074 224604 621076
rect 260004 621074 260604 621076
rect 296004 621074 296604 621076
rect 332004 621074 332604 621076
rect 368004 621074 368604 621076
rect 404004 621074 404604 621076
rect 440004 621074 440604 621076
rect 476004 621074 476604 621076
rect 512004 621074 512604 621076
rect 548004 621074 548604 621076
rect 589080 621074 589680 621076
rect -3876 618076 -3276 618078
rect 4404 618076 5004 618078
rect 40404 618076 41004 618078
rect 76404 618076 77004 618078
rect 112404 618076 113004 618078
rect 148404 618076 149004 618078
rect 184404 618076 185004 618078
rect 220404 618076 221004 618078
rect 256404 618076 257004 618078
rect 292404 618076 293004 618078
rect 328404 618076 329004 618078
rect 364404 618076 365004 618078
rect 400404 618076 401004 618078
rect 436404 618076 437004 618078
rect 472404 618076 473004 618078
rect 508404 618076 509004 618078
rect 544404 618076 545004 618078
rect 580404 618076 581004 618078
rect 587200 618076 587800 618078
rect -4816 618054 588740 618076
rect -4816 617818 -3694 618054
rect -3458 617818 4586 618054
rect 4822 617818 40586 618054
rect 40822 617818 76586 618054
rect 76822 617818 112586 618054
rect 112822 617818 148586 618054
rect 148822 617818 184586 618054
rect 184822 617818 220586 618054
rect 220822 617818 256586 618054
rect 256822 617818 292586 618054
rect 292822 617818 328586 618054
rect 328822 617818 364586 618054
rect 364822 617818 400586 618054
rect 400822 617818 436586 618054
rect 436822 617818 472586 618054
rect 472822 617818 508586 618054
rect 508822 617818 544586 618054
rect 544822 617818 580586 618054
rect 580822 617818 587382 618054
rect 587618 617818 588740 618054
rect -4816 617734 588740 617818
rect -4816 617498 -3694 617734
rect -3458 617498 4586 617734
rect 4822 617498 40586 617734
rect 40822 617498 76586 617734
rect 76822 617498 112586 617734
rect 112822 617498 148586 617734
rect 148822 617498 184586 617734
rect 184822 617498 220586 617734
rect 220822 617498 256586 617734
rect 256822 617498 292586 617734
rect 292822 617498 328586 617734
rect 328822 617498 364586 617734
rect 364822 617498 400586 617734
rect 400822 617498 436586 617734
rect 436822 617498 472586 617734
rect 472822 617498 508586 617734
rect 508822 617498 544586 617734
rect 544822 617498 580586 617734
rect 580822 617498 587382 617734
rect 587618 617498 588740 617734
rect -4816 617476 588740 617498
rect -3876 617474 -3276 617476
rect 4404 617474 5004 617476
rect 40404 617474 41004 617476
rect 76404 617474 77004 617476
rect 112404 617474 113004 617476
rect 148404 617474 149004 617476
rect 184404 617474 185004 617476
rect 220404 617474 221004 617476
rect 256404 617474 257004 617476
rect 292404 617474 293004 617476
rect 328404 617474 329004 617476
rect 364404 617474 365004 617476
rect 400404 617474 401004 617476
rect 436404 617474 437004 617476
rect 472404 617474 473004 617476
rect 508404 617474 509004 617476
rect 544404 617474 545004 617476
rect 580404 617474 581004 617476
rect 587200 617474 587800 617476
rect -1996 614476 -1396 614478
rect 804 614476 1404 614478
rect 36804 614476 37404 614478
rect 72804 614476 73404 614478
rect 108804 614476 109404 614478
rect 144804 614476 145404 614478
rect 180804 614476 181404 614478
rect 216804 614476 217404 614478
rect 252804 614476 253404 614478
rect 288804 614476 289404 614478
rect 324804 614476 325404 614478
rect 360804 614476 361404 614478
rect 396804 614476 397404 614478
rect 432804 614476 433404 614478
rect 468804 614476 469404 614478
rect 504804 614476 505404 614478
rect 540804 614476 541404 614478
rect 576804 614476 577404 614478
rect 585320 614476 585920 614478
rect -2936 614454 586860 614476
rect -2936 614218 -1814 614454
rect -1578 614218 986 614454
rect 1222 614218 36986 614454
rect 37222 614218 72986 614454
rect 73222 614218 108986 614454
rect 109222 614218 144986 614454
rect 145222 614218 180986 614454
rect 181222 614218 216986 614454
rect 217222 614218 252986 614454
rect 253222 614218 288986 614454
rect 289222 614218 324986 614454
rect 325222 614218 360986 614454
rect 361222 614218 396986 614454
rect 397222 614218 432986 614454
rect 433222 614218 468986 614454
rect 469222 614218 504986 614454
rect 505222 614218 540986 614454
rect 541222 614218 576986 614454
rect 577222 614218 585502 614454
rect 585738 614218 586860 614454
rect -2936 614134 586860 614218
rect -2936 613898 -1814 614134
rect -1578 613898 986 614134
rect 1222 613898 36986 614134
rect 37222 613898 72986 614134
rect 73222 613898 108986 614134
rect 109222 613898 144986 614134
rect 145222 613898 180986 614134
rect 181222 613898 216986 614134
rect 217222 613898 252986 614134
rect 253222 613898 288986 614134
rect 289222 613898 324986 614134
rect 325222 613898 360986 614134
rect 361222 613898 396986 614134
rect 397222 613898 432986 614134
rect 433222 613898 468986 614134
rect 469222 613898 504986 614134
rect 505222 613898 540986 614134
rect 541222 613898 576986 614134
rect 577222 613898 585502 614134
rect 585738 613898 586860 614134
rect -2936 613876 586860 613898
rect -1996 613874 -1396 613876
rect 804 613874 1404 613876
rect 36804 613874 37404 613876
rect 72804 613874 73404 613876
rect 108804 613874 109404 613876
rect 144804 613874 145404 613876
rect 180804 613874 181404 613876
rect 216804 613874 217404 613876
rect 252804 613874 253404 613876
rect 288804 613874 289404 613876
rect 324804 613874 325404 613876
rect 360804 613874 361404 613876
rect 396804 613874 397404 613876
rect 432804 613874 433404 613876
rect 468804 613874 469404 613876
rect 504804 613874 505404 613876
rect 540804 613874 541404 613876
rect 576804 613874 577404 613876
rect 585320 613874 585920 613876
rect -8576 607276 -7976 607278
rect 29604 607276 30204 607278
rect 65604 607276 66204 607278
rect 101604 607276 102204 607278
rect 137604 607276 138204 607278
rect 173604 607276 174204 607278
rect 209604 607276 210204 607278
rect 245604 607276 246204 607278
rect 281604 607276 282204 607278
rect 317604 607276 318204 607278
rect 353604 607276 354204 607278
rect 389604 607276 390204 607278
rect 425604 607276 426204 607278
rect 461604 607276 462204 607278
rect 497604 607276 498204 607278
rect 533604 607276 534204 607278
rect 569604 607276 570204 607278
rect 591900 607276 592500 607278
rect -8576 607254 592500 607276
rect -8576 607018 -8394 607254
rect -8158 607018 29786 607254
rect 30022 607018 65786 607254
rect 66022 607018 101786 607254
rect 102022 607018 137786 607254
rect 138022 607018 173786 607254
rect 174022 607018 209786 607254
rect 210022 607018 245786 607254
rect 246022 607018 281786 607254
rect 282022 607018 317786 607254
rect 318022 607018 353786 607254
rect 354022 607018 389786 607254
rect 390022 607018 425786 607254
rect 426022 607018 461786 607254
rect 462022 607018 497786 607254
rect 498022 607018 533786 607254
rect 534022 607018 569786 607254
rect 570022 607018 592082 607254
rect 592318 607018 592500 607254
rect -8576 606934 592500 607018
rect -8576 606698 -8394 606934
rect -8158 606698 29786 606934
rect 30022 606698 65786 606934
rect 66022 606698 101786 606934
rect 102022 606698 137786 606934
rect 138022 606698 173786 606934
rect 174022 606698 209786 606934
rect 210022 606698 245786 606934
rect 246022 606698 281786 606934
rect 282022 606698 317786 606934
rect 318022 606698 353786 606934
rect 354022 606698 389786 606934
rect 390022 606698 425786 606934
rect 426022 606698 461786 606934
rect 462022 606698 497786 606934
rect 498022 606698 533786 606934
rect 534022 606698 569786 606934
rect 570022 606698 592082 606934
rect 592318 606698 592500 606934
rect -8576 606676 592500 606698
rect -8576 606674 -7976 606676
rect 29604 606674 30204 606676
rect 65604 606674 66204 606676
rect 101604 606674 102204 606676
rect 137604 606674 138204 606676
rect 173604 606674 174204 606676
rect 209604 606674 210204 606676
rect 245604 606674 246204 606676
rect 281604 606674 282204 606676
rect 317604 606674 318204 606676
rect 353604 606674 354204 606676
rect 389604 606674 390204 606676
rect 425604 606674 426204 606676
rect 461604 606674 462204 606676
rect 497604 606674 498204 606676
rect 533604 606674 534204 606676
rect 569604 606674 570204 606676
rect 591900 606674 592500 606676
rect -6696 603676 -6096 603678
rect 26004 603676 26604 603678
rect 62004 603676 62604 603678
rect 98004 603676 98604 603678
rect 134004 603676 134604 603678
rect 170004 603676 170604 603678
rect 206004 603676 206604 603678
rect 242004 603676 242604 603678
rect 278004 603676 278604 603678
rect 314004 603676 314604 603678
rect 350004 603676 350604 603678
rect 386004 603676 386604 603678
rect 422004 603676 422604 603678
rect 458004 603676 458604 603678
rect 494004 603676 494604 603678
rect 530004 603676 530604 603678
rect 566004 603676 566604 603678
rect 590020 603676 590620 603678
rect -6696 603654 590620 603676
rect -6696 603418 -6514 603654
rect -6278 603418 26186 603654
rect 26422 603418 62186 603654
rect 62422 603418 98186 603654
rect 98422 603418 134186 603654
rect 134422 603418 170186 603654
rect 170422 603418 206186 603654
rect 206422 603418 242186 603654
rect 242422 603418 278186 603654
rect 278422 603418 314186 603654
rect 314422 603418 350186 603654
rect 350422 603418 386186 603654
rect 386422 603418 422186 603654
rect 422422 603418 458186 603654
rect 458422 603418 494186 603654
rect 494422 603418 530186 603654
rect 530422 603418 566186 603654
rect 566422 603418 590202 603654
rect 590438 603418 590620 603654
rect -6696 603334 590620 603418
rect -6696 603098 -6514 603334
rect -6278 603098 26186 603334
rect 26422 603098 62186 603334
rect 62422 603098 98186 603334
rect 98422 603098 134186 603334
rect 134422 603098 170186 603334
rect 170422 603098 206186 603334
rect 206422 603098 242186 603334
rect 242422 603098 278186 603334
rect 278422 603098 314186 603334
rect 314422 603098 350186 603334
rect 350422 603098 386186 603334
rect 386422 603098 422186 603334
rect 422422 603098 458186 603334
rect 458422 603098 494186 603334
rect 494422 603098 530186 603334
rect 530422 603098 566186 603334
rect 566422 603098 590202 603334
rect 590438 603098 590620 603334
rect -6696 603076 590620 603098
rect -6696 603074 -6096 603076
rect 26004 603074 26604 603076
rect 62004 603074 62604 603076
rect 98004 603074 98604 603076
rect 134004 603074 134604 603076
rect 170004 603074 170604 603076
rect 206004 603074 206604 603076
rect 242004 603074 242604 603076
rect 278004 603074 278604 603076
rect 314004 603074 314604 603076
rect 350004 603074 350604 603076
rect 386004 603074 386604 603076
rect 422004 603074 422604 603076
rect 458004 603074 458604 603076
rect 494004 603074 494604 603076
rect 530004 603074 530604 603076
rect 566004 603074 566604 603076
rect 590020 603074 590620 603076
rect -4816 600076 -4216 600078
rect 22404 600076 23004 600078
rect 58404 600076 59004 600078
rect 94404 600076 95004 600078
rect 130404 600076 131004 600078
rect 166404 600076 167004 600078
rect 202404 600076 203004 600078
rect 238404 600076 239004 600078
rect 274404 600076 275004 600078
rect 310404 600076 311004 600078
rect 346404 600076 347004 600078
rect 382404 600076 383004 600078
rect 418404 600076 419004 600078
rect 454404 600076 455004 600078
rect 490404 600076 491004 600078
rect 526404 600076 527004 600078
rect 562404 600076 563004 600078
rect 588140 600076 588740 600078
rect -4816 600054 588740 600076
rect -4816 599818 -4634 600054
rect -4398 599818 22586 600054
rect 22822 599818 58586 600054
rect 58822 599818 94586 600054
rect 94822 599818 130586 600054
rect 130822 599818 166586 600054
rect 166822 599818 202586 600054
rect 202822 599818 238586 600054
rect 238822 599818 274586 600054
rect 274822 599818 310586 600054
rect 310822 599818 346586 600054
rect 346822 599818 382586 600054
rect 382822 599818 418586 600054
rect 418822 599818 454586 600054
rect 454822 599818 490586 600054
rect 490822 599818 526586 600054
rect 526822 599818 562586 600054
rect 562822 599818 588322 600054
rect 588558 599818 588740 600054
rect -4816 599734 588740 599818
rect -4816 599498 -4634 599734
rect -4398 599498 22586 599734
rect 22822 599498 58586 599734
rect 58822 599498 94586 599734
rect 94822 599498 130586 599734
rect 130822 599498 166586 599734
rect 166822 599498 202586 599734
rect 202822 599498 238586 599734
rect 238822 599498 274586 599734
rect 274822 599498 310586 599734
rect 310822 599498 346586 599734
rect 346822 599498 382586 599734
rect 382822 599498 418586 599734
rect 418822 599498 454586 599734
rect 454822 599498 490586 599734
rect 490822 599498 526586 599734
rect 526822 599498 562586 599734
rect 562822 599498 588322 599734
rect 588558 599498 588740 599734
rect -4816 599476 588740 599498
rect -4816 599474 -4216 599476
rect 22404 599474 23004 599476
rect 58404 599474 59004 599476
rect 94404 599474 95004 599476
rect 130404 599474 131004 599476
rect 166404 599474 167004 599476
rect 202404 599474 203004 599476
rect 238404 599474 239004 599476
rect 274404 599474 275004 599476
rect 310404 599474 311004 599476
rect 346404 599474 347004 599476
rect 382404 599474 383004 599476
rect 418404 599474 419004 599476
rect 454404 599474 455004 599476
rect 490404 599474 491004 599476
rect 526404 599474 527004 599476
rect 562404 599474 563004 599476
rect 588140 599474 588740 599476
rect -2936 596476 -2336 596478
rect 18804 596476 19404 596478
rect 54804 596476 55404 596478
rect 90804 596476 91404 596478
rect 126804 596476 127404 596478
rect 162804 596476 163404 596478
rect 198804 596476 199404 596478
rect 234804 596476 235404 596478
rect 270804 596476 271404 596478
rect 306804 596476 307404 596478
rect 342804 596476 343404 596478
rect 378804 596476 379404 596478
rect 414804 596476 415404 596478
rect 450804 596476 451404 596478
rect 486804 596476 487404 596478
rect 522804 596476 523404 596478
rect 558804 596476 559404 596478
rect 586260 596476 586860 596478
rect -2936 596454 586860 596476
rect -2936 596218 -2754 596454
rect -2518 596218 18986 596454
rect 19222 596218 54986 596454
rect 55222 596218 90986 596454
rect 91222 596218 126986 596454
rect 127222 596218 162986 596454
rect 163222 596218 198986 596454
rect 199222 596218 234986 596454
rect 235222 596218 270986 596454
rect 271222 596218 306986 596454
rect 307222 596218 342986 596454
rect 343222 596218 378986 596454
rect 379222 596218 414986 596454
rect 415222 596218 450986 596454
rect 451222 596218 486986 596454
rect 487222 596218 522986 596454
rect 523222 596218 558986 596454
rect 559222 596218 586442 596454
rect 586678 596218 586860 596454
rect -2936 596134 586860 596218
rect -2936 595898 -2754 596134
rect -2518 595898 18986 596134
rect 19222 595898 54986 596134
rect 55222 595898 90986 596134
rect 91222 595898 126986 596134
rect 127222 595898 162986 596134
rect 163222 595898 198986 596134
rect 199222 595898 234986 596134
rect 235222 595898 270986 596134
rect 271222 595898 306986 596134
rect 307222 595898 342986 596134
rect 343222 595898 378986 596134
rect 379222 595898 414986 596134
rect 415222 595898 450986 596134
rect 451222 595898 486986 596134
rect 487222 595898 522986 596134
rect 523222 595898 558986 596134
rect 559222 595898 586442 596134
rect 586678 595898 586860 596134
rect -2936 595876 586860 595898
rect -2936 595874 -2336 595876
rect 18804 595874 19404 595876
rect 54804 595874 55404 595876
rect 90804 595874 91404 595876
rect 126804 595874 127404 595876
rect 162804 595874 163404 595876
rect 198804 595874 199404 595876
rect 234804 595874 235404 595876
rect 270804 595874 271404 595876
rect 306804 595874 307404 595876
rect 342804 595874 343404 595876
rect 378804 595874 379404 595876
rect 414804 595874 415404 595876
rect 450804 595874 451404 595876
rect 486804 595874 487404 595876
rect 522804 595874 523404 595876
rect 558804 595874 559404 595876
rect 586260 595874 586860 595876
rect -7636 589276 -7036 589278
rect 11604 589276 12204 589278
rect 47604 589276 48204 589278
rect 83604 589276 84204 589278
rect 119604 589276 120204 589278
rect 155604 589276 156204 589278
rect 191604 589276 192204 589278
rect 227604 589276 228204 589278
rect 263604 589276 264204 589278
rect 299604 589276 300204 589278
rect 335604 589276 336204 589278
rect 371604 589276 372204 589278
rect 407604 589276 408204 589278
rect 443604 589276 444204 589278
rect 479604 589276 480204 589278
rect 515604 589276 516204 589278
rect 551604 589276 552204 589278
rect 590960 589276 591560 589278
rect -8576 589254 592500 589276
rect -8576 589018 -7454 589254
rect -7218 589018 11786 589254
rect 12022 589018 47786 589254
rect 48022 589018 83786 589254
rect 84022 589018 119786 589254
rect 120022 589018 155786 589254
rect 156022 589018 191786 589254
rect 192022 589018 227786 589254
rect 228022 589018 263786 589254
rect 264022 589018 299786 589254
rect 300022 589018 335786 589254
rect 336022 589018 371786 589254
rect 372022 589018 407786 589254
rect 408022 589018 443786 589254
rect 444022 589018 479786 589254
rect 480022 589018 515786 589254
rect 516022 589018 551786 589254
rect 552022 589018 591142 589254
rect 591378 589018 592500 589254
rect -8576 588934 592500 589018
rect -8576 588698 -7454 588934
rect -7218 588698 11786 588934
rect 12022 588698 47786 588934
rect 48022 588698 83786 588934
rect 84022 588698 119786 588934
rect 120022 588698 155786 588934
rect 156022 588698 191786 588934
rect 192022 588698 227786 588934
rect 228022 588698 263786 588934
rect 264022 588698 299786 588934
rect 300022 588698 335786 588934
rect 336022 588698 371786 588934
rect 372022 588698 407786 588934
rect 408022 588698 443786 588934
rect 444022 588698 479786 588934
rect 480022 588698 515786 588934
rect 516022 588698 551786 588934
rect 552022 588698 591142 588934
rect 591378 588698 592500 588934
rect -8576 588676 592500 588698
rect -7636 588674 -7036 588676
rect 11604 588674 12204 588676
rect 47604 588674 48204 588676
rect 83604 588674 84204 588676
rect 119604 588674 120204 588676
rect 155604 588674 156204 588676
rect 191604 588674 192204 588676
rect 227604 588674 228204 588676
rect 263604 588674 264204 588676
rect 299604 588674 300204 588676
rect 335604 588674 336204 588676
rect 371604 588674 372204 588676
rect 407604 588674 408204 588676
rect 443604 588674 444204 588676
rect 479604 588674 480204 588676
rect 515604 588674 516204 588676
rect 551604 588674 552204 588676
rect 590960 588674 591560 588676
rect -5756 585676 -5156 585678
rect 8004 585676 8604 585678
rect 44004 585676 44604 585678
rect 80004 585676 80604 585678
rect 116004 585676 116604 585678
rect 152004 585676 152604 585678
rect 188004 585676 188604 585678
rect 224004 585676 224604 585678
rect 260004 585676 260604 585678
rect 296004 585676 296604 585678
rect 332004 585676 332604 585678
rect 368004 585676 368604 585678
rect 404004 585676 404604 585678
rect 440004 585676 440604 585678
rect 476004 585676 476604 585678
rect 512004 585676 512604 585678
rect 548004 585676 548604 585678
rect 589080 585676 589680 585678
rect -6696 585654 590620 585676
rect -6696 585418 -5574 585654
rect -5338 585418 8186 585654
rect 8422 585418 44186 585654
rect 44422 585418 80186 585654
rect 80422 585418 116186 585654
rect 116422 585418 152186 585654
rect 152422 585418 188186 585654
rect 188422 585418 224186 585654
rect 224422 585418 260186 585654
rect 260422 585418 296186 585654
rect 296422 585418 332186 585654
rect 332422 585418 368186 585654
rect 368422 585418 404186 585654
rect 404422 585418 440186 585654
rect 440422 585418 476186 585654
rect 476422 585418 512186 585654
rect 512422 585418 548186 585654
rect 548422 585418 589262 585654
rect 589498 585418 590620 585654
rect -6696 585334 590620 585418
rect -6696 585098 -5574 585334
rect -5338 585098 8186 585334
rect 8422 585098 44186 585334
rect 44422 585098 80186 585334
rect 80422 585098 116186 585334
rect 116422 585098 152186 585334
rect 152422 585098 188186 585334
rect 188422 585098 224186 585334
rect 224422 585098 260186 585334
rect 260422 585098 296186 585334
rect 296422 585098 332186 585334
rect 332422 585098 368186 585334
rect 368422 585098 404186 585334
rect 404422 585098 440186 585334
rect 440422 585098 476186 585334
rect 476422 585098 512186 585334
rect 512422 585098 548186 585334
rect 548422 585098 589262 585334
rect 589498 585098 590620 585334
rect -6696 585076 590620 585098
rect -5756 585074 -5156 585076
rect 8004 585074 8604 585076
rect 44004 585074 44604 585076
rect 80004 585074 80604 585076
rect 116004 585074 116604 585076
rect 152004 585074 152604 585076
rect 188004 585074 188604 585076
rect 224004 585074 224604 585076
rect 260004 585074 260604 585076
rect 296004 585074 296604 585076
rect 332004 585074 332604 585076
rect 368004 585074 368604 585076
rect 404004 585074 404604 585076
rect 440004 585074 440604 585076
rect 476004 585074 476604 585076
rect 512004 585074 512604 585076
rect 548004 585074 548604 585076
rect 589080 585074 589680 585076
rect -3876 582076 -3276 582078
rect 4404 582076 5004 582078
rect 40404 582076 41004 582078
rect 76404 582076 77004 582078
rect 112404 582076 113004 582078
rect 148404 582076 149004 582078
rect 184404 582076 185004 582078
rect 220404 582076 221004 582078
rect 256404 582076 257004 582078
rect 292404 582076 293004 582078
rect 328404 582076 329004 582078
rect 364404 582076 365004 582078
rect 400404 582076 401004 582078
rect 436404 582076 437004 582078
rect 472404 582076 473004 582078
rect 508404 582076 509004 582078
rect 544404 582076 545004 582078
rect 580404 582076 581004 582078
rect 587200 582076 587800 582078
rect -4816 582054 588740 582076
rect -4816 581818 -3694 582054
rect -3458 581818 4586 582054
rect 4822 581818 40586 582054
rect 40822 581818 76586 582054
rect 76822 581818 112586 582054
rect 112822 581818 148586 582054
rect 148822 581818 184586 582054
rect 184822 581818 220586 582054
rect 220822 581818 256586 582054
rect 256822 581818 292586 582054
rect 292822 581818 328586 582054
rect 328822 581818 364586 582054
rect 364822 581818 400586 582054
rect 400822 581818 436586 582054
rect 436822 581818 472586 582054
rect 472822 581818 508586 582054
rect 508822 581818 544586 582054
rect 544822 581818 580586 582054
rect 580822 581818 587382 582054
rect 587618 581818 588740 582054
rect -4816 581734 588740 581818
rect -4816 581498 -3694 581734
rect -3458 581498 4586 581734
rect 4822 581498 40586 581734
rect 40822 581498 76586 581734
rect 76822 581498 112586 581734
rect 112822 581498 148586 581734
rect 148822 581498 184586 581734
rect 184822 581498 220586 581734
rect 220822 581498 256586 581734
rect 256822 581498 292586 581734
rect 292822 581498 328586 581734
rect 328822 581498 364586 581734
rect 364822 581498 400586 581734
rect 400822 581498 436586 581734
rect 436822 581498 472586 581734
rect 472822 581498 508586 581734
rect 508822 581498 544586 581734
rect 544822 581498 580586 581734
rect 580822 581498 587382 581734
rect 587618 581498 588740 581734
rect -4816 581476 588740 581498
rect -3876 581474 -3276 581476
rect 4404 581474 5004 581476
rect 40404 581474 41004 581476
rect 76404 581474 77004 581476
rect 112404 581474 113004 581476
rect 148404 581474 149004 581476
rect 184404 581474 185004 581476
rect 220404 581474 221004 581476
rect 256404 581474 257004 581476
rect 292404 581474 293004 581476
rect 328404 581474 329004 581476
rect 364404 581474 365004 581476
rect 400404 581474 401004 581476
rect 436404 581474 437004 581476
rect 472404 581474 473004 581476
rect 508404 581474 509004 581476
rect 544404 581474 545004 581476
rect 580404 581474 581004 581476
rect 587200 581474 587800 581476
rect -1996 578476 -1396 578478
rect 804 578476 1404 578478
rect 36804 578476 37404 578478
rect 72804 578476 73404 578478
rect 108804 578476 109404 578478
rect 144804 578476 145404 578478
rect 180804 578476 181404 578478
rect 216804 578476 217404 578478
rect 252804 578476 253404 578478
rect 288804 578476 289404 578478
rect 324804 578476 325404 578478
rect 360804 578476 361404 578478
rect 396804 578476 397404 578478
rect 432804 578476 433404 578478
rect 468804 578476 469404 578478
rect 504804 578476 505404 578478
rect 540804 578476 541404 578478
rect 576804 578476 577404 578478
rect 585320 578476 585920 578478
rect -2936 578454 586860 578476
rect -2936 578218 -1814 578454
rect -1578 578218 986 578454
rect 1222 578218 36986 578454
rect 37222 578218 72986 578454
rect 73222 578218 108986 578454
rect 109222 578218 144986 578454
rect 145222 578218 180986 578454
rect 181222 578218 216986 578454
rect 217222 578218 252986 578454
rect 253222 578218 288986 578454
rect 289222 578218 324986 578454
rect 325222 578218 360986 578454
rect 361222 578218 396986 578454
rect 397222 578218 432986 578454
rect 433222 578218 468986 578454
rect 469222 578218 504986 578454
rect 505222 578218 540986 578454
rect 541222 578218 576986 578454
rect 577222 578218 585502 578454
rect 585738 578218 586860 578454
rect -2936 578134 586860 578218
rect -2936 577898 -1814 578134
rect -1578 577898 986 578134
rect 1222 577898 36986 578134
rect 37222 577898 72986 578134
rect 73222 577898 108986 578134
rect 109222 577898 144986 578134
rect 145222 577898 180986 578134
rect 181222 577898 216986 578134
rect 217222 577898 252986 578134
rect 253222 577898 288986 578134
rect 289222 577898 324986 578134
rect 325222 577898 360986 578134
rect 361222 577898 396986 578134
rect 397222 577898 432986 578134
rect 433222 577898 468986 578134
rect 469222 577898 504986 578134
rect 505222 577898 540986 578134
rect 541222 577898 576986 578134
rect 577222 577898 585502 578134
rect 585738 577898 586860 578134
rect -2936 577876 586860 577898
rect -1996 577874 -1396 577876
rect 804 577874 1404 577876
rect 36804 577874 37404 577876
rect 72804 577874 73404 577876
rect 108804 577874 109404 577876
rect 144804 577874 145404 577876
rect 180804 577874 181404 577876
rect 216804 577874 217404 577876
rect 252804 577874 253404 577876
rect 288804 577874 289404 577876
rect 324804 577874 325404 577876
rect 360804 577874 361404 577876
rect 396804 577874 397404 577876
rect 432804 577874 433404 577876
rect 468804 577874 469404 577876
rect 504804 577874 505404 577876
rect 540804 577874 541404 577876
rect 576804 577874 577404 577876
rect 585320 577874 585920 577876
rect -8576 571276 -7976 571278
rect 29604 571276 30204 571278
rect 65604 571276 66204 571278
rect 101604 571276 102204 571278
rect 137604 571276 138204 571278
rect 173604 571276 174204 571278
rect 209604 571276 210204 571278
rect 245604 571276 246204 571278
rect 281604 571276 282204 571278
rect 317604 571276 318204 571278
rect 353604 571276 354204 571278
rect 389604 571276 390204 571278
rect 425604 571276 426204 571278
rect 461604 571276 462204 571278
rect 497604 571276 498204 571278
rect 533604 571276 534204 571278
rect 569604 571276 570204 571278
rect 591900 571276 592500 571278
rect -8576 571254 592500 571276
rect -8576 571018 -8394 571254
rect -8158 571018 29786 571254
rect 30022 571018 65786 571254
rect 66022 571018 101786 571254
rect 102022 571018 137786 571254
rect 138022 571018 173786 571254
rect 174022 571018 209786 571254
rect 210022 571018 245786 571254
rect 246022 571018 281786 571254
rect 282022 571018 317786 571254
rect 318022 571018 353786 571254
rect 354022 571018 389786 571254
rect 390022 571018 425786 571254
rect 426022 571018 461786 571254
rect 462022 571018 497786 571254
rect 498022 571018 533786 571254
rect 534022 571018 569786 571254
rect 570022 571018 592082 571254
rect 592318 571018 592500 571254
rect -8576 570934 592500 571018
rect -8576 570698 -8394 570934
rect -8158 570698 29786 570934
rect 30022 570698 65786 570934
rect 66022 570698 101786 570934
rect 102022 570698 137786 570934
rect 138022 570698 173786 570934
rect 174022 570698 209786 570934
rect 210022 570698 245786 570934
rect 246022 570698 281786 570934
rect 282022 570698 317786 570934
rect 318022 570698 353786 570934
rect 354022 570698 389786 570934
rect 390022 570698 425786 570934
rect 426022 570698 461786 570934
rect 462022 570698 497786 570934
rect 498022 570698 533786 570934
rect 534022 570698 569786 570934
rect 570022 570698 592082 570934
rect 592318 570698 592500 570934
rect -8576 570676 592500 570698
rect -8576 570674 -7976 570676
rect 29604 570674 30204 570676
rect 65604 570674 66204 570676
rect 101604 570674 102204 570676
rect 137604 570674 138204 570676
rect 173604 570674 174204 570676
rect 209604 570674 210204 570676
rect 245604 570674 246204 570676
rect 281604 570674 282204 570676
rect 317604 570674 318204 570676
rect 353604 570674 354204 570676
rect 389604 570674 390204 570676
rect 425604 570674 426204 570676
rect 461604 570674 462204 570676
rect 497604 570674 498204 570676
rect 533604 570674 534204 570676
rect 569604 570674 570204 570676
rect 591900 570674 592500 570676
rect -6696 567676 -6096 567678
rect 26004 567676 26604 567678
rect 62004 567676 62604 567678
rect 98004 567676 98604 567678
rect 134004 567676 134604 567678
rect 170004 567676 170604 567678
rect 206004 567676 206604 567678
rect 242004 567676 242604 567678
rect 278004 567676 278604 567678
rect 314004 567676 314604 567678
rect 350004 567676 350604 567678
rect 386004 567676 386604 567678
rect 422004 567676 422604 567678
rect 458004 567676 458604 567678
rect 494004 567676 494604 567678
rect 530004 567676 530604 567678
rect 566004 567676 566604 567678
rect 590020 567676 590620 567678
rect -6696 567654 590620 567676
rect -6696 567418 -6514 567654
rect -6278 567418 26186 567654
rect 26422 567418 62186 567654
rect 62422 567418 98186 567654
rect 98422 567418 134186 567654
rect 134422 567418 170186 567654
rect 170422 567418 206186 567654
rect 206422 567418 242186 567654
rect 242422 567418 278186 567654
rect 278422 567418 314186 567654
rect 314422 567418 350186 567654
rect 350422 567418 386186 567654
rect 386422 567418 422186 567654
rect 422422 567418 458186 567654
rect 458422 567418 494186 567654
rect 494422 567418 530186 567654
rect 530422 567418 566186 567654
rect 566422 567418 590202 567654
rect 590438 567418 590620 567654
rect -6696 567334 590620 567418
rect -6696 567098 -6514 567334
rect -6278 567098 26186 567334
rect 26422 567098 62186 567334
rect 62422 567098 98186 567334
rect 98422 567098 134186 567334
rect 134422 567098 170186 567334
rect 170422 567098 206186 567334
rect 206422 567098 242186 567334
rect 242422 567098 278186 567334
rect 278422 567098 314186 567334
rect 314422 567098 350186 567334
rect 350422 567098 386186 567334
rect 386422 567098 422186 567334
rect 422422 567098 458186 567334
rect 458422 567098 494186 567334
rect 494422 567098 530186 567334
rect 530422 567098 566186 567334
rect 566422 567098 590202 567334
rect 590438 567098 590620 567334
rect -6696 567076 590620 567098
rect -6696 567074 -6096 567076
rect 26004 567074 26604 567076
rect 62004 567074 62604 567076
rect 98004 567074 98604 567076
rect 134004 567074 134604 567076
rect 170004 567074 170604 567076
rect 206004 567074 206604 567076
rect 242004 567074 242604 567076
rect 278004 567074 278604 567076
rect 314004 567074 314604 567076
rect 350004 567074 350604 567076
rect 386004 567074 386604 567076
rect 422004 567074 422604 567076
rect 458004 567074 458604 567076
rect 494004 567074 494604 567076
rect 530004 567074 530604 567076
rect 566004 567074 566604 567076
rect 590020 567074 590620 567076
rect -4816 564076 -4216 564078
rect 22404 564076 23004 564078
rect 58404 564076 59004 564078
rect 94404 564076 95004 564078
rect 130404 564076 131004 564078
rect 166404 564076 167004 564078
rect 202404 564076 203004 564078
rect 238404 564076 239004 564078
rect 274404 564076 275004 564078
rect 310404 564076 311004 564078
rect 346404 564076 347004 564078
rect 382404 564076 383004 564078
rect 418404 564076 419004 564078
rect 454404 564076 455004 564078
rect 490404 564076 491004 564078
rect 526404 564076 527004 564078
rect 562404 564076 563004 564078
rect 588140 564076 588740 564078
rect -4816 564054 588740 564076
rect -4816 563818 -4634 564054
rect -4398 563818 22586 564054
rect 22822 563818 58586 564054
rect 58822 563818 94586 564054
rect 94822 563818 130586 564054
rect 130822 563818 166586 564054
rect 166822 563818 202586 564054
rect 202822 563818 238586 564054
rect 238822 563818 274586 564054
rect 274822 563818 310586 564054
rect 310822 563818 346586 564054
rect 346822 563818 382586 564054
rect 382822 563818 418586 564054
rect 418822 563818 454586 564054
rect 454822 563818 490586 564054
rect 490822 563818 526586 564054
rect 526822 563818 562586 564054
rect 562822 563818 588322 564054
rect 588558 563818 588740 564054
rect -4816 563734 588740 563818
rect -4816 563498 -4634 563734
rect -4398 563498 22586 563734
rect 22822 563498 58586 563734
rect 58822 563498 94586 563734
rect 94822 563498 130586 563734
rect 130822 563498 166586 563734
rect 166822 563498 202586 563734
rect 202822 563498 238586 563734
rect 238822 563498 274586 563734
rect 274822 563498 310586 563734
rect 310822 563498 346586 563734
rect 346822 563498 382586 563734
rect 382822 563498 418586 563734
rect 418822 563498 454586 563734
rect 454822 563498 490586 563734
rect 490822 563498 526586 563734
rect 526822 563498 562586 563734
rect 562822 563498 588322 563734
rect 588558 563498 588740 563734
rect -4816 563476 588740 563498
rect -4816 563474 -4216 563476
rect 22404 563474 23004 563476
rect 58404 563474 59004 563476
rect 94404 563474 95004 563476
rect 130404 563474 131004 563476
rect 166404 563474 167004 563476
rect 202404 563474 203004 563476
rect 238404 563474 239004 563476
rect 274404 563474 275004 563476
rect 310404 563474 311004 563476
rect 346404 563474 347004 563476
rect 382404 563474 383004 563476
rect 418404 563474 419004 563476
rect 454404 563474 455004 563476
rect 490404 563474 491004 563476
rect 526404 563474 527004 563476
rect 562404 563474 563004 563476
rect 588140 563474 588740 563476
rect -2936 560476 -2336 560478
rect 18804 560476 19404 560478
rect 54804 560476 55404 560478
rect 90804 560476 91404 560478
rect 126804 560476 127404 560478
rect 162804 560476 163404 560478
rect 198804 560476 199404 560478
rect 234804 560476 235404 560478
rect 270804 560476 271404 560478
rect 306804 560476 307404 560478
rect 342804 560476 343404 560478
rect 378804 560476 379404 560478
rect 414804 560476 415404 560478
rect 450804 560476 451404 560478
rect 486804 560476 487404 560478
rect 522804 560476 523404 560478
rect 558804 560476 559404 560478
rect 586260 560476 586860 560478
rect -2936 560454 586860 560476
rect -2936 560218 -2754 560454
rect -2518 560218 18986 560454
rect 19222 560218 54986 560454
rect 55222 560218 90986 560454
rect 91222 560218 126986 560454
rect 127222 560218 162986 560454
rect 163222 560218 198986 560454
rect 199222 560218 234986 560454
rect 235222 560218 270986 560454
rect 271222 560218 306986 560454
rect 307222 560218 342986 560454
rect 343222 560218 378986 560454
rect 379222 560218 414986 560454
rect 415222 560218 450986 560454
rect 451222 560218 486986 560454
rect 487222 560218 522986 560454
rect 523222 560218 558986 560454
rect 559222 560218 586442 560454
rect 586678 560218 586860 560454
rect -2936 560134 586860 560218
rect -2936 559898 -2754 560134
rect -2518 559898 18986 560134
rect 19222 559898 54986 560134
rect 55222 559898 90986 560134
rect 91222 559898 126986 560134
rect 127222 559898 162986 560134
rect 163222 559898 198986 560134
rect 199222 559898 234986 560134
rect 235222 559898 270986 560134
rect 271222 559898 306986 560134
rect 307222 559898 342986 560134
rect 343222 559898 378986 560134
rect 379222 559898 414986 560134
rect 415222 559898 450986 560134
rect 451222 559898 486986 560134
rect 487222 559898 522986 560134
rect 523222 559898 558986 560134
rect 559222 559898 586442 560134
rect 586678 559898 586860 560134
rect -2936 559876 586860 559898
rect -2936 559874 -2336 559876
rect 18804 559874 19404 559876
rect 54804 559874 55404 559876
rect 90804 559874 91404 559876
rect 126804 559874 127404 559876
rect 162804 559874 163404 559876
rect 198804 559874 199404 559876
rect 234804 559874 235404 559876
rect 270804 559874 271404 559876
rect 306804 559874 307404 559876
rect 342804 559874 343404 559876
rect 378804 559874 379404 559876
rect 414804 559874 415404 559876
rect 450804 559874 451404 559876
rect 486804 559874 487404 559876
rect 522804 559874 523404 559876
rect 558804 559874 559404 559876
rect 586260 559874 586860 559876
rect -7636 553276 -7036 553278
rect 11604 553276 12204 553278
rect 47604 553276 48204 553278
rect 83604 553276 84204 553278
rect 119604 553276 120204 553278
rect 155604 553276 156204 553278
rect 191604 553276 192204 553278
rect 227604 553276 228204 553278
rect 263604 553276 264204 553278
rect 299604 553276 300204 553278
rect 335604 553276 336204 553278
rect 371604 553276 372204 553278
rect 407604 553276 408204 553278
rect 443604 553276 444204 553278
rect 479604 553276 480204 553278
rect 515604 553276 516204 553278
rect 551604 553276 552204 553278
rect 590960 553276 591560 553278
rect -8576 553254 592500 553276
rect -8576 553018 -7454 553254
rect -7218 553018 11786 553254
rect 12022 553018 47786 553254
rect 48022 553018 83786 553254
rect 84022 553018 119786 553254
rect 120022 553018 155786 553254
rect 156022 553018 191786 553254
rect 192022 553018 227786 553254
rect 228022 553018 263786 553254
rect 264022 553018 299786 553254
rect 300022 553018 335786 553254
rect 336022 553018 371786 553254
rect 372022 553018 407786 553254
rect 408022 553018 443786 553254
rect 444022 553018 479786 553254
rect 480022 553018 515786 553254
rect 516022 553018 551786 553254
rect 552022 553018 591142 553254
rect 591378 553018 592500 553254
rect -8576 552934 592500 553018
rect -8576 552698 -7454 552934
rect -7218 552698 11786 552934
rect 12022 552698 47786 552934
rect 48022 552698 83786 552934
rect 84022 552698 119786 552934
rect 120022 552698 155786 552934
rect 156022 552698 191786 552934
rect 192022 552698 227786 552934
rect 228022 552698 263786 552934
rect 264022 552698 299786 552934
rect 300022 552698 335786 552934
rect 336022 552698 371786 552934
rect 372022 552698 407786 552934
rect 408022 552698 443786 552934
rect 444022 552698 479786 552934
rect 480022 552698 515786 552934
rect 516022 552698 551786 552934
rect 552022 552698 591142 552934
rect 591378 552698 592500 552934
rect -8576 552676 592500 552698
rect -7636 552674 -7036 552676
rect 11604 552674 12204 552676
rect 47604 552674 48204 552676
rect 83604 552674 84204 552676
rect 119604 552674 120204 552676
rect 155604 552674 156204 552676
rect 191604 552674 192204 552676
rect 227604 552674 228204 552676
rect 263604 552674 264204 552676
rect 299604 552674 300204 552676
rect 335604 552674 336204 552676
rect 371604 552674 372204 552676
rect 407604 552674 408204 552676
rect 443604 552674 444204 552676
rect 479604 552674 480204 552676
rect 515604 552674 516204 552676
rect 551604 552674 552204 552676
rect 590960 552674 591560 552676
rect -5756 549676 -5156 549678
rect 8004 549676 8604 549678
rect 44004 549676 44604 549678
rect 80004 549676 80604 549678
rect 116004 549676 116604 549678
rect 152004 549676 152604 549678
rect 188004 549676 188604 549678
rect 224004 549676 224604 549678
rect 260004 549676 260604 549678
rect 296004 549676 296604 549678
rect 332004 549676 332604 549678
rect 368004 549676 368604 549678
rect 404004 549676 404604 549678
rect 440004 549676 440604 549678
rect 476004 549676 476604 549678
rect 512004 549676 512604 549678
rect 548004 549676 548604 549678
rect 589080 549676 589680 549678
rect -6696 549654 590620 549676
rect -6696 549418 -5574 549654
rect -5338 549418 8186 549654
rect 8422 549418 44186 549654
rect 44422 549418 80186 549654
rect 80422 549418 116186 549654
rect 116422 549418 152186 549654
rect 152422 549418 188186 549654
rect 188422 549418 224186 549654
rect 224422 549418 260186 549654
rect 260422 549418 296186 549654
rect 296422 549418 332186 549654
rect 332422 549418 368186 549654
rect 368422 549418 404186 549654
rect 404422 549418 440186 549654
rect 440422 549418 476186 549654
rect 476422 549418 512186 549654
rect 512422 549418 548186 549654
rect 548422 549418 589262 549654
rect 589498 549418 590620 549654
rect -6696 549334 590620 549418
rect -6696 549098 -5574 549334
rect -5338 549098 8186 549334
rect 8422 549098 44186 549334
rect 44422 549098 80186 549334
rect 80422 549098 116186 549334
rect 116422 549098 152186 549334
rect 152422 549098 188186 549334
rect 188422 549098 224186 549334
rect 224422 549098 260186 549334
rect 260422 549098 296186 549334
rect 296422 549098 332186 549334
rect 332422 549098 368186 549334
rect 368422 549098 404186 549334
rect 404422 549098 440186 549334
rect 440422 549098 476186 549334
rect 476422 549098 512186 549334
rect 512422 549098 548186 549334
rect 548422 549098 589262 549334
rect 589498 549098 590620 549334
rect -6696 549076 590620 549098
rect -5756 549074 -5156 549076
rect 8004 549074 8604 549076
rect 44004 549074 44604 549076
rect 80004 549074 80604 549076
rect 116004 549074 116604 549076
rect 152004 549074 152604 549076
rect 188004 549074 188604 549076
rect 224004 549074 224604 549076
rect 260004 549074 260604 549076
rect 296004 549074 296604 549076
rect 332004 549074 332604 549076
rect 368004 549074 368604 549076
rect 404004 549074 404604 549076
rect 440004 549074 440604 549076
rect 476004 549074 476604 549076
rect 512004 549074 512604 549076
rect 548004 549074 548604 549076
rect 589080 549074 589680 549076
rect -3876 546076 -3276 546078
rect 4404 546076 5004 546078
rect 40404 546076 41004 546078
rect 76404 546076 77004 546078
rect 112404 546076 113004 546078
rect 148404 546076 149004 546078
rect 184404 546076 185004 546078
rect 220404 546076 221004 546078
rect 256404 546076 257004 546078
rect 292404 546076 293004 546078
rect 328404 546076 329004 546078
rect 364404 546076 365004 546078
rect 400404 546076 401004 546078
rect 436404 546076 437004 546078
rect 472404 546076 473004 546078
rect 508404 546076 509004 546078
rect 544404 546076 545004 546078
rect 580404 546076 581004 546078
rect 587200 546076 587800 546078
rect -4816 546054 588740 546076
rect -4816 545818 -3694 546054
rect -3458 545818 4586 546054
rect 4822 545818 40586 546054
rect 40822 545818 76586 546054
rect 76822 545818 112586 546054
rect 112822 545818 148586 546054
rect 148822 545818 184586 546054
rect 184822 545818 220586 546054
rect 220822 545818 256586 546054
rect 256822 545818 292586 546054
rect 292822 545818 328586 546054
rect 328822 545818 364586 546054
rect 364822 545818 400586 546054
rect 400822 545818 436586 546054
rect 436822 545818 472586 546054
rect 472822 545818 508586 546054
rect 508822 545818 544586 546054
rect 544822 545818 580586 546054
rect 580822 545818 587382 546054
rect 587618 545818 588740 546054
rect -4816 545734 588740 545818
rect -4816 545498 -3694 545734
rect -3458 545498 4586 545734
rect 4822 545498 40586 545734
rect 40822 545498 76586 545734
rect 76822 545498 112586 545734
rect 112822 545498 148586 545734
rect 148822 545498 184586 545734
rect 184822 545498 220586 545734
rect 220822 545498 256586 545734
rect 256822 545498 292586 545734
rect 292822 545498 328586 545734
rect 328822 545498 364586 545734
rect 364822 545498 400586 545734
rect 400822 545498 436586 545734
rect 436822 545498 472586 545734
rect 472822 545498 508586 545734
rect 508822 545498 544586 545734
rect 544822 545498 580586 545734
rect 580822 545498 587382 545734
rect 587618 545498 588740 545734
rect -4816 545476 588740 545498
rect -3876 545474 -3276 545476
rect 4404 545474 5004 545476
rect 40404 545474 41004 545476
rect 76404 545474 77004 545476
rect 112404 545474 113004 545476
rect 148404 545474 149004 545476
rect 184404 545474 185004 545476
rect 220404 545474 221004 545476
rect 256404 545474 257004 545476
rect 292404 545474 293004 545476
rect 328404 545474 329004 545476
rect 364404 545474 365004 545476
rect 400404 545474 401004 545476
rect 436404 545474 437004 545476
rect 472404 545474 473004 545476
rect 508404 545474 509004 545476
rect 544404 545474 545004 545476
rect 580404 545474 581004 545476
rect 587200 545474 587800 545476
rect -1996 542476 -1396 542478
rect 804 542476 1404 542478
rect 36804 542476 37404 542478
rect 72804 542476 73404 542478
rect 108804 542476 109404 542478
rect 144804 542476 145404 542478
rect 180804 542476 181404 542478
rect 216804 542476 217404 542478
rect 252804 542476 253404 542478
rect 288804 542476 289404 542478
rect 324804 542476 325404 542478
rect 360804 542476 361404 542478
rect 396804 542476 397404 542478
rect 432804 542476 433404 542478
rect 468804 542476 469404 542478
rect 504804 542476 505404 542478
rect 540804 542476 541404 542478
rect 576804 542476 577404 542478
rect 585320 542476 585920 542478
rect -2936 542454 586860 542476
rect -2936 542218 -1814 542454
rect -1578 542218 986 542454
rect 1222 542218 36986 542454
rect 37222 542218 72986 542454
rect 73222 542218 108986 542454
rect 109222 542218 144986 542454
rect 145222 542218 180986 542454
rect 181222 542218 216986 542454
rect 217222 542218 252986 542454
rect 253222 542218 288986 542454
rect 289222 542218 324986 542454
rect 325222 542218 360986 542454
rect 361222 542218 396986 542454
rect 397222 542218 432986 542454
rect 433222 542218 468986 542454
rect 469222 542218 504986 542454
rect 505222 542218 540986 542454
rect 541222 542218 576986 542454
rect 577222 542218 585502 542454
rect 585738 542218 586860 542454
rect -2936 542134 586860 542218
rect -2936 541898 -1814 542134
rect -1578 541898 986 542134
rect 1222 541898 36986 542134
rect 37222 541898 72986 542134
rect 73222 541898 108986 542134
rect 109222 541898 144986 542134
rect 145222 541898 180986 542134
rect 181222 541898 216986 542134
rect 217222 541898 252986 542134
rect 253222 541898 288986 542134
rect 289222 541898 324986 542134
rect 325222 541898 360986 542134
rect 361222 541898 396986 542134
rect 397222 541898 432986 542134
rect 433222 541898 468986 542134
rect 469222 541898 504986 542134
rect 505222 541898 540986 542134
rect 541222 541898 576986 542134
rect 577222 541898 585502 542134
rect 585738 541898 586860 542134
rect -2936 541876 586860 541898
rect -1996 541874 -1396 541876
rect 804 541874 1404 541876
rect 36804 541874 37404 541876
rect 72804 541874 73404 541876
rect 108804 541874 109404 541876
rect 144804 541874 145404 541876
rect 180804 541874 181404 541876
rect 216804 541874 217404 541876
rect 252804 541874 253404 541876
rect 288804 541874 289404 541876
rect 324804 541874 325404 541876
rect 360804 541874 361404 541876
rect 396804 541874 397404 541876
rect 432804 541874 433404 541876
rect 468804 541874 469404 541876
rect 504804 541874 505404 541876
rect 540804 541874 541404 541876
rect 576804 541874 577404 541876
rect 585320 541874 585920 541876
rect -8576 535276 -7976 535278
rect 29604 535276 30204 535278
rect 65604 535276 66204 535278
rect 101604 535276 102204 535278
rect 137604 535276 138204 535278
rect 173604 535276 174204 535278
rect 209604 535276 210204 535278
rect 245604 535276 246204 535278
rect 281604 535276 282204 535278
rect 317604 535276 318204 535278
rect 353604 535276 354204 535278
rect 389604 535276 390204 535278
rect 425604 535276 426204 535278
rect 461604 535276 462204 535278
rect 497604 535276 498204 535278
rect 533604 535276 534204 535278
rect 569604 535276 570204 535278
rect 591900 535276 592500 535278
rect -8576 535254 592500 535276
rect -8576 535018 -8394 535254
rect -8158 535018 29786 535254
rect 30022 535018 65786 535254
rect 66022 535018 101786 535254
rect 102022 535018 137786 535254
rect 138022 535018 173786 535254
rect 174022 535018 209786 535254
rect 210022 535018 245786 535254
rect 246022 535018 281786 535254
rect 282022 535018 317786 535254
rect 318022 535018 353786 535254
rect 354022 535018 389786 535254
rect 390022 535018 425786 535254
rect 426022 535018 461786 535254
rect 462022 535018 497786 535254
rect 498022 535018 533786 535254
rect 534022 535018 569786 535254
rect 570022 535018 592082 535254
rect 592318 535018 592500 535254
rect -8576 534934 592500 535018
rect -8576 534698 -8394 534934
rect -8158 534698 29786 534934
rect 30022 534698 65786 534934
rect 66022 534698 101786 534934
rect 102022 534698 137786 534934
rect 138022 534698 173786 534934
rect 174022 534698 209786 534934
rect 210022 534698 245786 534934
rect 246022 534698 281786 534934
rect 282022 534698 317786 534934
rect 318022 534698 353786 534934
rect 354022 534698 389786 534934
rect 390022 534698 425786 534934
rect 426022 534698 461786 534934
rect 462022 534698 497786 534934
rect 498022 534698 533786 534934
rect 534022 534698 569786 534934
rect 570022 534698 592082 534934
rect 592318 534698 592500 534934
rect -8576 534676 592500 534698
rect -8576 534674 -7976 534676
rect 29604 534674 30204 534676
rect 65604 534674 66204 534676
rect 101604 534674 102204 534676
rect 137604 534674 138204 534676
rect 173604 534674 174204 534676
rect 209604 534674 210204 534676
rect 245604 534674 246204 534676
rect 281604 534674 282204 534676
rect 317604 534674 318204 534676
rect 353604 534674 354204 534676
rect 389604 534674 390204 534676
rect 425604 534674 426204 534676
rect 461604 534674 462204 534676
rect 497604 534674 498204 534676
rect 533604 534674 534204 534676
rect 569604 534674 570204 534676
rect 591900 534674 592500 534676
rect -6696 531676 -6096 531678
rect 26004 531676 26604 531678
rect 62004 531676 62604 531678
rect 98004 531676 98604 531678
rect 134004 531676 134604 531678
rect 170004 531676 170604 531678
rect 206004 531676 206604 531678
rect 242004 531676 242604 531678
rect 278004 531676 278604 531678
rect 314004 531676 314604 531678
rect 350004 531676 350604 531678
rect 386004 531676 386604 531678
rect 422004 531676 422604 531678
rect 458004 531676 458604 531678
rect 494004 531676 494604 531678
rect 530004 531676 530604 531678
rect 566004 531676 566604 531678
rect 590020 531676 590620 531678
rect -6696 531654 590620 531676
rect -6696 531418 -6514 531654
rect -6278 531418 26186 531654
rect 26422 531418 62186 531654
rect 62422 531418 98186 531654
rect 98422 531418 134186 531654
rect 134422 531418 170186 531654
rect 170422 531418 206186 531654
rect 206422 531418 242186 531654
rect 242422 531418 278186 531654
rect 278422 531418 314186 531654
rect 314422 531418 350186 531654
rect 350422 531418 386186 531654
rect 386422 531418 422186 531654
rect 422422 531418 458186 531654
rect 458422 531418 494186 531654
rect 494422 531418 530186 531654
rect 530422 531418 566186 531654
rect 566422 531418 590202 531654
rect 590438 531418 590620 531654
rect -6696 531334 590620 531418
rect -6696 531098 -6514 531334
rect -6278 531098 26186 531334
rect 26422 531098 62186 531334
rect 62422 531098 98186 531334
rect 98422 531098 134186 531334
rect 134422 531098 170186 531334
rect 170422 531098 206186 531334
rect 206422 531098 242186 531334
rect 242422 531098 278186 531334
rect 278422 531098 314186 531334
rect 314422 531098 350186 531334
rect 350422 531098 386186 531334
rect 386422 531098 422186 531334
rect 422422 531098 458186 531334
rect 458422 531098 494186 531334
rect 494422 531098 530186 531334
rect 530422 531098 566186 531334
rect 566422 531098 590202 531334
rect 590438 531098 590620 531334
rect -6696 531076 590620 531098
rect -6696 531074 -6096 531076
rect 26004 531074 26604 531076
rect 62004 531074 62604 531076
rect 98004 531074 98604 531076
rect 134004 531074 134604 531076
rect 170004 531074 170604 531076
rect 206004 531074 206604 531076
rect 242004 531074 242604 531076
rect 278004 531074 278604 531076
rect 314004 531074 314604 531076
rect 350004 531074 350604 531076
rect 386004 531074 386604 531076
rect 422004 531074 422604 531076
rect 458004 531074 458604 531076
rect 494004 531074 494604 531076
rect 530004 531074 530604 531076
rect 566004 531074 566604 531076
rect 590020 531074 590620 531076
rect -4816 528076 -4216 528078
rect 22404 528076 23004 528078
rect 58404 528076 59004 528078
rect 94404 528076 95004 528078
rect 130404 528076 131004 528078
rect 166404 528076 167004 528078
rect 202404 528076 203004 528078
rect 238404 528076 239004 528078
rect 274404 528076 275004 528078
rect 310404 528076 311004 528078
rect 346404 528076 347004 528078
rect 382404 528076 383004 528078
rect 418404 528076 419004 528078
rect 454404 528076 455004 528078
rect 490404 528076 491004 528078
rect 526404 528076 527004 528078
rect 562404 528076 563004 528078
rect 588140 528076 588740 528078
rect -4816 528054 588740 528076
rect -4816 527818 -4634 528054
rect -4398 527818 22586 528054
rect 22822 527818 58586 528054
rect 58822 527818 94586 528054
rect 94822 527818 130586 528054
rect 130822 527818 166586 528054
rect 166822 527818 202586 528054
rect 202822 527818 238586 528054
rect 238822 527818 274586 528054
rect 274822 527818 310586 528054
rect 310822 527818 346586 528054
rect 346822 527818 382586 528054
rect 382822 527818 418586 528054
rect 418822 527818 454586 528054
rect 454822 527818 490586 528054
rect 490822 527818 526586 528054
rect 526822 527818 562586 528054
rect 562822 527818 588322 528054
rect 588558 527818 588740 528054
rect -4816 527734 588740 527818
rect -4816 527498 -4634 527734
rect -4398 527498 22586 527734
rect 22822 527498 58586 527734
rect 58822 527498 94586 527734
rect 94822 527498 130586 527734
rect 130822 527498 166586 527734
rect 166822 527498 202586 527734
rect 202822 527498 238586 527734
rect 238822 527498 274586 527734
rect 274822 527498 310586 527734
rect 310822 527498 346586 527734
rect 346822 527498 382586 527734
rect 382822 527498 418586 527734
rect 418822 527498 454586 527734
rect 454822 527498 490586 527734
rect 490822 527498 526586 527734
rect 526822 527498 562586 527734
rect 562822 527498 588322 527734
rect 588558 527498 588740 527734
rect -4816 527476 588740 527498
rect -4816 527474 -4216 527476
rect 22404 527474 23004 527476
rect 58404 527474 59004 527476
rect 94404 527474 95004 527476
rect 130404 527474 131004 527476
rect 166404 527474 167004 527476
rect 202404 527474 203004 527476
rect 238404 527474 239004 527476
rect 274404 527474 275004 527476
rect 310404 527474 311004 527476
rect 346404 527474 347004 527476
rect 382404 527474 383004 527476
rect 418404 527474 419004 527476
rect 454404 527474 455004 527476
rect 490404 527474 491004 527476
rect 526404 527474 527004 527476
rect 562404 527474 563004 527476
rect 588140 527474 588740 527476
rect -2936 524476 -2336 524478
rect 18804 524476 19404 524478
rect 54804 524476 55404 524478
rect 90804 524476 91404 524478
rect 126804 524476 127404 524478
rect 162804 524476 163404 524478
rect 198804 524476 199404 524478
rect 234804 524476 235404 524478
rect 270804 524476 271404 524478
rect 306804 524476 307404 524478
rect 342804 524476 343404 524478
rect 378804 524476 379404 524478
rect 414804 524476 415404 524478
rect 450804 524476 451404 524478
rect 486804 524476 487404 524478
rect 522804 524476 523404 524478
rect 558804 524476 559404 524478
rect 586260 524476 586860 524478
rect -2936 524454 586860 524476
rect -2936 524218 -2754 524454
rect -2518 524218 18986 524454
rect 19222 524218 54986 524454
rect 55222 524218 90986 524454
rect 91222 524218 126986 524454
rect 127222 524218 162986 524454
rect 163222 524218 198986 524454
rect 199222 524218 234986 524454
rect 235222 524218 270986 524454
rect 271222 524218 306986 524454
rect 307222 524218 342986 524454
rect 343222 524218 378986 524454
rect 379222 524218 414986 524454
rect 415222 524218 450986 524454
rect 451222 524218 486986 524454
rect 487222 524218 522986 524454
rect 523222 524218 558986 524454
rect 559222 524218 586442 524454
rect 586678 524218 586860 524454
rect -2936 524134 586860 524218
rect -2936 523898 -2754 524134
rect -2518 523898 18986 524134
rect 19222 523898 54986 524134
rect 55222 523898 90986 524134
rect 91222 523898 126986 524134
rect 127222 523898 162986 524134
rect 163222 523898 198986 524134
rect 199222 523898 234986 524134
rect 235222 523898 270986 524134
rect 271222 523898 306986 524134
rect 307222 523898 342986 524134
rect 343222 523898 378986 524134
rect 379222 523898 414986 524134
rect 415222 523898 450986 524134
rect 451222 523898 486986 524134
rect 487222 523898 522986 524134
rect 523222 523898 558986 524134
rect 559222 523898 586442 524134
rect 586678 523898 586860 524134
rect -2936 523876 586860 523898
rect -2936 523874 -2336 523876
rect 18804 523874 19404 523876
rect 54804 523874 55404 523876
rect 90804 523874 91404 523876
rect 126804 523874 127404 523876
rect 162804 523874 163404 523876
rect 198804 523874 199404 523876
rect 234804 523874 235404 523876
rect 270804 523874 271404 523876
rect 306804 523874 307404 523876
rect 342804 523874 343404 523876
rect 378804 523874 379404 523876
rect 414804 523874 415404 523876
rect 450804 523874 451404 523876
rect 486804 523874 487404 523876
rect 522804 523874 523404 523876
rect 558804 523874 559404 523876
rect 586260 523874 586860 523876
rect -7636 517276 -7036 517278
rect 11604 517276 12204 517278
rect 47604 517276 48204 517278
rect 83604 517276 84204 517278
rect 119604 517276 120204 517278
rect 155604 517276 156204 517278
rect 191604 517276 192204 517278
rect 227604 517276 228204 517278
rect 263604 517276 264204 517278
rect 299604 517276 300204 517278
rect 335604 517276 336204 517278
rect 371604 517276 372204 517278
rect 407604 517276 408204 517278
rect 443604 517276 444204 517278
rect 479604 517276 480204 517278
rect 515604 517276 516204 517278
rect 551604 517276 552204 517278
rect 590960 517276 591560 517278
rect -8576 517254 592500 517276
rect -8576 517018 -7454 517254
rect -7218 517018 11786 517254
rect 12022 517018 47786 517254
rect 48022 517018 83786 517254
rect 84022 517018 119786 517254
rect 120022 517018 155786 517254
rect 156022 517018 191786 517254
rect 192022 517018 227786 517254
rect 228022 517018 263786 517254
rect 264022 517018 299786 517254
rect 300022 517018 335786 517254
rect 336022 517018 371786 517254
rect 372022 517018 407786 517254
rect 408022 517018 443786 517254
rect 444022 517018 479786 517254
rect 480022 517018 515786 517254
rect 516022 517018 551786 517254
rect 552022 517018 591142 517254
rect 591378 517018 592500 517254
rect -8576 516934 592500 517018
rect -8576 516698 -7454 516934
rect -7218 516698 11786 516934
rect 12022 516698 47786 516934
rect 48022 516698 83786 516934
rect 84022 516698 119786 516934
rect 120022 516698 155786 516934
rect 156022 516698 191786 516934
rect 192022 516698 227786 516934
rect 228022 516698 263786 516934
rect 264022 516698 299786 516934
rect 300022 516698 335786 516934
rect 336022 516698 371786 516934
rect 372022 516698 407786 516934
rect 408022 516698 443786 516934
rect 444022 516698 479786 516934
rect 480022 516698 515786 516934
rect 516022 516698 551786 516934
rect 552022 516698 591142 516934
rect 591378 516698 592500 516934
rect -8576 516676 592500 516698
rect -7636 516674 -7036 516676
rect 11604 516674 12204 516676
rect 47604 516674 48204 516676
rect 83604 516674 84204 516676
rect 119604 516674 120204 516676
rect 155604 516674 156204 516676
rect 191604 516674 192204 516676
rect 227604 516674 228204 516676
rect 263604 516674 264204 516676
rect 299604 516674 300204 516676
rect 335604 516674 336204 516676
rect 371604 516674 372204 516676
rect 407604 516674 408204 516676
rect 443604 516674 444204 516676
rect 479604 516674 480204 516676
rect 515604 516674 516204 516676
rect 551604 516674 552204 516676
rect 590960 516674 591560 516676
rect -5756 513676 -5156 513678
rect 8004 513676 8604 513678
rect 44004 513676 44604 513678
rect 80004 513676 80604 513678
rect 116004 513676 116604 513678
rect 152004 513676 152604 513678
rect 188004 513676 188604 513678
rect 224004 513676 224604 513678
rect 260004 513676 260604 513678
rect 296004 513676 296604 513678
rect 332004 513676 332604 513678
rect 368004 513676 368604 513678
rect 404004 513676 404604 513678
rect 440004 513676 440604 513678
rect 476004 513676 476604 513678
rect 512004 513676 512604 513678
rect 548004 513676 548604 513678
rect 589080 513676 589680 513678
rect -6696 513654 590620 513676
rect -6696 513418 -5574 513654
rect -5338 513418 8186 513654
rect 8422 513418 44186 513654
rect 44422 513418 80186 513654
rect 80422 513418 116186 513654
rect 116422 513418 152186 513654
rect 152422 513418 188186 513654
rect 188422 513418 224186 513654
rect 224422 513418 260186 513654
rect 260422 513418 296186 513654
rect 296422 513418 332186 513654
rect 332422 513418 368186 513654
rect 368422 513418 404186 513654
rect 404422 513418 440186 513654
rect 440422 513418 476186 513654
rect 476422 513418 512186 513654
rect 512422 513418 548186 513654
rect 548422 513418 589262 513654
rect 589498 513418 590620 513654
rect -6696 513334 590620 513418
rect -6696 513098 -5574 513334
rect -5338 513098 8186 513334
rect 8422 513098 44186 513334
rect 44422 513098 80186 513334
rect 80422 513098 116186 513334
rect 116422 513098 152186 513334
rect 152422 513098 188186 513334
rect 188422 513098 224186 513334
rect 224422 513098 260186 513334
rect 260422 513098 296186 513334
rect 296422 513098 332186 513334
rect 332422 513098 368186 513334
rect 368422 513098 404186 513334
rect 404422 513098 440186 513334
rect 440422 513098 476186 513334
rect 476422 513098 512186 513334
rect 512422 513098 548186 513334
rect 548422 513098 589262 513334
rect 589498 513098 590620 513334
rect -6696 513076 590620 513098
rect -5756 513074 -5156 513076
rect 8004 513074 8604 513076
rect 44004 513074 44604 513076
rect 80004 513074 80604 513076
rect 116004 513074 116604 513076
rect 152004 513074 152604 513076
rect 188004 513074 188604 513076
rect 224004 513074 224604 513076
rect 260004 513074 260604 513076
rect 296004 513074 296604 513076
rect 332004 513074 332604 513076
rect 368004 513074 368604 513076
rect 404004 513074 404604 513076
rect 440004 513074 440604 513076
rect 476004 513074 476604 513076
rect 512004 513074 512604 513076
rect 548004 513074 548604 513076
rect 589080 513074 589680 513076
rect -3876 510076 -3276 510078
rect 4404 510076 5004 510078
rect 40404 510076 41004 510078
rect 76404 510076 77004 510078
rect 112404 510076 113004 510078
rect 148404 510076 149004 510078
rect 184404 510076 185004 510078
rect 220404 510076 221004 510078
rect 256404 510076 257004 510078
rect 292404 510076 293004 510078
rect 328404 510076 329004 510078
rect 364404 510076 365004 510078
rect 400404 510076 401004 510078
rect 436404 510076 437004 510078
rect 472404 510076 473004 510078
rect 508404 510076 509004 510078
rect 544404 510076 545004 510078
rect 580404 510076 581004 510078
rect 587200 510076 587800 510078
rect -4816 510054 588740 510076
rect -4816 509818 -3694 510054
rect -3458 509818 4586 510054
rect 4822 509818 40586 510054
rect 40822 509818 76586 510054
rect 76822 509818 112586 510054
rect 112822 509818 148586 510054
rect 148822 509818 184586 510054
rect 184822 509818 220586 510054
rect 220822 509818 256586 510054
rect 256822 509818 292586 510054
rect 292822 509818 328586 510054
rect 328822 509818 364586 510054
rect 364822 509818 400586 510054
rect 400822 509818 436586 510054
rect 436822 509818 472586 510054
rect 472822 509818 508586 510054
rect 508822 509818 544586 510054
rect 544822 509818 580586 510054
rect 580822 509818 587382 510054
rect 587618 509818 588740 510054
rect -4816 509734 588740 509818
rect -4816 509498 -3694 509734
rect -3458 509498 4586 509734
rect 4822 509498 40586 509734
rect 40822 509498 76586 509734
rect 76822 509498 112586 509734
rect 112822 509498 148586 509734
rect 148822 509498 184586 509734
rect 184822 509498 220586 509734
rect 220822 509498 256586 509734
rect 256822 509498 292586 509734
rect 292822 509498 328586 509734
rect 328822 509498 364586 509734
rect 364822 509498 400586 509734
rect 400822 509498 436586 509734
rect 436822 509498 472586 509734
rect 472822 509498 508586 509734
rect 508822 509498 544586 509734
rect 544822 509498 580586 509734
rect 580822 509498 587382 509734
rect 587618 509498 588740 509734
rect -4816 509476 588740 509498
rect -3876 509474 -3276 509476
rect 4404 509474 5004 509476
rect 40404 509474 41004 509476
rect 76404 509474 77004 509476
rect 112404 509474 113004 509476
rect 148404 509474 149004 509476
rect 184404 509474 185004 509476
rect 220404 509474 221004 509476
rect 256404 509474 257004 509476
rect 292404 509474 293004 509476
rect 328404 509474 329004 509476
rect 364404 509474 365004 509476
rect 400404 509474 401004 509476
rect 436404 509474 437004 509476
rect 472404 509474 473004 509476
rect 508404 509474 509004 509476
rect 544404 509474 545004 509476
rect 580404 509474 581004 509476
rect 587200 509474 587800 509476
rect -1996 506476 -1396 506478
rect 804 506476 1404 506478
rect 36804 506476 37404 506478
rect 72804 506476 73404 506478
rect 108804 506476 109404 506478
rect 144804 506476 145404 506478
rect 180804 506476 181404 506478
rect 216804 506476 217404 506478
rect 252804 506476 253404 506478
rect 288804 506476 289404 506478
rect 324804 506476 325404 506478
rect 360804 506476 361404 506478
rect 396804 506476 397404 506478
rect 432804 506476 433404 506478
rect 468804 506476 469404 506478
rect 504804 506476 505404 506478
rect 540804 506476 541404 506478
rect 576804 506476 577404 506478
rect 585320 506476 585920 506478
rect -2936 506454 586860 506476
rect -2936 506218 -1814 506454
rect -1578 506218 986 506454
rect 1222 506218 36986 506454
rect 37222 506218 72986 506454
rect 73222 506218 108986 506454
rect 109222 506218 144986 506454
rect 145222 506218 180986 506454
rect 181222 506218 216986 506454
rect 217222 506218 252986 506454
rect 253222 506218 288986 506454
rect 289222 506218 324986 506454
rect 325222 506218 360986 506454
rect 361222 506218 396986 506454
rect 397222 506218 432986 506454
rect 433222 506218 468986 506454
rect 469222 506218 504986 506454
rect 505222 506218 540986 506454
rect 541222 506218 576986 506454
rect 577222 506218 585502 506454
rect 585738 506218 586860 506454
rect -2936 506134 586860 506218
rect -2936 505898 -1814 506134
rect -1578 505898 986 506134
rect 1222 505898 36986 506134
rect 37222 505898 72986 506134
rect 73222 505898 108986 506134
rect 109222 505898 144986 506134
rect 145222 505898 180986 506134
rect 181222 505898 216986 506134
rect 217222 505898 252986 506134
rect 253222 505898 288986 506134
rect 289222 505898 324986 506134
rect 325222 505898 360986 506134
rect 361222 505898 396986 506134
rect 397222 505898 432986 506134
rect 433222 505898 468986 506134
rect 469222 505898 504986 506134
rect 505222 505898 540986 506134
rect 541222 505898 576986 506134
rect 577222 505898 585502 506134
rect 585738 505898 586860 506134
rect -2936 505876 586860 505898
rect -1996 505874 -1396 505876
rect 804 505874 1404 505876
rect 36804 505874 37404 505876
rect 72804 505874 73404 505876
rect 108804 505874 109404 505876
rect 144804 505874 145404 505876
rect 180804 505874 181404 505876
rect 216804 505874 217404 505876
rect 252804 505874 253404 505876
rect 288804 505874 289404 505876
rect 324804 505874 325404 505876
rect 360804 505874 361404 505876
rect 396804 505874 397404 505876
rect 432804 505874 433404 505876
rect 468804 505874 469404 505876
rect 504804 505874 505404 505876
rect 540804 505874 541404 505876
rect 576804 505874 577404 505876
rect 585320 505874 585920 505876
rect -8576 499276 -7976 499278
rect 29604 499276 30204 499278
rect 65604 499276 66204 499278
rect 101604 499276 102204 499278
rect 137604 499276 138204 499278
rect 173604 499276 174204 499278
rect 209604 499276 210204 499278
rect 245604 499276 246204 499278
rect 281604 499276 282204 499278
rect 317604 499276 318204 499278
rect 353604 499276 354204 499278
rect 389604 499276 390204 499278
rect 425604 499276 426204 499278
rect 461604 499276 462204 499278
rect 497604 499276 498204 499278
rect 533604 499276 534204 499278
rect 569604 499276 570204 499278
rect 591900 499276 592500 499278
rect -8576 499254 592500 499276
rect -8576 499018 -8394 499254
rect -8158 499018 29786 499254
rect 30022 499018 65786 499254
rect 66022 499018 101786 499254
rect 102022 499018 137786 499254
rect 138022 499018 173786 499254
rect 174022 499018 209786 499254
rect 210022 499018 245786 499254
rect 246022 499018 281786 499254
rect 282022 499018 317786 499254
rect 318022 499018 353786 499254
rect 354022 499018 389786 499254
rect 390022 499018 425786 499254
rect 426022 499018 461786 499254
rect 462022 499018 497786 499254
rect 498022 499018 533786 499254
rect 534022 499018 569786 499254
rect 570022 499018 592082 499254
rect 592318 499018 592500 499254
rect -8576 498934 592500 499018
rect -8576 498698 -8394 498934
rect -8158 498698 29786 498934
rect 30022 498698 65786 498934
rect 66022 498698 101786 498934
rect 102022 498698 137786 498934
rect 138022 498698 173786 498934
rect 174022 498698 209786 498934
rect 210022 498698 245786 498934
rect 246022 498698 281786 498934
rect 282022 498698 317786 498934
rect 318022 498698 353786 498934
rect 354022 498698 389786 498934
rect 390022 498698 425786 498934
rect 426022 498698 461786 498934
rect 462022 498698 497786 498934
rect 498022 498698 533786 498934
rect 534022 498698 569786 498934
rect 570022 498698 592082 498934
rect 592318 498698 592500 498934
rect -8576 498676 592500 498698
rect -8576 498674 -7976 498676
rect 29604 498674 30204 498676
rect 65604 498674 66204 498676
rect 101604 498674 102204 498676
rect 137604 498674 138204 498676
rect 173604 498674 174204 498676
rect 209604 498674 210204 498676
rect 245604 498674 246204 498676
rect 281604 498674 282204 498676
rect 317604 498674 318204 498676
rect 353604 498674 354204 498676
rect 389604 498674 390204 498676
rect 425604 498674 426204 498676
rect 461604 498674 462204 498676
rect 497604 498674 498204 498676
rect 533604 498674 534204 498676
rect 569604 498674 570204 498676
rect 591900 498674 592500 498676
rect -6696 495676 -6096 495678
rect 26004 495676 26604 495678
rect 62004 495676 62604 495678
rect 98004 495676 98604 495678
rect 134004 495676 134604 495678
rect 170004 495676 170604 495678
rect 206004 495676 206604 495678
rect 242004 495676 242604 495678
rect 278004 495676 278604 495678
rect 314004 495676 314604 495678
rect 350004 495676 350604 495678
rect 386004 495676 386604 495678
rect 422004 495676 422604 495678
rect 458004 495676 458604 495678
rect 494004 495676 494604 495678
rect 530004 495676 530604 495678
rect 566004 495676 566604 495678
rect 590020 495676 590620 495678
rect -6696 495654 590620 495676
rect -6696 495418 -6514 495654
rect -6278 495418 26186 495654
rect 26422 495418 62186 495654
rect 62422 495418 98186 495654
rect 98422 495418 134186 495654
rect 134422 495418 170186 495654
rect 170422 495418 206186 495654
rect 206422 495418 242186 495654
rect 242422 495418 278186 495654
rect 278422 495418 314186 495654
rect 314422 495418 350186 495654
rect 350422 495418 386186 495654
rect 386422 495418 422186 495654
rect 422422 495418 458186 495654
rect 458422 495418 494186 495654
rect 494422 495418 530186 495654
rect 530422 495418 566186 495654
rect 566422 495418 590202 495654
rect 590438 495418 590620 495654
rect -6696 495334 590620 495418
rect -6696 495098 -6514 495334
rect -6278 495098 26186 495334
rect 26422 495098 62186 495334
rect 62422 495098 98186 495334
rect 98422 495098 134186 495334
rect 134422 495098 170186 495334
rect 170422 495098 206186 495334
rect 206422 495098 242186 495334
rect 242422 495098 278186 495334
rect 278422 495098 314186 495334
rect 314422 495098 350186 495334
rect 350422 495098 386186 495334
rect 386422 495098 422186 495334
rect 422422 495098 458186 495334
rect 458422 495098 494186 495334
rect 494422 495098 530186 495334
rect 530422 495098 566186 495334
rect 566422 495098 590202 495334
rect 590438 495098 590620 495334
rect -6696 495076 590620 495098
rect -6696 495074 -6096 495076
rect 26004 495074 26604 495076
rect 62004 495074 62604 495076
rect 98004 495074 98604 495076
rect 134004 495074 134604 495076
rect 170004 495074 170604 495076
rect 206004 495074 206604 495076
rect 242004 495074 242604 495076
rect 278004 495074 278604 495076
rect 314004 495074 314604 495076
rect 350004 495074 350604 495076
rect 386004 495074 386604 495076
rect 422004 495074 422604 495076
rect 458004 495074 458604 495076
rect 494004 495074 494604 495076
rect 530004 495074 530604 495076
rect 566004 495074 566604 495076
rect 590020 495074 590620 495076
rect -4816 492076 -4216 492078
rect 22404 492076 23004 492078
rect 58404 492076 59004 492078
rect 94404 492076 95004 492078
rect 130404 492076 131004 492078
rect 166404 492076 167004 492078
rect 202404 492076 203004 492078
rect 238404 492076 239004 492078
rect 274404 492076 275004 492078
rect 310404 492076 311004 492078
rect 346404 492076 347004 492078
rect 382404 492076 383004 492078
rect 418404 492076 419004 492078
rect 454404 492076 455004 492078
rect 490404 492076 491004 492078
rect 526404 492076 527004 492078
rect 562404 492076 563004 492078
rect 588140 492076 588740 492078
rect -4816 492054 588740 492076
rect -4816 491818 -4634 492054
rect -4398 491818 22586 492054
rect 22822 491818 58586 492054
rect 58822 491818 94586 492054
rect 94822 491818 130586 492054
rect 130822 491818 166586 492054
rect 166822 491818 202586 492054
rect 202822 491818 238586 492054
rect 238822 491818 274586 492054
rect 274822 491818 310586 492054
rect 310822 491818 346586 492054
rect 346822 491818 382586 492054
rect 382822 491818 418586 492054
rect 418822 491818 454586 492054
rect 454822 491818 490586 492054
rect 490822 491818 526586 492054
rect 526822 491818 562586 492054
rect 562822 491818 588322 492054
rect 588558 491818 588740 492054
rect -4816 491734 588740 491818
rect -4816 491498 -4634 491734
rect -4398 491498 22586 491734
rect 22822 491498 58586 491734
rect 58822 491498 94586 491734
rect 94822 491498 130586 491734
rect 130822 491498 166586 491734
rect 166822 491498 202586 491734
rect 202822 491498 238586 491734
rect 238822 491498 274586 491734
rect 274822 491498 310586 491734
rect 310822 491498 346586 491734
rect 346822 491498 382586 491734
rect 382822 491498 418586 491734
rect 418822 491498 454586 491734
rect 454822 491498 490586 491734
rect 490822 491498 526586 491734
rect 526822 491498 562586 491734
rect 562822 491498 588322 491734
rect 588558 491498 588740 491734
rect -4816 491476 588740 491498
rect -4816 491474 -4216 491476
rect 22404 491474 23004 491476
rect 58404 491474 59004 491476
rect 94404 491474 95004 491476
rect 130404 491474 131004 491476
rect 166404 491474 167004 491476
rect 202404 491474 203004 491476
rect 238404 491474 239004 491476
rect 274404 491474 275004 491476
rect 310404 491474 311004 491476
rect 346404 491474 347004 491476
rect 382404 491474 383004 491476
rect 418404 491474 419004 491476
rect 454404 491474 455004 491476
rect 490404 491474 491004 491476
rect 526404 491474 527004 491476
rect 562404 491474 563004 491476
rect 588140 491474 588740 491476
rect -2936 488476 -2336 488478
rect 18804 488476 19404 488478
rect 54804 488476 55404 488478
rect 90804 488476 91404 488478
rect 126804 488476 127404 488478
rect 162804 488476 163404 488478
rect 198804 488476 199404 488478
rect 234804 488476 235404 488478
rect 270804 488476 271404 488478
rect 306804 488476 307404 488478
rect 342804 488476 343404 488478
rect 378804 488476 379404 488478
rect 414804 488476 415404 488478
rect 450804 488476 451404 488478
rect 486804 488476 487404 488478
rect 522804 488476 523404 488478
rect 558804 488476 559404 488478
rect 586260 488476 586860 488478
rect -2936 488454 586860 488476
rect -2936 488218 -2754 488454
rect -2518 488218 18986 488454
rect 19222 488218 54986 488454
rect 55222 488218 90986 488454
rect 91222 488218 126986 488454
rect 127222 488218 162986 488454
rect 163222 488218 198986 488454
rect 199222 488218 234986 488454
rect 235222 488218 270986 488454
rect 271222 488218 306986 488454
rect 307222 488218 342986 488454
rect 343222 488218 378986 488454
rect 379222 488218 414986 488454
rect 415222 488218 450986 488454
rect 451222 488218 486986 488454
rect 487222 488218 522986 488454
rect 523222 488218 558986 488454
rect 559222 488218 586442 488454
rect 586678 488218 586860 488454
rect -2936 488134 586860 488218
rect -2936 487898 -2754 488134
rect -2518 487898 18986 488134
rect 19222 487898 54986 488134
rect 55222 487898 90986 488134
rect 91222 487898 126986 488134
rect 127222 487898 162986 488134
rect 163222 487898 198986 488134
rect 199222 487898 234986 488134
rect 235222 487898 270986 488134
rect 271222 487898 306986 488134
rect 307222 487898 342986 488134
rect 343222 487898 378986 488134
rect 379222 487898 414986 488134
rect 415222 487898 450986 488134
rect 451222 487898 486986 488134
rect 487222 487898 522986 488134
rect 523222 487898 558986 488134
rect 559222 487898 586442 488134
rect 586678 487898 586860 488134
rect -2936 487876 586860 487898
rect -2936 487874 -2336 487876
rect 18804 487874 19404 487876
rect 54804 487874 55404 487876
rect 90804 487874 91404 487876
rect 126804 487874 127404 487876
rect 162804 487874 163404 487876
rect 198804 487874 199404 487876
rect 234804 487874 235404 487876
rect 270804 487874 271404 487876
rect 306804 487874 307404 487876
rect 342804 487874 343404 487876
rect 378804 487874 379404 487876
rect 414804 487874 415404 487876
rect 450804 487874 451404 487876
rect 486804 487874 487404 487876
rect 522804 487874 523404 487876
rect 558804 487874 559404 487876
rect 586260 487874 586860 487876
rect -7636 481276 -7036 481278
rect 11604 481276 12204 481278
rect 47604 481276 48204 481278
rect 83604 481276 84204 481278
rect 119604 481276 120204 481278
rect 155604 481276 156204 481278
rect 191604 481276 192204 481278
rect 227604 481276 228204 481278
rect 263604 481276 264204 481278
rect 299604 481276 300204 481278
rect 335604 481276 336204 481278
rect 371604 481276 372204 481278
rect 407604 481276 408204 481278
rect 443604 481276 444204 481278
rect 479604 481276 480204 481278
rect 515604 481276 516204 481278
rect 551604 481276 552204 481278
rect 590960 481276 591560 481278
rect -8576 481254 592500 481276
rect -8576 481018 -7454 481254
rect -7218 481018 11786 481254
rect 12022 481018 47786 481254
rect 48022 481018 83786 481254
rect 84022 481018 119786 481254
rect 120022 481018 155786 481254
rect 156022 481018 191786 481254
rect 192022 481018 227786 481254
rect 228022 481018 263786 481254
rect 264022 481018 299786 481254
rect 300022 481018 335786 481254
rect 336022 481018 371786 481254
rect 372022 481018 407786 481254
rect 408022 481018 443786 481254
rect 444022 481018 479786 481254
rect 480022 481018 515786 481254
rect 516022 481018 551786 481254
rect 552022 481018 591142 481254
rect 591378 481018 592500 481254
rect -8576 480934 592500 481018
rect -8576 480698 -7454 480934
rect -7218 480698 11786 480934
rect 12022 480698 47786 480934
rect 48022 480698 83786 480934
rect 84022 480698 119786 480934
rect 120022 480698 155786 480934
rect 156022 480698 191786 480934
rect 192022 480698 227786 480934
rect 228022 480698 263786 480934
rect 264022 480698 299786 480934
rect 300022 480698 335786 480934
rect 336022 480698 371786 480934
rect 372022 480698 407786 480934
rect 408022 480698 443786 480934
rect 444022 480698 479786 480934
rect 480022 480698 515786 480934
rect 516022 480698 551786 480934
rect 552022 480698 591142 480934
rect 591378 480698 592500 480934
rect -8576 480676 592500 480698
rect -7636 480674 -7036 480676
rect 11604 480674 12204 480676
rect 47604 480674 48204 480676
rect 83604 480674 84204 480676
rect 119604 480674 120204 480676
rect 155604 480674 156204 480676
rect 191604 480674 192204 480676
rect 227604 480674 228204 480676
rect 263604 480674 264204 480676
rect 299604 480674 300204 480676
rect 335604 480674 336204 480676
rect 371604 480674 372204 480676
rect 407604 480674 408204 480676
rect 443604 480674 444204 480676
rect 479604 480674 480204 480676
rect 515604 480674 516204 480676
rect 551604 480674 552204 480676
rect 590960 480674 591560 480676
rect -5756 477676 -5156 477678
rect 8004 477676 8604 477678
rect 44004 477676 44604 477678
rect 80004 477676 80604 477678
rect 116004 477676 116604 477678
rect 152004 477676 152604 477678
rect 188004 477676 188604 477678
rect 224004 477676 224604 477678
rect 260004 477676 260604 477678
rect 296004 477676 296604 477678
rect 332004 477676 332604 477678
rect 368004 477676 368604 477678
rect 404004 477676 404604 477678
rect 440004 477676 440604 477678
rect 476004 477676 476604 477678
rect 512004 477676 512604 477678
rect 548004 477676 548604 477678
rect 589080 477676 589680 477678
rect -6696 477654 590620 477676
rect -6696 477418 -5574 477654
rect -5338 477418 8186 477654
rect 8422 477418 44186 477654
rect 44422 477418 80186 477654
rect 80422 477418 116186 477654
rect 116422 477418 152186 477654
rect 152422 477418 188186 477654
rect 188422 477418 224186 477654
rect 224422 477418 260186 477654
rect 260422 477418 296186 477654
rect 296422 477418 332186 477654
rect 332422 477418 368186 477654
rect 368422 477418 404186 477654
rect 404422 477418 440186 477654
rect 440422 477418 476186 477654
rect 476422 477418 512186 477654
rect 512422 477418 548186 477654
rect 548422 477418 589262 477654
rect 589498 477418 590620 477654
rect -6696 477334 590620 477418
rect -6696 477098 -5574 477334
rect -5338 477098 8186 477334
rect 8422 477098 44186 477334
rect 44422 477098 80186 477334
rect 80422 477098 116186 477334
rect 116422 477098 152186 477334
rect 152422 477098 188186 477334
rect 188422 477098 224186 477334
rect 224422 477098 260186 477334
rect 260422 477098 296186 477334
rect 296422 477098 332186 477334
rect 332422 477098 368186 477334
rect 368422 477098 404186 477334
rect 404422 477098 440186 477334
rect 440422 477098 476186 477334
rect 476422 477098 512186 477334
rect 512422 477098 548186 477334
rect 548422 477098 589262 477334
rect 589498 477098 590620 477334
rect -6696 477076 590620 477098
rect -5756 477074 -5156 477076
rect 8004 477074 8604 477076
rect 44004 477074 44604 477076
rect 80004 477074 80604 477076
rect 116004 477074 116604 477076
rect 152004 477074 152604 477076
rect 188004 477074 188604 477076
rect 224004 477074 224604 477076
rect 260004 477074 260604 477076
rect 296004 477074 296604 477076
rect 332004 477074 332604 477076
rect 368004 477074 368604 477076
rect 404004 477074 404604 477076
rect 440004 477074 440604 477076
rect 476004 477074 476604 477076
rect 512004 477074 512604 477076
rect 548004 477074 548604 477076
rect 589080 477074 589680 477076
rect -3876 474076 -3276 474078
rect 4404 474076 5004 474078
rect 40404 474076 41004 474078
rect 76404 474076 77004 474078
rect 112404 474076 113004 474078
rect 148404 474076 149004 474078
rect 184404 474076 185004 474078
rect 220404 474076 221004 474078
rect 256404 474076 257004 474078
rect 292404 474076 293004 474078
rect 328404 474076 329004 474078
rect 364404 474076 365004 474078
rect 400404 474076 401004 474078
rect 436404 474076 437004 474078
rect 472404 474076 473004 474078
rect 508404 474076 509004 474078
rect 544404 474076 545004 474078
rect 580404 474076 581004 474078
rect 587200 474076 587800 474078
rect -4816 474054 588740 474076
rect -4816 473818 -3694 474054
rect -3458 473818 4586 474054
rect 4822 473818 40586 474054
rect 40822 473818 76586 474054
rect 76822 473818 112586 474054
rect 112822 473818 148586 474054
rect 148822 473818 184586 474054
rect 184822 473818 220586 474054
rect 220822 473818 256586 474054
rect 256822 473818 292586 474054
rect 292822 473818 328586 474054
rect 328822 473818 364586 474054
rect 364822 473818 400586 474054
rect 400822 473818 436586 474054
rect 436822 473818 472586 474054
rect 472822 473818 508586 474054
rect 508822 473818 544586 474054
rect 544822 473818 580586 474054
rect 580822 473818 587382 474054
rect 587618 473818 588740 474054
rect -4816 473734 588740 473818
rect -4816 473498 -3694 473734
rect -3458 473498 4586 473734
rect 4822 473498 40586 473734
rect 40822 473498 76586 473734
rect 76822 473498 112586 473734
rect 112822 473498 148586 473734
rect 148822 473498 184586 473734
rect 184822 473498 220586 473734
rect 220822 473498 256586 473734
rect 256822 473498 292586 473734
rect 292822 473498 328586 473734
rect 328822 473498 364586 473734
rect 364822 473498 400586 473734
rect 400822 473498 436586 473734
rect 436822 473498 472586 473734
rect 472822 473498 508586 473734
rect 508822 473498 544586 473734
rect 544822 473498 580586 473734
rect 580822 473498 587382 473734
rect 587618 473498 588740 473734
rect -4816 473476 588740 473498
rect -3876 473474 -3276 473476
rect 4404 473474 5004 473476
rect 40404 473474 41004 473476
rect 76404 473474 77004 473476
rect 112404 473474 113004 473476
rect 148404 473474 149004 473476
rect 184404 473474 185004 473476
rect 220404 473474 221004 473476
rect 256404 473474 257004 473476
rect 292404 473474 293004 473476
rect 328404 473474 329004 473476
rect 364404 473474 365004 473476
rect 400404 473474 401004 473476
rect 436404 473474 437004 473476
rect 472404 473474 473004 473476
rect 508404 473474 509004 473476
rect 544404 473474 545004 473476
rect 580404 473474 581004 473476
rect 587200 473474 587800 473476
rect -1996 470476 -1396 470478
rect 804 470476 1404 470478
rect 36804 470476 37404 470478
rect 72804 470476 73404 470478
rect 108804 470476 109404 470478
rect 144804 470476 145404 470478
rect 180804 470476 181404 470478
rect 216804 470476 217404 470478
rect 252804 470476 253404 470478
rect 288804 470476 289404 470478
rect 324804 470476 325404 470478
rect 360804 470476 361404 470478
rect 396804 470476 397404 470478
rect 432804 470476 433404 470478
rect 468804 470476 469404 470478
rect 504804 470476 505404 470478
rect 540804 470476 541404 470478
rect 576804 470476 577404 470478
rect 585320 470476 585920 470478
rect -2936 470454 586860 470476
rect -2936 470218 -1814 470454
rect -1578 470218 986 470454
rect 1222 470218 36986 470454
rect 37222 470218 72986 470454
rect 73222 470218 108986 470454
rect 109222 470218 144986 470454
rect 145222 470218 180986 470454
rect 181222 470218 216986 470454
rect 217222 470218 252986 470454
rect 253222 470218 288986 470454
rect 289222 470218 324986 470454
rect 325222 470218 360986 470454
rect 361222 470218 396986 470454
rect 397222 470218 432986 470454
rect 433222 470218 468986 470454
rect 469222 470218 504986 470454
rect 505222 470218 540986 470454
rect 541222 470218 576986 470454
rect 577222 470218 585502 470454
rect 585738 470218 586860 470454
rect -2936 470134 586860 470218
rect -2936 469898 -1814 470134
rect -1578 469898 986 470134
rect 1222 469898 36986 470134
rect 37222 469898 72986 470134
rect 73222 469898 108986 470134
rect 109222 469898 144986 470134
rect 145222 469898 180986 470134
rect 181222 469898 216986 470134
rect 217222 469898 252986 470134
rect 253222 469898 288986 470134
rect 289222 469898 324986 470134
rect 325222 469898 360986 470134
rect 361222 469898 396986 470134
rect 397222 469898 432986 470134
rect 433222 469898 468986 470134
rect 469222 469898 504986 470134
rect 505222 469898 540986 470134
rect 541222 469898 576986 470134
rect 577222 469898 585502 470134
rect 585738 469898 586860 470134
rect -2936 469876 586860 469898
rect -1996 469874 -1396 469876
rect 804 469874 1404 469876
rect 36804 469874 37404 469876
rect 72804 469874 73404 469876
rect 108804 469874 109404 469876
rect 144804 469874 145404 469876
rect 180804 469874 181404 469876
rect 216804 469874 217404 469876
rect 252804 469874 253404 469876
rect 288804 469874 289404 469876
rect 324804 469874 325404 469876
rect 360804 469874 361404 469876
rect 396804 469874 397404 469876
rect 432804 469874 433404 469876
rect 468804 469874 469404 469876
rect 504804 469874 505404 469876
rect 540804 469874 541404 469876
rect 576804 469874 577404 469876
rect 585320 469874 585920 469876
rect -8576 463276 -7976 463278
rect 29604 463276 30204 463278
rect 65604 463276 66204 463278
rect 101604 463276 102204 463278
rect 137604 463276 138204 463278
rect 173604 463276 174204 463278
rect 209604 463276 210204 463278
rect 245604 463276 246204 463278
rect 281604 463276 282204 463278
rect 317604 463276 318204 463278
rect 353604 463276 354204 463278
rect 389604 463276 390204 463278
rect 425604 463276 426204 463278
rect 461604 463276 462204 463278
rect 497604 463276 498204 463278
rect 533604 463276 534204 463278
rect 569604 463276 570204 463278
rect 591900 463276 592500 463278
rect -8576 463254 592500 463276
rect -8576 463018 -8394 463254
rect -8158 463018 29786 463254
rect 30022 463018 65786 463254
rect 66022 463018 101786 463254
rect 102022 463018 137786 463254
rect 138022 463018 173786 463254
rect 174022 463018 209786 463254
rect 210022 463018 245786 463254
rect 246022 463018 281786 463254
rect 282022 463018 317786 463254
rect 318022 463018 353786 463254
rect 354022 463018 389786 463254
rect 390022 463018 425786 463254
rect 426022 463018 461786 463254
rect 462022 463018 497786 463254
rect 498022 463018 533786 463254
rect 534022 463018 569786 463254
rect 570022 463018 592082 463254
rect 592318 463018 592500 463254
rect -8576 462934 592500 463018
rect -8576 462698 -8394 462934
rect -8158 462698 29786 462934
rect 30022 462698 65786 462934
rect 66022 462698 101786 462934
rect 102022 462698 137786 462934
rect 138022 462698 173786 462934
rect 174022 462698 209786 462934
rect 210022 462698 245786 462934
rect 246022 462698 281786 462934
rect 282022 462698 317786 462934
rect 318022 462698 353786 462934
rect 354022 462698 389786 462934
rect 390022 462698 425786 462934
rect 426022 462698 461786 462934
rect 462022 462698 497786 462934
rect 498022 462698 533786 462934
rect 534022 462698 569786 462934
rect 570022 462698 592082 462934
rect 592318 462698 592500 462934
rect -8576 462676 592500 462698
rect -8576 462674 -7976 462676
rect 29604 462674 30204 462676
rect 65604 462674 66204 462676
rect 101604 462674 102204 462676
rect 137604 462674 138204 462676
rect 173604 462674 174204 462676
rect 209604 462674 210204 462676
rect 245604 462674 246204 462676
rect 281604 462674 282204 462676
rect 317604 462674 318204 462676
rect 353604 462674 354204 462676
rect 389604 462674 390204 462676
rect 425604 462674 426204 462676
rect 461604 462674 462204 462676
rect 497604 462674 498204 462676
rect 533604 462674 534204 462676
rect 569604 462674 570204 462676
rect 591900 462674 592500 462676
rect -6696 459676 -6096 459678
rect 26004 459676 26604 459678
rect 62004 459676 62604 459678
rect 98004 459676 98604 459678
rect 134004 459676 134604 459678
rect 170004 459676 170604 459678
rect 206004 459676 206604 459678
rect 242004 459676 242604 459678
rect 278004 459676 278604 459678
rect 314004 459676 314604 459678
rect 350004 459676 350604 459678
rect 386004 459676 386604 459678
rect 422004 459676 422604 459678
rect 458004 459676 458604 459678
rect 494004 459676 494604 459678
rect 530004 459676 530604 459678
rect 566004 459676 566604 459678
rect 590020 459676 590620 459678
rect -6696 459654 590620 459676
rect -6696 459418 -6514 459654
rect -6278 459418 26186 459654
rect 26422 459418 62186 459654
rect 62422 459418 98186 459654
rect 98422 459418 134186 459654
rect 134422 459418 170186 459654
rect 170422 459418 206186 459654
rect 206422 459418 242186 459654
rect 242422 459418 278186 459654
rect 278422 459418 314186 459654
rect 314422 459418 350186 459654
rect 350422 459418 386186 459654
rect 386422 459418 422186 459654
rect 422422 459418 458186 459654
rect 458422 459418 494186 459654
rect 494422 459418 530186 459654
rect 530422 459418 566186 459654
rect 566422 459418 590202 459654
rect 590438 459418 590620 459654
rect -6696 459334 590620 459418
rect -6696 459098 -6514 459334
rect -6278 459098 26186 459334
rect 26422 459098 62186 459334
rect 62422 459098 98186 459334
rect 98422 459098 134186 459334
rect 134422 459098 170186 459334
rect 170422 459098 206186 459334
rect 206422 459098 242186 459334
rect 242422 459098 278186 459334
rect 278422 459098 314186 459334
rect 314422 459098 350186 459334
rect 350422 459098 386186 459334
rect 386422 459098 422186 459334
rect 422422 459098 458186 459334
rect 458422 459098 494186 459334
rect 494422 459098 530186 459334
rect 530422 459098 566186 459334
rect 566422 459098 590202 459334
rect 590438 459098 590620 459334
rect -6696 459076 590620 459098
rect -6696 459074 -6096 459076
rect 26004 459074 26604 459076
rect 62004 459074 62604 459076
rect 98004 459074 98604 459076
rect 134004 459074 134604 459076
rect 170004 459074 170604 459076
rect 206004 459074 206604 459076
rect 242004 459074 242604 459076
rect 278004 459074 278604 459076
rect 314004 459074 314604 459076
rect 350004 459074 350604 459076
rect 386004 459074 386604 459076
rect 422004 459074 422604 459076
rect 458004 459074 458604 459076
rect 494004 459074 494604 459076
rect 530004 459074 530604 459076
rect 566004 459074 566604 459076
rect 590020 459074 590620 459076
rect -4816 456076 -4216 456078
rect 22404 456076 23004 456078
rect 58404 456076 59004 456078
rect 94404 456076 95004 456078
rect 130404 456076 131004 456078
rect 166404 456076 167004 456078
rect 202404 456076 203004 456078
rect 238404 456076 239004 456078
rect 274404 456076 275004 456078
rect 310404 456076 311004 456078
rect 346404 456076 347004 456078
rect 382404 456076 383004 456078
rect 418404 456076 419004 456078
rect 454404 456076 455004 456078
rect 490404 456076 491004 456078
rect 526404 456076 527004 456078
rect 562404 456076 563004 456078
rect 588140 456076 588740 456078
rect -4816 456054 588740 456076
rect -4816 455818 -4634 456054
rect -4398 455818 22586 456054
rect 22822 455818 58586 456054
rect 58822 455818 94586 456054
rect 94822 455818 130586 456054
rect 130822 455818 166586 456054
rect 166822 455818 202586 456054
rect 202822 455818 238586 456054
rect 238822 455818 274586 456054
rect 274822 455818 310586 456054
rect 310822 455818 346586 456054
rect 346822 455818 382586 456054
rect 382822 455818 418586 456054
rect 418822 455818 454586 456054
rect 454822 455818 490586 456054
rect 490822 455818 526586 456054
rect 526822 455818 562586 456054
rect 562822 455818 588322 456054
rect 588558 455818 588740 456054
rect -4816 455734 588740 455818
rect -4816 455498 -4634 455734
rect -4398 455498 22586 455734
rect 22822 455498 58586 455734
rect 58822 455498 94586 455734
rect 94822 455498 130586 455734
rect 130822 455498 166586 455734
rect 166822 455498 202586 455734
rect 202822 455498 238586 455734
rect 238822 455498 274586 455734
rect 274822 455498 310586 455734
rect 310822 455498 346586 455734
rect 346822 455498 382586 455734
rect 382822 455498 418586 455734
rect 418822 455498 454586 455734
rect 454822 455498 490586 455734
rect 490822 455498 526586 455734
rect 526822 455498 562586 455734
rect 562822 455498 588322 455734
rect 588558 455498 588740 455734
rect -4816 455476 588740 455498
rect -4816 455474 -4216 455476
rect 22404 455474 23004 455476
rect 58404 455474 59004 455476
rect 94404 455474 95004 455476
rect 130404 455474 131004 455476
rect 166404 455474 167004 455476
rect 202404 455474 203004 455476
rect 238404 455474 239004 455476
rect 274404 455474 275004 455476
rect 310404 455474 311004 455476
rect 346404 455474 347004 455476
rect 382404 455474 383004 455476
rect 418404 455474 419004 455476
rect 454404 455474 455004 455476
rect 490404 455474 491004 455476
rect 526404 455474 527004 455476
rect 562404 455474 563004 455476
rect 588140 455474 588740 455476
rect -2936 452476 -2336 452478
rect 18804 452476 19404 452478
rect 54804 452476 55404 452478
rect 90804 452476 91404 452478
rect 126804 452476 127404 452478
rect 162804 452476 163404 452478
rect 198804 452476 199404 452478
rect 234804 452476 235404 452478
rect 270804 452476 271404 452478
rect 306804 452476 307404 452478
rect 342804 452476 343404 452478
rect 378804 452476 379404 452478
rect 414804 452476 415404 452478
rect 450804 452476 451404 452478
rect 486804 452476 487404 452478
rect 522804 452476 523404 452478
rect 558804 452476 559404 452478
rect 586260 452476 586860 452478
rect -2936 452454 586860 452476
rect -2936 452218 -2754 452454
rect -2518 452218 18986 452454
rect 19222 452218 54986 452454
rect 55222 452218 90986 452454
rect 91222 452218 126986 452454
rect 127222 452218 162986 452454
rect 163222 452218 198986 452454
rect 199222 452218 234986 452454
rect 235222 452218 270986 452454
rect 271222 452218 306986 452454
rect 307222 452218 342986 452454
rect 343222 452218 378986 452454
rect 379222 452218 414986 452454
rect 415222 452218 450986 452454
rect 451222 452218 486986 452454
rect 487222 452218 522986 452454
rect 523222 452218 558986 452454
rect 559222 452218 586442 452454
rect 586678 452218 586860 452454
rect -2936 452134 586860 452218
rect -2936 451898 -2754 452134
rect -2518 451898 18986 452134
rect 19222 451898 54986 452134
rect 55222 451898 90986 452134
rect 91222 451898 126986 452134
rect 127222 451898 162986 452134
rect 163222 451898 198986 452134
rect 199222 451898 234986 452134
rect 235222 451898 270986 452134
rect 271222 451898 306986 452134
rect 307222 451898 342986 452134
rect 343222 451898 378986 452134
rect 379222 451898 414986 452134
rect 415222 451898 450986 452134
rect 451222 451898 486986 452134
rect 487222 451898 522986 452134
rect 523222 451898 558986 452134
rect 559222 451898 586442 452134
rect 586678 451898 586860 452134
rect -2936 451876 586860 451898
rect -2936 451874 -2336 451876
rect 18804 451874 19404 451876
rect 54804 451874 55404 451876
rect 90804 451874 91404 451876
rect 126804 451874 127404 451876
rect 162804 451874 163404 451876
rect 198804 451874 199404 451876
rect 234804 451874 235404 451876
rect 270804 451874 271404 451876
rect 306804 451874 307404 451876
rect 342804 451874 343404 451876
rect 378804 451874 379404 451876
rect 414804 451874 415404 451876
rect 450804 451874 451404 451876
rect 486804 451874 487404 451876
rect 522804 451874 523404 451876
rect 558804 451874 559404 451876
rect 586260 451874 586860 451876
rect -7636 445276 -7036 445278
rect 11604 445276 12204 445278
rect 47604 445276 48204 445278
rect 83604 445276 84204 445278
rect 119604 445276 120204 445278
rect 155604 445276 156204 445278
rect 191604 445276 192204 445278
rect 227604 445276 228204 445278
rect 263604 445276 264204 445278
rect 299604 445276 300204 445278
rect 335604 445276 336204 445278
rect 371604 445276 372204 445278
rect 407604 445276 408204 445278
rect 443604 445276 444204 445278
rect 479604 445276 480204 445278
rect 515604 445276 516204 445278
rect 551604 445276 552204 445278
rect 590960 445276 591560 445278
rect -8576 445254 592500 445276
rect -8576 445018 -7454 445254
rect -7218 445018 11786 445254
rect 12022 445018 47786 445254
rect 48022 445018 83786 445254
rect 84022 445018 119786 445254
rect 120022 445018 155786 445254
rect 156022 445018 191786 445254
rect 192022 445018 227786 445254
rect 228022 445018 263786 445254
rect 264022 445018 299786 445254
rect 300022 445018 335786 445254
rect 336022 445018 371786 445254
rect 372022 445018 407786 445254
rect 408022 445018 443786 445254
rect 444022 445018 479786 445254
rect 480022 445018 515786 445254
rect 516022 445018 551786 445254
rect 552022 445018 591142 445254
rect 591378 445018 592500 445254
rect -8576 444934 592500 445018
rect -8576 444698 -7454 444934
rect -7218 444698 11786 444934
rect 12022 444698 47786 444934
rect 48022 444698 83786 444934
rect 84022 444698 119786 444934
rect 120022 444698 155786 444934
rect 156022 444698 191786 444934
rect 192022 444698 227786 444934
rect 228022 444698 263786 444934
rect 264022 444698 299786 444934
rect 300022 444698 335786 444934
rect 336022 444698 371786 444934
rect 372022 444698 407786 444934
rect 408022 444698 443786 444934
rect 444022 444698 479786 444934
rect 480022 444698 515786 444934
rect 516022 444698 551786 444934
rect 552022 444698 591142 444934
rect 591378 444698 592500 444934
rect -8576 444676 592500 444698
rect -7636 444674 -7036 444676
rect 11604 444674 12204 444676
rect 47604 444674 48204 444676
rect 83604 444674 84204 444676
rect 119604 444674 120204 444676
rect 155604 444674 156204 444676
rect 191604 444674 192204 444676
rect 227604 444674 228204 444676
rect 263604 444674 264204 444676
rect 299604 444674 300204 444676
rect 335604 444674 336204 444676
rect 371604 444674 372204 444676
rect 407604 444674 408204 444676
rect 443604 444674 444204 444676
rect 479604 444674 480204 444676
rect 515604 444674 516204 444676
rect 551604 444674 552204 444676
rect 590960 444674 591560 444676
rect -5756 441676 -5156 441678
rect 8004 441676 8604 441678
rect 44004 441676 44604 441678
rect 80004 441676 80604 441678
rect 116004 441676 116604 441678
rect 152004 441676 152604 441678
rect 188004 441676 188604 441678
rect 224004 441676 224604 441678
rect 260004 441676 260604 441678
rect 296004 441676 296604 441678
rect 332004 441676 332604 441678
rect 368004 441676 368604 441678
rect 404004 441676 404604 441678
rect 440004 441676 440604 441678
rect 476004 441676 476604 441678
rect 512004 441676 512604 441678
rect 548004 441676 548604 441678
rect 589080 441676 589680 441678
rect -6696 441654 590620 441676
rect -6696 441418 -5574 441654
rect -5338 441418 8186 441654
rect 8422 441418 44186 441654
rect 44422 441418 80186 441654
rect 80422 441418 116186 441654
rect 116422 441418 152186 441654
rect 152422 441418 188186 441654
rect 188422 441418 224186 441654
rect 224422 441418 260186 441654
rect 260422 441418 296186 441654
rect 296422 441418 332186 441654
rect 332422 441418 368186 441654
rect 368422 441418 404186 441654
rect 404422 441418 440186 441654
rect 440422 441418 476186 441654
rect 476422 441418 512186 441654
rect 512422 441418 548186 441654
rect 548422 441418 589262 441654
rect 589498 441418 590620 441654
rect -6696 441334 590620 441418
rect -6696 441098 -5574 441334
rect -5338 441098 8186 441334
rect 8422 441098 44186 441334
rect 44422 441098 80186 441334
rect 80422 441098 116186 441334
rect 116422 441098 152186 441334
rect 152422 441098 188186 441334
rect 188422 441098 224186 441334
rect 224422 441098 260186 441334
rect 260422 441098 296186 441334
rect 296422 441098 332186 441334
rect 332422 441098 368186 441334
rect 368422 441098 404186 441334
rect 404422 441098 440186 441334
rect 440422 441098 476186 441334
rect 476422 441098 512186 441334
rect 512422 441098 548186 441334
rect 548422 441098 589262 441334
rect 589498 441098 590620 441334
rect -6696 441076 590620 441098
rect -5756 441074 -5156 441076
rect 8004 441074 8604 441076
rect 44004 441074 44604 441076
rect 80004 441074 80604 441076
rect 116004 441074 116604 441076
rect 152004 441074 152604 441076
rect 188004 441074 188604 441076
rect 224004 441074 224604 441076
rect 260004 441074 260604 441076
rect 296004 441074 296604 441076
rect 332004 441074 332604 441076
rect 368004 441074 368604 441076
rect 404004 441074 404604 441076
rect 440004 441074 440604 441076
rect 476004 441074 476604 441076
rect 512004 441074 512604 441076
rect 548004 441074 548604 441076
rect 589080 441074 589680 441076
rect -3876 438076 -3276 438078
rect 4404 438076 5004 438078
rect 40404 438076 41004 438078
rect 76404 438076 77004 438078
rect 112404 438076 113004 438078
rect 148404 438076 149004 438078
rect 184404 438076 185004 438078
rect 220404 438076 221004 438078
rect 256404 438076 257004 438078
rect 292404 438076 293004 438078
rect 328404 438076 329004 438078
rect 364404 438076 365004 438078
rect 400404 438076 401004 438078
rect 436404 438076 437004 438078
rect 472404 438076 473004 438078
rect 508404 438076 509004 438078
rect 544404 438076 545004 438078
rect 580404 438076 581004 438078
rect 587200 438076 587800 438078
rect -4816 438054 588740 438076
rect -4816 437818 -3694 438054
rect -3458 437818 4586 438054
rect 4822 437818 40586 438054
rect 40822 437818 76586 438054
rect 76822 437818 112586 438054
rect 112822 437818 148586 438054
rect 148822 437818 184586 438054
rect 184822 437818 220586 438054
rect 220822 437818 256586 438054
rect 256822 437818 292586 438054
rect 292822 437818 328586 438054
rect 328822 437818 364586 438054
rect 364822 437818 400586 438054
rect 400822 437818 436586 438054
rect 436822 437818 472586 438054
rect 472822 437818 508586 438054
rect 508822 437818 544586 438054
rect 544822 437818 580586 438054
rect 580822 437818 587382 438054
rect 587618 437818 588740 438054
rect -4816 437734 588740 437818
rect -4816 437498 -3694 437734
rect -3458 437498 4586 437734
rect 4822 437498 40586 437734
rect 40822 437498 76586 437734
rect 76822 437498 112586 437734
rect 112822 437498 148586 437734
rect 148822 437498 184586 437734
rect 184822 437498 220586 437734
rect 220822 437498 256586 437734
rect 256822 437498 292586 437734
rect 292822 437498 328586 437734
rect 328822 437498 364586 437734
rect 364822 437498 400586 437734
rect 400822 437498 436586 437734
rect 436822 437498 472586 437734
rect 472822 437498 508586 437734
rect 508822 437498 544586 437734
rect 544822 437498 580586 437734
rect 580822 437498 587382 437734
rect 587618 437498 588740 437734
rect -4816 437476 588740 437498
rect -3876 437474 -3276 437476
rect 4404 437474 5004 437476
rect 40404 437474 41004 437476
rect 76404 437474 77004 437476
rect 112404 437474 113004 437476
rect 148404 437474 149004 437476
rect 184404 437474 185004 437476
rect 220404 437474 221004 437476
rect 256404 437474 257004 437476
rect 292404 437474 293004 437476
rect 328404 437474 329004 437476
rect 364404 437474 365004 437476
rect 400404 437474 401004 437476
rect 436404 437474 437004 437476
rect 472404 437474 473004 437476
rect 508404 437474 509004 437476
rect 544404 437474 545004 437476
rect 580404 437474 581004 437476
rect 587200 437474 587800 437476
rect -1996 434476 -1396 434478
rect 804 434476 1404 434478
rect 36804 434476 37404 434478
rect 72804 434476 73404 434478
rect 108804 434476 109404 434478
rect 144804 434476 145404 434478
rect 180804 434476 181404 434478
rect 216804 434476 217404 434478
rect 252804 434476 253404 434478
rect 288804 434476 289404 434478
rect 324804 434476 325404 434478
rect 360804 434476 361404 434478
rect 396804 434476 397404 434478
rect 432804 434476 433404 434478
rect 468804 434476 469404 434478
rect 504804 434476 505404 434478
rect 540804 434476 541404 434478
rect 576804 434476 577404 434478
rect 585320 434476 585920 434478
rect -2936 434454 586860 434476
rect -2936 434218 -1814 434454
rect -1578 434218 986 434454
rect 1222 434218 36986 434454
rect 37222 434218 72986 434454
rect 73222 434218 108986 434454
rect 109222 434218 144986 434454
rect 145222 434218 180986 434454
rect 181222 434218 216986 434454
rect 217222 434218 252986 434454
rect 253222 434218 288986 434454
rect 289222 434218 324986 434454
rect 325222 434218 360986 434454
rect 361222 434218 396986 434454
rect 397222 434218 432986 434454
rect 433222 434218 468986 434454
rect 469222 434218 504986 434454
rect 505222 434218 540986 434454
rect 541222 434218 576986 434454
rect 577222 434218 585502 434454
rect 585738 434218 586860 434454
rect -2936 434134 586860 434218
rect -2936 433898 -1814 434134
rect -1578 433898 986 434134
rect 1222 433898 36986 434134
rect 37222 433898 72986 434134
rect 73222 433898 108986 434134
rect 109222 433898 144986 434134
rect 145222 433898 180986 434134
rect 181222 433898 216986 434134
rect 217222 433898 252986 434134
rect 253222 433898 288986 434134
rect 289222 433898 324986 434134
rect 325222 433898 360986 434134
rect 361222 433898 396986 434134
rect 397222 433898 432986 434134
rect 433222 433898 468986 434134
rect 469222 433898 504986 434134
rect 505222 433898 540986 434134
rect 541222 433898 576986 434134
rect 577222 433898 585502 434134
rect 585738 433898 586860 434134
rect -2936 433876 586860 433898
rect -1996 433874 -1396 433876
rect 804 433874 1404 433876
rect 36804 433874 37404 433876
rect 72804 433874 73404 433876
rect 108804 433874 109404 433876
rect 144804 433874 145404 433876
rect 180804 433874 181404 433876
rect 216804 433874 217404 433876
rect 252804 433874 253404 433876
rect 288804 433874 289404 433876
rect 324804 433874 325404 433876
rect 360804 433874 361404 433876
rect 396804 433874 397404 433876
rect 432804 433874 433404 433876
rect 468804 433874 469404 433876
rect 504804 433874 505404 433876
rect 540804 433874 541404 433876
rect 576804 433874 577404 433876
rect 585320 433874 585920 433876
rect -8576 427276 -7976 427278
rect 29604 427276 30204 427278
rect 65604 427276 66204 427278
rect 101604 427276 102204 427278
rect 137604 427276 138204 427278
rect 173604 427276 174204 427278
rect 209604 427276 210204 427278
rect 245604 427276 246204 427278
rect 281604 427276 282204 427278
rect 317604 427276 318204 427278
rect 353604 427276 354204 427278
rect 389604 427276 390204 427278
rect 425604 427276 426204 427278
rect 461604 427276 462204 427278
rect 497604 427276 498204 427278
rect 533604 427276 534204 427278
rect 569604 427276 570204 427278
rect 591900 427276 592500 427278
rect -8576 427254 592500 427276
rect -8576 427018 -8394 427254
rect -8158 427018 29786 427254
rect 30022 427018 65786 427254
rect 66022 427018 101786 427254
rect 102022 427018 137786 427254
rect 138022 427018 173786 427254
rect 174022 427018 209786 427254
rect 210022 427018 245786 427254
rect 246022 427018 281786 427254
rect 282022 427018 317786 427254
rect 318022 427018 353786 427254
rect 354022 427018 389786 427254
rect 390022 427018 425786 427254
rect 426022 427018 461786 427254
rect 462022 427018 497786 427254
rect 498022 427018 533786 427254
rect 534022 427018 569786 427254
rect 570022 427018 592082 427254
rect 592318 427018 592500 427254
rect -8576 426934 592500 427018
rect -8576 426698 -8394 426934
rect -8158 426698 29786 426934
rect 30022 426698 65786 426934
rect 66022 426698 101786 426934
rect 102022 426698 137786 426934
rect 138022 426698 173786 426934
rect 174022 426698 209786 426934
rect 210022 426698 245786 426934
rect 246022 426698 281786 426934
rect 282022 426698 317786 426934
rect 318022 426698 353786 426934
rect 354022 426698 389786 426934
rect 390022 426698 425786 426934
rect 426022 426698 461786 426934
rect 462022 426698 497786 426934
rect 498022 426698 533786 426934
rect 534022 426698 569786 426934
rect 570022 426698 592082 426934
rect 592318 426698 592500 426934
rect -8576 426676 592500 426698
rect -8576 426674 -7976 426676
rect 29604 426674 30204 426676
rect 65604 426674 66204 426676
rect 101604 426674 102204 426676
rect 137604 426674 138204 426676
rect 173604 426674 174204 426676
rect 209604 426674 210204 426676
rect 245604 426674 246204 426676
rect 281604 426674 282204 426676
rect 317604 426674 318204 426676
rect 353604 426674 354204 426676
rect 389604 426674 390204 426676
rect 425604 426674 426204 426676
rect 461604 426674 462204 426676
rect 497604 426674 498204 426676
rect 533604 426674 534204 426676
rect 569604 426674 570204 426676
rect 591900 426674 592500 426676
rect -6696 423676 -6096 423678
rect 26004 423676 26604 423678
rect 62004 423676 62604 423678
rect 98004 423676 98604 423678
rect 134004 423676 134604 423678
rect 170004 423676 170604 423678
rect 206004 423676 206604 423678
rect 242004 423676 242604 423678
rect 278004 423676 278604 423678
rect 314004 423676 314604 423678
rect 350004 423676 350604 423678
rect 386004 423676 386604 423678
rect 422004 423676 422604 423678
rect 458004 423676 458604 423678
rect 494004 423676 494604 423678
rect 530004 423676 530604 423678
rect 566004 423676 566604 423678
rect 590020 423676 590620 423678
rect -6696 423654 590620 423676
rect -6696 423418 -6514 423654
rect -6278 423418 26186 423654
rect 26422 423418 62186 423654
rect 62422 423418 98186 423654
rect 98422 423418 134186 423654
rect 134422 423418 170186 423654
rect 170422 423418 206186 423654
rect 206422 423418 242186 423654
rect 242422 423418 278186 423654
rect 278422 423418 314186 423654
rect 314422 423418 350186 423654
rect 350422 423418 386186 423654
rect 386422 423418 422186 423654
rect 422422 423418 458186 423654
rect 458422 423418 494186 423654
rect 494422 423418 530186 423654
rect 530422 423418 566186 423654
rect 566422 423418 590202 423654
rect 590438 423418 590620 423654
rect -6696 423334 590620 423418
rect -6696 423098 -6514 423334
rect -6278 423098 26186 423334
rect 26422 423098 62186 423334
rect 62422 423098 98186 423334
rect 98422 423098 134186 423334
rect 134422 423098 170186 423334
rect 170422 423098 206186 423334
rect 206422 423098 242186 423334
rect 242422 423098 278186 423334
rect 278422 423098 314186 423334
rect 314422 423098 350186 423334
rect 350422 423098 386186 423334
rect 386422 423098 422186 423334
rect 422422 423098 458186 423334
rect 458422 423098 494186 423334
rect 494422 423098 530186 423334
rect 530422 423098 566186 423334
rect 566422 423098 590202 423334
rect 590438 423098 590620 423334
rect -6696 423076 590620 423098
rect -6696 423074 -6096 423076
rect 26004 423074 26604 423076
rect 62004 423074 62604 423076
rect 98004 423074 98604 423076
rect 134004 423074 134604 423076
rect 170004 423074 170604 423076
rect 206004 423074 206604 423076
rect 242004 423074 242604 423076
rect 278004 423074 278604 423076
rect 314004 423074 314604 423076
rect 350004 423074 350604 423076
rect 386004 423074 386604 423076
rect 422004 423074 422604 423076
rect 458004 423074 458604 423076
rect 494004 423074 494604 423076
rect 530004 423074 530604 423076
rect 566004 423074 566604 423076
rect 590020 423074 590620 423076
rect -4816 420076 -4216 420078
rect 22404 420076 23004 420078
rect 58404 420076 59004 420078
rect 94404 420076 95004 420078
rect 130404 420076 131004 420078
rect 166404 420076 167004 420078
rect 202404 420076 203004 420078
rect 238404 420076 239004 420078
rect 274404 420076 275004 420078
rect 310404 420076 311004 420078
rect 346404 420076 347004 420078
rect 382404 420076 383004 420078
rect 418404 420076 419004 420078
rect 454404 420076 455004 420078
rect 490404 420076 491004 420078
rect 526404 420076 527004 420078
rect 562404 420076 563004 420078
rect 588140 420076 588740 420078
rect -4816 420054 588740 420076
rect -4816 419818 -4634 420054
rect -4398 419818 22586 420054
rect 22822 419818 58586 420054
rect 58822 419818 94586 420054
rect 94822 419818 130586 420054
rect 130822 419818 166586 420054
rect 166822 419818 202586 420054
rect 202822 419818 238586 420054
rect 238822 419818 274586 420054
rect 274822 419818 310586 420054
rect 310822 419818 346586 420054
rect 346822 419818 382586 420054
rect 382822 419818 418586 420054
rect 418822 419818 454586 420054
rect 454822 419818 490586 420054
rect 490822 419818 526586 420054
rect 526822 419818 562586 420054
rect 562822 419818 588322 420054
rect 588558 419818 588740 420054
rect -4816 419734 588740 419818
rect -4816 419498 -4634 419734
rect -4398 419498 22586 419734
rect 22822 419498 58586 419734
rect 58822 419498 94586 419734
rect 94822 419498 130586 419734
rect 130822 419498 166586 419734
rect 166822 419498 202586 419734
rect 202822 419498 238586 419734
rect 238822 419498 274586 419734
rect 274822 419498 310586 419734
rect 310822 419498 346586 419734
rect 346822 419498 382586 419734
rect 382822 419498 418586 419734
rect 418822 419498 454586 419734
rect 454822 419498 490586 419734
rect 490822 419498 526586 419734
rect 526822 419498 562586 419734
rect 562822 419498 588322 419734
rect 588558 419498 588740 419734
rect -4816 419476 588740 419498
rect -4816 419474 -4216 419476
rect 22404 419474 23004 419476
rect 58404 419474 59004 419476
rect 94404 419474 95004 419476
rect 130404 419474 131004 419476
rect 166404 419474 167004 419476
rect 202404 419474 203004 419476
rect 238404 419474 239004 419476
rect 274404 419474 275004 419476
rect 310404 419474 311004 419476
rect 346404 419474 347004 419476
rect 382404 419474 383004 419476
rect 418404 419474 419004 419476
rect 454404 419474 455004 419476
rect 490404 419474 491004 419476
rect 526404 419474 527004 419476
rect 562404 419474 563004 419476
rect 588140 419474 588740 419476
rect -2936 416476 -2336 416478
rect 18804 416476 19404 416478
rect 54804 416476 55404 416478
rect 90804 416476 91404 416478
rect 126804 416476 127404 416478
rect 162804 416476 163404 416478
rect 198804 416476 199404 416478
rect 234804 416476 235404 416478
rect 270804 416476 271404 416478
rect 306804 416476 307404 416478
rect 342804 416476 343404 416478
rect 378804 416476 379404 416478
rect 414804 416476 415404 416478
rect 450804 416476 451404 416478
rect 486804 416476 487404 416478
rect 522804 416476 523404 416478
rect 558804 416476 559404 416478
rect 586260 416476 586860 416478
rect -2936 416454 586860 416476
rect -2936 416218 -2754 416454
rect -2518 416218 18986 416454
rect 19222 416218 54986 416454
rect 55222 416218 90986 416454
rect 91222 416218 126986 416454
rect 127222 416218 162986 416454
rect 163222 416218 198986 416454
rect 199222 416218 234986 416454
rect 235222 416218 270986 416454
rect 271222 416218 306986 416454
rect 307222 416218 342986 416454
rect 343222 416218 378986 416454
rect 379222 416218 414986 416454
rect 415222 416218 450986 416454
rect 451222 416218 486986 416454
rect 487222 416218 522986 416454
rect 523222 416218 558986 416454
rect 559222 416218 586442 416454
rect 586678 416218 586860 416454
rect -2936 416134 586860 416218
rect -2936 415898 -2754 416134
rect -2518 415898 18986 416134
rect 19222 415898 54986 416134
rect 55222 415898 90986 416134
rect 91222 415898 126986 416134
rect 127222 415898 162986 416134
rect 163222 415898 198986 416134
rect 199222 415898 234986 416134
rect 235222 415898 270986 416134
rect 271222 415898 306986 416134
rect 307222 415898 342986 416134
rect 343222 415898 378986 416134
rect 379222 415898 414986 416134
rect 415222 415898 450986 416134
rect 451222 415898 486986 416134
rect 487222 415898 522986 416134
rect 523222 415898 558986 416134
rect 559222 415898 586442 416134
rect 586678 415898 586860 416134
rect -2936 415876 586860 415898
rect -2936 415874 -2336 415876
rect 18804 415874 19404 415876
rect 54804 415874 55404 415876
rect 90804 415874 91404 415876
rect 126804 415874 127404 415876
rect 162804 415874 163404 415876
rect 198804 415874 199404 415876
rect 234804 415874 235404 415876
rect 270804 415874 271404 415876
rect 306804 415874 307404 415876
rect 342804 415874 343404 415876
rect 378804 415874 379404 415876
rect 414804 415874 415404 415876
rect 450804 415874 451404 415876
rect 486804 415874 487404 415876
rect 522804 415874 523404 415876
rect 558804 415874 559404 415876
rect 586260 415874 586860 415876
rect -7636 409276 -7036 409278
rect 11604 409276 12204 409278
rect 47604 409276 48204 409278
rect 83604 409276 84204 409278
rect 119604 409276 120204 409278
rect 155604 409276 156204 409278
rect 191604 409276 192204 409278
rect 227604 409276 228204 409278
rect 263604 409276 264204 409278
rect 299604 409276 300204 409278
rect 335604 409276 336204 409278
rect 371604 409276 372204 409278
rect 407604 409276 408204 409278
rect 443604 409276 444204 409278
rect 479604 409276 480204 409278
rect 515604 409276 516204 409278
rect 551604 409276 552204 409278
rect 590960 409276 591560 409278
rect -8576 409254 592500 409276
rect -8576 409018 -7454 409254
rect -7218 409018 11786 409254
rect 12022 409018 47786 409254
rect 48022 409018 83786 409254
rect 84022 409018 119786 409254
rect 120022 409018 155786 409254
rect 156022 409018 191786 409254
rect 192022 409018 227786 409254
rect 228022 409018 263786 409254
rect 264022 409018 299786 409254
rect 300022 409018 335786 409254
rect 336022 409018 371786 409254
rect 372022 409018 407786 409254
rect 408022 409018 443786 409254
rect 444022 409018 479786 409254
rect 480022 409018 515786 409254
rect 516022 409018 551786 409254
rect 552022 409018 591142 409254
rect 591378 409018 592500 409254
rect -8576 408934 592500 409018
rect -8576 408698 -7454 408934
rect -7218 408698 11786 408934
rect 12022 408698 47786 408934
rect 48022 408698 83786 408934
rect 84022 408698 119786 408934
rect 120022 408698 155786 408934
rect 156022 408698 191786 408934
rect 192022 408698 227786 408934
rect 228022 408698 263786 408934
rect 264022 408698 299786 408934
rect 300022 408698 335786 408934
rect 336022 408698 371786 408934
rect 372022 408698 407786 408934
rect 408022 408698 443786 408934
rect 444022 408698 479786 408934
rect 480022 408698 515786 408934
rect 516022 408698 551786 408934
rect 552022 408698 591142 408934
rect 591378 408698 592500 408934
rect -8576 408676 592500 408698
rect -7636 408674 -7036 408676
rect 11604 408674 12204 408676
rect 47604 408674 48204 408676
rect 83604 408674 84204 408676
rect 119604 408674 120204 408676
rect 155604 408674 156204 408676
rect 191604 408674 192204 408676
rect 227604 408674 228204 408676
rect 263604 408674 264204 408676
rect 299604 408674 300204 408676
rect 335604 408674 336204 408676
rect 371604 408674 372204 408676
rect 407604 408674 408204 408676
rect 443604 408674 444204 408676
rect 479604 408674 480204 408676
rect 515604 408674 516204 408676
rect 551604 408674 552204 408676
rect 590960 408674 591560 408676
rect -5756 405676 -5156 405678
rect 8004 405676 8604 405678
rect 44004 405676 44604 405678
rect 80004 405676 80604 405678
rect 116004 405676 116604 405678
rect 152004 405676 152604 405678
rect 188004 405676 188604 405678
rect 224004 405676 224604 405678
rect 260004 405676 260604 405678
rect 296004 405676 296604 405678
rect 332004 405676 332604 405678
rect 368004 405676 368604 405678
rect 404004 405676 404604 405678
rect 440004 405676 440604 405678
rect 476004 405676 476604 405678
rect 512004 405676 512604 405678
rect 548004 405676 548604 405678
rect 589080 405676 589680 405678
rect -6696 405654 590620 405676
rect -6696 405418 -5574 405654
rect -5338 405418 8186 405654
rect 8422 405418 44186 405654
rect 44422 405418 80186 405654
rect 80422 405418 116186 405654
rect 116422 405418 152186 405654
rect 152422 405418 188186 405654
rect 188422 405418 224186 405654
rect 224422 405418 260186 405654
rect 260422 405418 296186 405654
rect 296422 405418 332186 405654
rect 332422 405418 368186 405654
rect 368422 405418 404186 405654
rect 404422 405418 440186 405654
rect 440422 405418 476186 405654
rect 476422 405418 512186 405654
rect 512422 405418 548186 405654
rect 548422 405418 589262 405654
rect 589498 405418 590620 405654
rect -6696 405334 590620 405418
rect -6696 405098 -5574 405334
rect -5338 405098 8186 405334
rect 8422 405098 44186 405334
rect 44422 405098 80186 405334
rect 80422 405098 116186 405334
rect 116422 405098 152186 405334
rect 152422 405098 188186 405334
rect 188422 405098 224186 405334
rect 224422 405098 260186 405334
rect 260422 405098 296186 405334
rect 296422 405098 332186 405334
rect 332422 405098 368186 405334
rect 368422 405098 404186 405334
rect 404422 405098 440186 405334
rect 440422 405098 476186 405334
rect 476422 405098 512186 405334
rect 512422 405098 548186 405334
rect 548422 405098 589262 405334
rect 589498 405098 590620 405334
rect -6696 405076 590620 405098
rect -5756 405074 -5156 405076
rect 8004 405074 8604 405076
rect 44004 405074 44604 405076
rect 80004 405074 80604 405076
rect 116004 405074 116604 405076
rect 152004 405074 152604 405076
rect 188004 405074 188604 405076
rect 224004 405074 224604 405076
rect 260004 405074 260604 405076
rect 296004 405074 296604 405076
rect 332004 405074 332604 405076
rect 368004 405074 368604 405076
rect 404004 405074 404604 405076
rect 440004 405074 440604 405076
rect 476004 405074 476604 405076
rect 512004 405074 512604 405076
rect 548004 405074 548604 405076
rect 589080 405074 589680 405076
rect -3876 402076 -3276 402078
rect 4404 402076 5004 402078
rect 40404 402076 41004 402078
rect 76404 402076 77004 402078
rect 112404 402076 113004 402078
rect 148404 402076 149004 402078
rect 184404 402076 185004 402078
rect 220404 402076 221004 402078
rect 256404 402076 257004 402078
rect 292404 402076 293004 402078
rect 328404 402076 329004 402078
rect 364404 402076 365004 402078
rect 400404 402076 401004 402078
rect 436404 402076 437004 402078
rect 472404 402076 473004 402078
rect 508404 402076 509004 402078
rect 544404 402076 545004 402078
rect 580404 402076 581004 402078
rect 587200 402076 587800 402078
rect -4816 402054 588740 402076
rect -4816 401818 -3694 402054
rect -3458 401818 4586 402054
rect 4822 401818 40586 402054
rect 40822 401818 76586 402054
rect 76822 401818 112586 402054
rect 112822 401818 148586 402054
rect 148822 401818 184586 402054
rect 184822 401818 220586 402054
rect 220822 401818 256586 402054
rect 256822 401818 292586 402054
rect 292822 401818 328586 402054
rect 328822 401818 364586 402054
rect 364822 401818 400586 402054
rect 400822 401818 436586 402054
rect 436822 401818 472586 402054
rect 472822 401818 508586 402054
rect 508822 401818 544586 402054
rect 544822 401818 580586 402054
rect 580822 401818 587382 402054
rect 587618 401818 588740 402054
rect -4816 401734 588740 401818
rect -4816 401498 -3694 401734
rect -3458 401498 4586 401734
rect 4822 401498 40586 401734
rect 40822 401498 76586 401734
rect 76822 401498 112586 401734
rect 112822 401498 148586 401734
rect 148822 401498 184586 401734
rect 184822 401498 220586 401734
rect 220822 401498 256586 401734
rect 256822 401498 292586 401734
rect 292822 401498 328586 401734
rect 328822 401498 364586 401734
rect 364822 401498 400586 401734
rect 400822 401498 436586 401734
rect 436822 401498 472586 401734
rect 472822 401498 508586 401734
rect 508822 401498 544586 401734
rect 544822 401498 580586 401734
rect 580822 401498 587382 401734
rect 587618 401498 588740 401734
rect -4816 401476 588740 401498
rect -3876 401474 -3276 401476
rect 4404 401474 5004 401476
rect 40404 401474 41004 401476
rect 76404 401474 77004 401476
rect 112404 401474 113004 401476
rect 148404 401474 149004 401476
rect 184404 401474 185004 401476
rect 220404 401474 221004 401476
rect 256404 401474 257004 401476
rect 292404 401474 293004 401476
rect 328404 401474 329004 401476
rect 364404 401474 365004 401476
rect 400404 401474 401004 401476
rect 436404 401474 437004 401476
rect 472404 401474 473004 401476
rect 508404 401474 509004 401476
rect 544404 401474 545004 401476
rect 580404 401474 581004 401476
rect 587200 401474 587800 401476
rect -1996 398476 -1396 398478
rect 804 398476 1404 398478
rect 36804 398476 37404 398478
rect 72804 398476 73404 398478
rect 108804 398476 109404 398478
rect 144804 398476 145404 398478
rect 180804 398476 181404 398478
rect 216804 398476 217404 398478
rect 252804 398476 253404 398478
rect 288804 398476 289404 398478
rect 324804 398476 325404 398478
rect 360804 398476 361404 398478
rect 396804 398476 397404 398478
rect 432804 398476 433404 398478
rect 468804 398476 469404 398478
rect 504804 398476 505404 398478
rect 540804 398476 541404 398478
rect 576804 398476 577404 398478
rect 585320 398476 585920 398478
rect -2936 398454 586860 398476
rect -2936 398218 -1814 398454
rect -1578 398218 986 398454
rect 1222 398218 36986 398454
rect 37222 398218 72986 398454
rect 73222 398218 108986 398454
rect 109222 398218 144986 398454
rect 145222 398218 180986 398454
rect 181222 398218 216986 398454
rect 217222 398218 252986 398454
rect 253222 398218 288986 398454
rect 289222 398218 324986 398454
rect 325222 398218 360986 398454
rect 361222 398218 396986 398454
rect 397222 398218 432986 398454
rect 433222 398218 468986 398454
rect 469222 398218 504986 398454
rect 505222 398218 540986 398454
rect 541222 398218 576986 398454
rect 577222 398218 585502 398454
rect 585738 398218 586860 398454
rect -2936 398134 586860 398218
rect -2936 397898 -1814 398134
rect -1578 397898 986 398134
rect 1222 397898 36986 398134
rect 37222 397898 72986 398134
rect 73222 397898 108986 398134
rect 109222 397898 144986 398134
rect 145222 397898 180986 398134
rect 181222 397898 216986 398134
rect 217222 397898 252986 398134
rect 253222 397898 288986 398134
rect 289222 397898 324986 398134
rect 325222 397898 360986 398134
rect 361222 397898 396986 398134
rect 397222 397898 432986 398134
rect 433222 397898 468986 398134
rect 469222 397898 504986 398134
rect 505222 397898 540986 398134
rect 541222 397898 576986 398134
rect 577222 397898 585502 398134
rect 585738 397898 586860 398134
rect -2936 397876 586860 397898
rect -1996 397874 -1396 397876
rect 804 397874 1404 397876
rect 36804 397874 37404 397876
rect 72804 397874 73404 397876
rect 108804 397874 109404 397876
rect 144804 397874 145404 397876
rect 180804 397874 181404 397876
rect 216804 397874 217404 397876
rect 252804 397874 253404 397876
rect 288804 397874 289404 397876
rect 324804 397874 325404 397876
rect 360804 397874 361404 397876
rect 396804 397874 397404 397876
rect 432804 397874 433404 397876
rect 468804 397874 469404 397876
rect 504804 397874 505404 397876
rect 540804 397874 541404 397876
rect 576804 397874 577404 397876
rect 585320 397874 585920 397876
rect -8576 391276 -7976 391278
rect 29604 391276 30204 391278
rect 65604 391276 66204 391278
rect 101604 391276 102204 391278
rect 137604 391276 138204 391278
rect 173604 391276 174204 391278
rect 209604 391276 210204 391278
rect 245604 391276 246204 391278
rect 281604 391276 282204 391278
rect 317604 391276 318204 391278
rect 353604 391276 354204 391278
rect 389604 391276 390204 391278
rect 425604 391276 426204 391278
rect 461604 391276 462204 391278
rect 497604 391276 498204 391278
rect 533604 391276 534204 391278
rect 569604 391276 570204 391278
rect 591900 391276 592500 391278
rect -8576 391254 592500 391276
rect -8576 391018 -8394 391254
rect -8158 391018 29786 391254
rect 30022 391018 65786 391254
rect 66022 391018 101786 391254
rect 102022 391018 137786 391254
rect 138022 391018 173786 391254
rect 174022 391018 209786 391254
rect 210022 391018 245786 391254
rect 246022 391018 281786 391254
rect 282022 391018 317786 391254
rect 318022 391018 353786 391254
rect 354022 391018 389786 391254
rect 390022 391018 425786 391254
rect 426022 391018 461786 391254
rect 462022 391018 497786 391254
rect 498022 391018 533786 391254
rect 534022 391018 569786 391254
rect 570022 391018 592082 391254
rect 592318 391018 592500 391254
rect -8576 390934 592500 391018
rect -8576 390698 -8394 390934
rect -8158 390698 29786 390934
rect 30022 390698 65786 390934
rect 66022 390698 101786 390934
rect 102022 390698 137786 390934
rect 138022 390698 173786 390934
rect 174022 390698 209786 390934
rect 210022 390698 245786 390934
rect 246022 390698 281786 390934
rect 282022 390698 317786 390934
rect 318022 390698 353786 390934
rect 354022 390698 389786 390934
rect 390022 390698 425786 390934
rect 426022 390698 461786 390934
rect 462022 390698 497786 390934
rect 498022 390698 533786 390934
rect 534022 390698 569786 390934
rect 570022 390698 592082 390934
rect 592318 390698 592500 390934
rect -8576 390676 592500 390698
rect -8576 390674 -7976 390676
rect 29604 390674 30204 390676
rect 65604 390674 66204 390676
rect 101604 390674 102204 390676
rect 137604 390674 138204 390676
rect 173604 390674 174204 390676
rect 209604 390674 210204 390676
rect 245604 390674 246204 390676
rect 281604 390674 282204 390676
rect 317604 390674 318204 390676
rect 353604 390674 354204 390676
rect 389604 390674 390204 390676
rect 425604 390674 426204 390676
rect 461604 390674 462204 390676
rect 497604 390674 498204 390676
rect 533604 390674 534204 390676
rect 569604 390674 570204 390676
rect 591900 390674 592500 390676
rect -6696 387676 -6096 387678
rect 26004 387676 26604 387678
rect 62004 387676 62604 387678
rect 98004 387676 98604 387678
rect 134004 387676 134604 387678
rect 170004 387676 170604 387678
rect 206004 387676 206604 387678
rect 242004 387676 242604 387678
rect 278004 387676 278604 387678
rect 314004 387676 314604 387678
rect 350004 387676 350604 387678
rect 386004 387676 386604 387678
rect 422004 387676 422604 387678
rect 458004 387676 458604 387678
rect 494004 387676 494604 387678
rect 530004 387676 530604 387678
rect 566004 387676 566604 387678
rect 590020 387676 590620 387678
rect -6696 387654 590620 387676
rect -6696 387418 -6514 387654
rect -6278 387418 26186 387654
rect 26422 387418 62186 387654
rect 62422 387418 98186 387654
rect 98422 387418 134186 387654
rect 134422 387418 170186 387654
rect 170422 387418 206186 387654
rect 206422 387418 242186 387654
rect 242422 387418 278186 387654
rect 278422 387418 314186 387654
rect 314422 387418 350186 387654
rect 350422 387418 386186 387654
rect 386422 387418 422186 387654
rect 422422 387418 458186 387654
rect 458422 387418 494186 387654
rect 494422 387418 530186 387654
rect 530422 387418 566186 387654
rect 566422 387418 590202 387654
rect 590438 387418 590620 387654
rect -6696 387334 590620 387418
rect -6696 387098 -6514 387334
rect -6278 387098 26186 387334
rect 26422 387098 62186 387334
rect 62422 387098 98186 387334
rect 98422 387098 134186 387334
rect 134422 387098 170186 387334
rect 170422 387098 206186 387334
rect 206422 387098 242186 387334
rect 242422 387098 278186 387334
rect 278422 387098 314186 387334
rect 314422 387098 350186 387334
rect 350422 387098 386186 387334
rect 386422 387098 422186 387334
rect 422422 387098 458186 387334
rect 458422 387098 494186 387334
rect 494422 387098 530186 387334
rect 530422 387098 566186 387334
rect 566422 387098 590202 387334
rect 590438 387098 590620 387334
rect -6696 387076 590620 387098
rect -6696 387074 -6096 387076
rect 26004 387074 26604 387076
rect 62004 387074 62604 387076
rect 98004 387074 98604 387076
rect 134004 387074 134604 387076
rect 170004 387074 170604 387076
rect 206004 387074 206604 387076
rect 242004 387074 242604 387076
rect 278004 387074 278604 387076
rect 314004 387074 314604 387076
rect 350004 387074 350604 387076
rect 386004 387074 386604 387076
rect 422004 387074 422604 387076
rect 458004 387074 458604 387076
rect 494004 387074 494604 387076
rect 530004 387074 530604 387076
rect 566004 387074 566604 387076
rect 590020 387074 590620 387076
rect -4816 384076 -4216 384078
rect 22404 384076 23004 384078
rect 58404 384076 59004 384078
rect 94404 384076 95004 384078
rect 130404 384076 131004 384078
rect 166404 384076 167004 384078
rect 202404 384076 203004 384078
rect 238404 384076 239004 384078
rect 274404 384076 275004 384078
rect 310404 384076 311004 384078
rect 346404 384076 347004 384078
rect 382404 384076 383004 384078
rect 418404 384076 419004 384078
rect 454404 384076 455004 384078
rect 490404 384076 491004 384078
rect 526404 384076 527004 384078
rect 562404 384076 563004 384078
rect 588140 384076 588740 384078
rect -4816 384054 588740 384076
rect -4816 383818 -4634 384054
rect -4398 383818 22586 384054
rect 22822 383818 58586 384054
rect 58822 383818 94586 384054
rect 94822 383818 130586 384054
rect 130822 383818 166586 384054
rect 166822 383818 202586 384054
rect 202822 383818 238586 384054
rect 238822 383818 274586 384054
rect 274822 383818 310586 384054
rect 310822 383818 346586 384054
rect 346822 383818 382586 384054
rect 382822 383818 418586 384054
rect 418822 383818 454586 384054
rect 454822 383818 490586 384054
rect 490822 383818 526586 384054
rect 526822 383818 562586 384054
rect 562822 383818 588322 384054
rect 588558 383818 588740 384054
rect -4816 383734 588740 383818
rect -4816 383498 -4634 383734
rect -4398 383498 22586 383734
rect 22822 383498 58586 383734
rect 58822 383498 94586 383734
rect 94822 383498 130586 383734
rect 130822 383498 166586 383734
rect 166822 383498 202586 383734
rect 202822 383498 238586 383734
rect 238822 383498 274586 383734
rect 274822 383498 310586 383734
rect 310822 383498 346586 383734
rect 346822 383498 382586 383734
rect 382822 383498 418586 383734
rect 418822 383498 454586 383734
rect 454822 383498 490586 383734
rect 490822 383498 526586 383734
rect 526822 383498 562586 383734
rect 562822 383498 588322 383734
rect 588558 383498 588740 383734
rect -4816 383476 588740 383498
rect -4816 383474 -4216 383476
rect 22404 383474 23004 383476
rect 58404 383474 59004 383476
rect 94404 383474 95004 383476
rect 130404 383474 131004 383476
rect 166404 383474 167004 383476
rect 202404 383474 203004 383476
rect 238404 383474 239004 383476
rect 274404 383474 275004 383476
rect 310404 383474 311004 383476
rect 346404 383474 347004 383476
rect 382404 383474 383004 383476
rect 418404 383474 419004 383476
rect 454404 383474 455004 383476
rect 490404 383474 491004 383476
rect 526404 383474 527004 383476
rect 562404 383474 563004 383476
rect 588140 383474 588740 383476
rect -2936 380476 -2336 380478
rect 18804 380476 19404 380478
rect 54804 380476 55404 380478
rect 90804 380476 91404 380478
rect 126804 380476 127404 380478
rect 162804 380476 163404 380478
rect 198804 380476 199404 380478
rect 234804 380476 235404 380478
rect 270804 380476 271404 380478
rect 306804 380476 307404 380478
rect 342804 380476 343404 380478
rect 378804 380476 379404 380478
rect 414804 380476 415404 380478
rect 450804 380476 451404 380478
rect 486804 380476 487404 380478
rect 522804 380476 523404 380478
rect 558804 380476 559404 380478
rect 586260 380476 586860 380478
rect -2936 380454 586860 380476
rect -2936 380218 -2754 380454
rect -2518 380218 18986 380454
rect 19222 380218 54986 380454
rect 55222 380218 90986 380454
rect 91222 380218 126986 380454
rect 127222 380218 162986 380454
rect 163222 380218 198986 380454
rect 199222 380218 234986 380454
rect 235222 380218 270986 380454
rect 271222 380218 306986 380454
rect 307222 380218 342986 380454
rect 343222 380218 378986 380454
rect 379222 380218 414986 380454
rect 415222 380218 450986 380454
rect 451222 380218 486986 380454
rect 487222 380218 522986 380454
rect 523222 380218 558986 380454
rect 559222 380218 586442 380454
rect 586678 380218 586860 380454
rect -2936 380134 586860 380218
rect -2936 379898 -2754 380134
rect -2518 379898 18986 380134
rect 19222 379898 54986 380134
rect 55222 379898 90986 380134
rect 91222 379898 126986 380134
rect 127222 379898 162986 380134
rect 163222 379898 198986 380134
rect 199222 379898 234986 380134
rect 235222 379898 270986 380134
rect 271222 379898 306986 380134
rect 307222 379898 342986 380134
rect 343222 379898 378986 380134
rect 379222 379898 414986 380134
rect 415222 379898 450986 380134
rect 451222 379898 486986 380134
rect 487222 379898 522986 380134
rect 523222 379898 558986 380134
rect 559222 379898 586442 380134
rect 586678 379898 586860 380134
rect -2936 379876 586860 379898
rect -2936 379874 -2336 379876
rect 18804 379874 19404 379876
rect 54804 379874 55404 379876
rect 90804 379874 91404 379876
rect 126804 379874 127404 379876
rect 162804 379874 163404 379876
rect 198804 379874 199404 379876
rect 234804 379874 235404 379876
rect 270804 379874 271404 379876
rect 306804 379874 307404 379876
rect 342804 379874 343404 379876
rect 378804 379874 379404 379876
rect 414804 379874 415404 379876
rect 450804 379874 451404 379876
rect 486804 379874 487404 379876
rect 522804 379874 523404 379876
rect 558804 379874 559404 379876
rect 586260 379874 586860 379876
rect -7636 373276 -7036 373278
rect 11604 373276 12204 373278
rect 47604 373276 48204 373278
rect 83604 373276 84204 373278
rect 119604 373276 120204 373278
rect 155604 373276 156204 373278
rect 191604 373276 192204 373278
rect 227604 373276 228204 373278
rect 263604 373276 264204 373278
rect 299604 373276 300204 373278
rect 335604 373276 336204 373278
rect 371604 373276 372204 373278
rect 407604 373276 408204 373278
rect 443604 373276 444204 373278
rect 479604 373276 480204 373278
rect 515604 373276 516204 373278
rect 551604 373276 552204 373278
rect 590960 373276 591560 373278
rect -8576 373254 592500 373276
rect -8576 373018 -7454 373254
rect -7218 373018 11786 373254
rect 12022 373018 47786 373254
rect 48022 373018 83786 373254
rect 84022 373018 119786 373254
rect 120022 373018 155786 373254
rect 156022 373018 191786 373254
rect 192022 373018 227786 373254
rect 228022 373018 263786 373254
rect 264022 373018 299786 373254
rect 300022 373018 335786 373254
rect 336022 373018 371786 373254
rect 372022 373018 407786 373254
rect 408022 373018 443786 373254
rect 444022 373018 479786 373254
rect 480022 373018 515786 373254
rect 516022 373018 551786 373254
rect 552022 373018 591142 373254
rect 591378 373018 592500 373254
rect -8576 372934 592500 373018
rect -8576 372698 -7454 372934
rect -7218 372698 11786 372934
rect 12022 372698 47786 372934
rect 48022 372698 83786 372934
rect 84022 372698 119786 372934
rect 120022 372698 155786 372934
rect 156022 372698 191786 372934
rect 192022 372698 227786 372934
rect 228022 372698 263786 372934
rect 264022 372698 299786 372934
rect 300022 372698 335786 372934
rect 336022 372698 371786 372934
rect 372022 372698 407786 372934
rect 408022 372698 443786 372934
rect 444022 372698 479786 372934
rect 480022 372698 515786 372934
rect 516022 372698 551786 372934
rect 552022 372698 591142 372934
rect 591378 372698 592500 372934
rect -8576 372676 592500 372698
rect -7636 372674 -7036 372676
rect 11604 372674 12204 372676
rect 47604 372674 48204 372676
rect 83604 372674 84204 372676
rect 119604 372674 120204 372676
rect 155604 372674 156204 372676
rect 191604 372674 192204 372676
rect 227604 372674 228204 372676
rect 263604 372674 264204 372676
rect 299604 372674 300204 372676
rect 335604 372674 336204 372676
rect 371604 372674 372204 372676
rect 407604 372674 408204 372676
rect 443604 372674 444204 372676
rect 479604 372674 480204 372676
rect 515604 372674 516204 372676
rect 551604 372674 552204 372676
rect 590960 372674 591560 372676
rect -5756 369676 -5156 369678
rect 8004 369676 8604 369678
rect 44004 369676 44604 369678
rect 80004 369676 80604 369678
rect 116004 369676 116604 369678
rect 152004 369676 152604 369678
rect 188004 369676 188604 369678
rect 224004 369676 224604 369678
rect 260004 369676 260604 369678
rect 296004 369676 296604 369678
rect 332004 369676 332604 369678
rect 368004 369676 368604 369678
rect 404004 369676 404604 369678
rect 440004 369676 440604 369678
rect 476004 369676 476604 369678
rect 512004 369676 512604 369678
rect 548004 369676 548604 369678
rect 589080 369676 589680 369678
rect -6696 369654 590620 369676
rect -6696 369418 -5574 369654
rect -5338 369418 8186 369654
rect 8422 369418 44186 369654
rect 44422 369418 80186 369654
rect 80422 369418 116186 369654
rect 116422 369418 152186 369654
rect 152422 369418 188186 369654
rect 188422 369418 224186 369654
rect 224422 369418 260186 369654
rect 260422 369418 296186 369654
rect 296422 369418 332186 369654
rect 332422 369418 368186 369654
rect 368422 369418 404186 369654
rect 404422 369418 440186 369654
rect 440422 369418 476186 369654
rect 476422 369418 512186 369654
rect 512422 369418 548186 369654
rect 548422 369418 589262 369654
rect 589498 369418 590620 369654
rect -6696 369334 590620 369418
rect -6696 369098 -5574 369334
rect -5338 369098 8186 369334
rect 8422 369098 44186 369334
rect 44422 369098 80186 369334
rect 80422 369098 116186 369334
rect 116422 369098 152186 369334
rect 152422 369098 188186 369334
rect 188422 369098 224186 369334
rect 224422 369098 260186 369334
rect 260422 369098 296186 369334
rect 296422 369098 332186 369334
rect 332422 369098 368186 369334
rect 368422 369098 404186 369334
rect 404422 369098 440186 369334
rect 440422 369098 476186 369334
rect 476422 369098 512186 369334
rect 512422 369098 548186 369334
rect 548422 369098 589262 369334
rect 589498 369098 590620 369334
rect -6696 369076 590620 369098
rect -5756 369074 -5156 369076
rect 8004 369074 8604 369076
rect 44004 369074 44604 369076
rect 80004 369074 80604 369076
rect 116004 369074 116604 369076
rect 152004 369074 152604 369076
rect 188004 369074 188604 369076
rect 224004 369074 224604 369076
rect 260004 369074 260604 369076
rect 296004 369074 296604 369076
rect 332004 369074 332604 369076
rect 368004 369074 368604 369076
rect 404004 369074 404604 369076
rect 440004 369074 440604 369076
rect 476004 369074 476604 369076
rect 512004 369074 512604 369076
rect 548004 369074 548604 369076
rect 589080 369074 589680 369076
rect -3876 366076 -3276 366078
rect 4404 366076 5004 366078
rect 40404 366076 41004 366078
rect 76404 366076 77004 366078
rect 112404 366076 113004 366078
rect 148404 366076 149004 366078
rect 184404 366076 185004 366078
rect 220404 366076 221004 366078
rect 256404 366076 257004 366078
rect 292404 366076 293004 366078
rect 328404 366076 329004 366078
rect 364404 366076 365004 366078
rect 400404 366076 401004 366078
rect 436404 366076 437004 366078
rect 472404 366076 473004 366078
rect 508404 366076 509004 366078
rect 544404 366076 545004 366078
rect 580404 366076 581004 366078
rect 587200 366076 587800 366078
rect -4816 366054 588740 366076
rect -4816 365818 -3694 366054
rect -3458 365818 4586 366054
rect 4822 365818 40586 366054
rect 40822 365818 76586 366054
rect 76822 365818 112586 366054
rect 112822 365818 148586 366054
rect 148822 365818 184586 366054
rect 184822 365818 220586 366054
rect 220822 365818 256586 366054
rect 256822 365818 292586 366054
rect 292822 365818 328586 366054
rect 328822 365818 364586 366054
rect 364822 365818 400586 366054
rect 400822 365818 436586 366054
rect 436822 365818 472586 366054
rect 472822 365818 508586 366054
rect 508822 365818 544586 366054
rect 544822 365818 580586 366054
rect 580822 365818 587382 366054
rect 587618 365818 588740 366054
rect -4816 365734 588740 365818
rect -4816 365498 -3694 365734
rect -3458 365498 4586 365734
rect 4822 365498 40586 365734
rect 40822 365498 76586 365734
rect 76822 365498 112586 365734
rect 112822 365498 148586 365734
rect 148822 365498 184586 365734
rect 184822 365498 220586 365734
rect 220822 365498 256586 365734
rect 256822 365498 292586 365734
rect 292822 365498 328586 365734
rect 328822 365498 364586 365734
rect 364822 365498 400586 365734
rect 400822 365498 436586 365734
rect 436822 365498 472586 365734
rect 472822 365498 508586 365734
rect 508822 365498 544586 365734
rect 544822 365498 580586 365734
rect 580822 365498 587382 365734
rect 587618 365498 588740 365734
rect -4816 365476 588740 365498
rect -3876 365474 -3276 365476
rect 4404 365474 5004 365476
rect 40404 365474 41004 365476
rect 76404 365474 77004 365476
rect 112404 365474 113004 365476
rect 148404 365474 149004 365476
rect 184404 365474 185004 365476
rect 220404 365474 221004 365476
rect 256404 365474 257004 365476
rect 292404 365474 293004 365476
rect 328404 365474 329004 365476
rect 364404 365474 365004 365476
rect 400404 365474 401004 365476
rect 436404 365474 437004 365476
rect 472404 365474 473004 365476
rect 508404 365474 509004 365476
rect 544404 365474 545004 365476
rect 580404 365474 581004 365476
rect 587200 365474 587800 365476
rect -1996 362476 -1396 362478
rect 804 362476 1404 362478
rect 36804 362476 37404 362478
rect 72804 362476 73404 362478
rect 108804 362476 109404 362478
rect 144804 362476 145404 362478
rect 180804 362476 181404 362478
rect 216804 362476 217404 362478
rect 252804 362476 253404 362478
rect 288804 362476 289404 362478
rect 324804 362476 325404 362478
rect 360804 362476 361404 362478
rect 396804 362476 397404 362478
rect 432804 362476 433404 362478
rect 468804 362476 469404 362478
rect 504804 362476 505404 362478
rect 540804 362476 541404 362478
rect 576804 362476 577404 362478
rect 585320 362476 585920 362478
rect -2936 362454 586860 362476
rect -2936 362218 -1814 362454
rect -1578 362218 986 362454
rect 1222 362218 36986 362454
rect 37222 362218 72986 362454
rect 73222 362218 108986 362454
rect 109222 362218 144986 362454
rect 145222 362218 180986 362454
rect 181222 362218 216986 362454
rect 217222 362218 252986 362454
rect 253222 362218 288986 362454
rect 289222 362218 324986 362454
rect 325222 362218 360986 362454
rect 361222 362218 396986 362454
rect 397222 362218 432986 362454
rect 433222 362218 468986 362454
rect 469222 362218 504986 362454
rect 505222 362218 540986 362454
rect 541222 362218 576986 362454
rect 577222 362218 585502 362454
rect 585738 362218 586860 362454
rect -2936 362134 586860 362218
rect -2936 361898 -1814 362134
rect -1578 361898 986 362134
rect 1222 361898 36986 362134
rect 37222 361898 72986 362134
rect 73222 361898 108986 362134
rect 109222 361898 144986 362134
rect 145222 361898 180986 362134
rect 181222 361898 216986 362134
rect 217222 361898 252986 362134
rect 253222 361898 288986 362134
rect 289222 361898 324986 362134
rect 325222 361898 360986 362134
rect 361222 361898 396986 362134
rect 397222 361898 432986 362134
rect 433222 361898 468986 362134
rect 469222 361898 504986 362134
rect 505222 361898 540986 362134
rect 541222 361898 576986 362134
rect 577222 361898 585502 362134
rect 585738 361898 586860 362134
rect -2936 361876 586860 361898
rect -1996 361874 -1396 361876
rect 804 361874 1404 361876
rect 36804 361874 37404 361876
rect 72804 361874 73404 361876
rect 108804 361874 109404 361876
rect 144804 361874 145404 361876
rect 180804 361874 181404 361876
rect 216804 361874 217404 361876
rect 252804 361874 253404 361876
rect 288804 361874 289404 361876
rect 324804 361874 325404 361876
rect 360804 361874 361404 361876
rect 396804 361874 397404 361876
rect 432804 361874 433404 361876
rect 468804 361874 469404 361876
rect 504804 361874 505404 361876
rect 540804 361874 541404 361876
rect 576804 361874 577404 361876
rect 585320 361874 585920 361876
rect -8576 355276 -7976 355278
rect 29604 355276 30204 355278
rect 65604 355276 66204 355278
rect 101604 355276 102204 355278
rect 137604 355276 138204 355278
rect 173604 355276 174204 355278
rect 209604 355276 210204 355278
rect 245604 355276 246204 355278
rect 281604 355276 282204 355278
rect 317604 355276 318204 355278
rect 353604 355276 354204 355278
rect 389604 355276 390204 355278
rect 425604 355276 426204 355278
rect 461604 355276 462204 355278
rect 497604 355276 498204 355278
rect 533604 355276 534204 355278
rect 569604 355276 570204 355278
rect 591900 355276 592500 355278
rect -8576 355254 592500 355276
rect -8576 355018 -8394 355254
rect -8158 355018 29786 355254
rect 30022 355018 65786 355254
rect 66022 355018 101786 355254
rect 102022 355018 137786 355254
rect 138022 355018 173786 355254
rect 174022 355018 209786 355254
rect 210022 355018 245786 355254
rect 246022 355018 281786 355254
rect 282022 355018 317786 355254
rect 318022 355018 353786 355254
rect 354022 355018 389786 355254
rect 390022 355018 425786 355254
rect 426022 355018 461786 355254
rect 462022 355018 497786 355254
rect 498022 355018 533786 355254
rect 534022 355018 569786 355254
rect 570022 355018 592082 355254
rect 592318 355018 592500 355254
rect -8576 354934 592500 355018
rect -8576 354698 -8394 354934
rect -8158 354698 29786 354934
rect 30022 354698 65786 354934
rect 66022 354698 101786 354934
rect 102022 354698 137786 354934
rect 138022 354698 173786 354934
rect 174022 354698 209786 354934
rect 210022 354698 245786 354934
rect 246022 354698 281786 354934
rect 282022 354698 317786 354934
rect 318022 354698 353786 354934
rect 354022 354698 389786 354934
rect 390022 354698 425786 354934
rect 426022 354698 461786 354934
rect 462022 354698 497786 354934
rect 498022 354698 533786 354934
rect 534022 354698 569786 354934
rect 570022 354698 592082 354934
rect 592318 354698 592500 354934
rect -8576 354676 592500 354698
rect -8576 354674 -7976 354676
rect 29604 354674 30204 354676
rect 65604 354674 66204 354676
rect 101604 354674 102204 354676
rect 137604 354674 138204 354676
rect 173604 354674 174204 354676
rect 209604 354674 210204 354676
rect 245604 354674 246204 354676
rect 281604 354674 282204 354676
rect 317604 354674 318204 354676
rect 353604 354674 354204 354676
rect 389604 354674 390204 354676
rect 425604 354674 426204 354676
rect 461604 354674 462204 354676
rect 497604 354674 498204 354676
rect 533604 354674 534204 354676
rect 569604 354674 570204 354676
rect 591900 354674 592500 354676
rect -6696 351676 -6096 351678
rect 26004 351676 26604 351678
rect 62004 351676 62604 351678
rect 98004 351676 98604 351678
rect 134004 351676 134604 351678
rect 170004 351676 170604 351678
rect 206004 351676 206604 351678
rect 242004 351676 242604 351678
rect 278004 351676 278604 351678
rect 314004 351676 314604 351678
rect 350004 351676 350604 351678
rect 386004 351676 386604 351678
rect 422004 351676 422604 351678
rect 458004 351676 458604 351678
rect 494004 351676 494604 351678
rect 530004 351676 530604 351678
rect 566004 351676 566604 351678
rect 590020 351676 590620 351678
rect -6696 351654 590620 351676
rect -6696 351418 -6514 351654
rect -6278 351418 26186 351654
rect 26422 351418 62186 351654
rect 62422 351418 98186 351654
rect 98422 351418 134186 351654
rect 134422 351418 170186 351654
rect 170422 351418 206186 351654
rect 206422 351418 242186 351654
rect 242422 351418 278186 351654
rect 278422 351418 314186 351654
rect 314422 351418 350186 351654
rect 350422 351418 386186 351654
rect 386422 351418 422186 351654
rect 422422 351418 458186 351654
rect 458422 351418 494186 351654
rect 494422 351418 530186 351654
rect 530422 351418 566186 351654
rect 566422 351418 590202 351654
rect 590438 351418 590620 351654
rect -6696 351334 590620 351418
rect -6696 351098 -6514 351334
rect -6278 351098 26186 351334
rect 26422 351098 62186 351334
rect 62422 351098 98186 351334
rect 98422 351098 134186 351334
rect 134422 351098 170186 351334
rect 170422 351098 206186 351334
rect 206422 351098 242186 351334
rect 242422 351098 278186 351334
rect 278422 351098 314186 351334
rect 314422 351098 350186 351334
rect 350422 351098 386186 351334
rect 386422 351098 422186 351334
rect 422422 351098 458186 351334
rect 458422 351098 494186 351334
rect 494422 351098 530186 351334
rect 530422 351098 566186 351334
rect 566422 351098 590202 351334
rect 590438 351098 590620 351334
rect -6696 351076 590620 351098
rect -6696 351074 -6096 351076
rect 26004 351074 26604 351076
rect 62004 351074 62604 351076
rect 98004 351074 98604 351076
rect 134004 351074 134604 351076
rect 170004 351074 170604 351076
rect 206004 351074 206604 351076
rect 242004 351074 242604 351076
rect 278004 351074 278604 351076
rect 314004 351074 314604 351076
rect 350004 351074 350604 351076
rect 386004 351074 386604 351076
rect 422004 351074 422604 351076
rect 458004 351074 458604 351076
rect 494004 351074 494604 351076
rect 530004 351074 530604 351076
rect 566004 351074 566604 351076
rect 590020 351074 590620 351076
rect -4816 348076 -4216 348078
rect 22404 348076 23004 348078
rect 58404 348076 59004 348078
rect 94404 348076 95004 348078
rect 130404 348076 131004 348078
rect 166404 348076 167004 348078
rect 202404 348076 203004 348078
rect 238404 348076 239004 348078
rect 274404 348076 275004 348078
rect 310404 348076 311004 348078
rect 346404 348076 347004 348078
rect 382404 348076 383004 348078
rect 418404 348076 419004 348078
rect 454404 348076 455004 348078
rect 490404 348076 491004 348078
rect 526404 348076 527004 348078
rect 562404 348076 563004 348078
rect 588140 348076 588740 348078
rect -4816 348054 588740 348076
rect -4816 347818 -4634 348054
rect -4398 347818 22586 348054
rect 22822 347818 58586 348054
rect 58822 347818 94586 348054
rect 94822 347818 130586 348054
rect 130822 347818 166586 348054
rect 166822 347818 202586 348054
rect 202822 347818 238586 348054
rect 238822 347818 274586 348054
rect 274822 347818 310586 348054
rect 310822 347818 346586 348054
rect 346822 347818 382586 348054
rect 382822 347818 418586 348054
rect 418822 347818 454586 348054
rect 454822 347818 490586 348054
rect 490822 347818 526586 348054
rect 526822 347818 562586 348054
rect 562822 347818 588322 348054
rect 588558 347818 588740 348054
rect -4816 347734 588740 347818
rect -4816 347498 -4634 347734
rect -4398 347498 22586 347734
rect 22822 347498 58586 347734
rect 58822 347498 94586 347734
rect 94822 347498 130586 347734
rect 130822 347498 166586 347734
rect 166822 347498 202586 347734
rect 202822 347498 238586 347734
rect 238822 347498 274586 347734
rect 274822 347498 310586 347734
rect 310822 347498 346586 347734
rect 346822 347498 382586 347734
rect 382822 347498 418586 347734
rect 418822 347498 454586 347734
rect 454822 347498 490586 347734
rect 490822 347498 526586 347734
rect 526822 347498 562586 347734
rect 562822 347498 588322 347734
rect 588558 347498 588740 347734
rect -4816 347476 588740 347498
rect -4816 347474 -4216 347476
rect 22404 347474 23004 347476
rect 58404 347474 59004 347476
rect 94404 347474 95004 347476
rect 130404 347474 131004 347476
rect 166404 347474 167004 347476
rect 202404 347474 203004 347476
rect 238404 347474 239004 347476
rect 274404 347474 275004 347476
rect 310404 347474 311004 347476
rect 346404 347474 347004 347476
rect 382404 347474 383004 347476
rect 418404 347474 419004 347476
rect 454404 347474 455004 347476
rect 490404 347474 491004 347476
rect 526404 347474 527004 347476
rect 562404 347474 563004 347476
rect 588140 347474 588740 347476
rect -2936 344476 -2336 344478
rect 18804 344476 19404 344478
rect 54804 344476 55404 344478
rect 90804 344476 91404 344478
rect 126804 344476 127404 344478
rect 162804 344476 163404 344478
rect 198804 344476 199404 344478
rect 234804 344476 235404 344478
rect 270804 344476 271404 344478
rect 306804 344476 307404 344478
rect 342804 344476 343404 344478
rect 378804 344476 379404 344478
rect 414804 344476 415404 344478
rect 450804 344476 451404 344478
rect 486804 344476 487404 344478
rect 522804 344476 523404 344478
rect 558804 344476 559404 344478
rect 586260 344476 586860 344478
rect -2936 344454 586860 344476
rect -2936 344218 -2754 344454
rect -2518 344218 18986 344454
rect 19222 344218 54986 344454
rect 55222 344218 90986 344454
rect 91222 344218 126986 344454
rect 127222 344218 162986 344454
rect 163222 344218 198986 344454
rect 199222 344218 234986 344454
rect 235222 344218 270986 344454
rect 271222 344218 306986 344454
rect 307222 344218 342986 344454
rect 343222 344218 378986 344454
rect 379222 344218 414986 344454
rect 415222 344218 450986 344454
rect 451222 344218 486986 344454
rect 487222 344218 522986 344454
rect 523222 344218 558986 344454
rect 559222 344218 586442 344454
rect 586678 344218 586860 344454
rect -2936 344134 586860 344218
rect -2936 343898 -2754 344134
rect -2518 343898 18986 344134
rect 19222 343898 54986 344134
rect 55222 343898 90986 344134
rect 91222 343898 126986 344134
rect 127222 343898 162986 344134
rect 163222 343898 198986 344134
rect 199222 343898 234986 344134
rect 235222 343898 270986 344134
rect 271222 343898 306986 344134
rect 307222 343898 342986 344134
rect 343222 343898 378986 344134
rect 379222 343898 414986 344134
rect 415222 343898 450986 344134
rect 451222 343898 486986 344134
rect 487222 343898 522986 344134
rect 523222 343898 558986 344134
rect 559222 343898 586442 344134
rect 586678 343898 586860 344134
rect -2936 343876 586860 343898
rect -2936 343874 -2336 343876
rect 18804 343874 19404 343876
rect 54804 343874 55404 343876
rect 90804 343874 91404 343876
rect 126804 343874 127404 343876
rect 162804 343874 163404 343876
rect 198804 343874 199404 343876
rect 234804 343874 235404 343876
rect 270804 343874 271404 343876
rect 306804 343874 307404 343876
rect 342804 343874 343404 343876
rect 378804 343874 379404 343876
rect 414804 343874 415404 343876
rect 450804 343874 451404 343876
rect 486804 343874 487404 343876
rect 522804 343874 523404 343876
rect 558804 343874 559404 343876
rect 586260 343874 586860 343876
rect -7636 337276 -7036 337278
rect 11604 337276 12204 337278
rect 47604 337276 48204 337278
rect 83604 337276 84204 337278
rect 119604 337276 120204 337278
rect 155604 337276 156204 337278
rect 191604 337276 192204 337278
rect 227604 337276 228204 337278
rect 263604 337276 264204 337278
rect 299604 337276 300204 337278
rect 335604 337276 336204 337278
rect 371604 337276 372204 337278
rect 407604 337276 408204 337278
rect 443604 337276 444204 337278
rect 479604 337276 480204 337278
rect 515604 337276 516204 337278
rect 551604 337276 552204 337278
rect 590960 337276 591560 337278
rect -8576 337254 592500 337276
rect -8576 337018 -7454 337254
rect -7218 337018 11786 337254
rect 12022 337018 47786 337254
rect 48022 337018 83786 337254
rect 84022 337018 119786 337254
rect 120022 337018 155786 337254
rect 156022 337018 191786 337254
rect 192022 337018 227786 337254
rect 228022 337018 263786 337254
rect 264022 337018 299786 337254
rect 300022 337018 335786 337254
rect 336022 337018 371786 337254
rect 372022 337018 407786 337254
rect 408022 337018 443786 337254
rect 444022 337018 479786 337254
rect 480022 337018 515786 337254
rect 516022 337018 551786 337254
rect 552022 337018 591142 337254
rect 591378 337018 592500 337254
rect -8576 336934 592500 337018
rect -8576 336698 -7454 336934
rect -7218 336698 11786 336934
rect 12022 336698 47786 336934
rect 48022 336698 83786 336934
rect 84022 336698 119786 336934
rect 120022 336698 155786 336934
rect 156022 336698 191786 336934
rect 192022 336698 227786 336934
rect 228022 336698 263786 336934
rect 264022 336698 299786 336934
rect 300022 336698 335786 336934
rect 336022 336698 371786 336934
rect 372022 336698 407786 336934
rect 408022 336698 443786 336934
rect 444022 336698 479786 336934
rect 480022 336698 515786 336934
rect 516022 336698 551786 336934
rect 552022 336698 591142 336934
rect 591378 336698 592500 336934
rect -8576 336676 592500 336698
rect -7636 336674 -7036 336676
rect 11604 336674 12204 336676
rect 47604 336674 48204 336676
rect 83604 336674 84204 336676
rect 119604 336674 120204 336676
rect 155604 336674 156204 336676
rect 191604 336674 192204 336676
rect 227604 336674 228204 336676
rect 263604 336674 264204 336676
rect 299604 336674 300204 336676
rect 335604 336674 336204 336676
rect 371604 336674 372204 336676
rect 407604 336674 408204 336676
rect 443604 336674 444204 336676
rect 479604 336674 480204 336676
rect 515604 336674 516204 336676
rect 551604 336674 552204 336676
rect 590960 336674 591560 336676
rect -5756 333676 -5156 333678
rect 8004 333676 8604 333678
rect 44004 333676 44604 333678
rect 80004 333676 80604 333678
rect 116004 333676 116604 333678
rect 152004 333676 152604 333678
rect 188004 333676 188604 333678
rect 224004 333676 224604 333678
rect 260004 333676 260604 333678
rect 296004 333676 296604 333678
rect 332004 333676 332604 333678
rect 368004 333676 368604 333678
rect 404004 333676 404604 333678
rect 440004 333676 440604 333678
rect 476004 333676 476604 333678
rect 512004 333676 512604 333678
rect 548004 333676 548604 333678
rect 589080 333676 589680 333678
rect -6696 333654 590620 333676
rect -6696 333418 -5574 333654
rect -5338 333418 8186 333654
rect 8422 333418 44186 333654
rect 44422 333418 80186 333654
rect 80422 333418 116186 333654
rect 116422 333418 152186 333654
rect 152422 333418 188186 333654
rect 188422 333418 224186 333654
rect 224422 333418 260186 333654
rect 260422 333418 296186 333654
rect 296422 333418 332186 333654
rect 332422 333418 368186 333654
rect 368422 333418 404186 333654
rect 404422 333418 440186 333654
rect 440422 333418 476186 333654
rect 476422 333418 512186 333654
rect 512422 333418 548186 333654
rect 548422 333418 589262 333654
rect 589498 333418 590620 333654
rect -6696 333334 590620 333418
rect -6696 333098 -5574 333334
rect -5338 333098 8186 333334
rect 8422 333098 44186 333334
rect 44422 333098 80186 333334
rect 80422 333098 116186 333334
rect 116422 333098 152186 333334
rect 152422 333098 188186 333334
rect 188422 333098 224186 333334
rect 224422 333098 260186 333334
rect 260422 333098 296186 333334
rect 296422 333098 332186 333334
rect 332422 333098 368186 333334
rect 368422 333098 404186 333334
rect 404422 333098 440186 333334
rect 440422 333098 476186 333334
rect 476422 333098 512186 333334
rect 512422 333098 548186 333334
rect 548422 333098 589262 333334
rect 589498 333098 590620 333334
rect -6696 333076 590620 333098
rect -5756 333074 -5156 333076
rect 8004 333074 8604 333076
rect 44004 333074 44604 333076
rect 80004 333074 80604 333076
rect 116004 333074 116604 333076
rect 152004 333074 152604 333076
rect 188004 333074 188604 333076
rect 224004 333074 224604 333076
rect 260004 333074 260604 333076
rect 296004 333074 296604 333076
rect 332004 333074 332604 333076
rect 368004 333074 368604 333076
rect 404004 333074 404604 333076
rect 440004 333074 440604 333076
rect 476004 333074 476604 333076
rect 512004 333074 512604 333076
rect 548004 333074 548604 333076
rect 589080 333074 589680 333076
rect -3876 330076 -3276 330078
rect 4404 330076 5004 330078
rect 40404 330076 41004 330078
rect 76404 330076 77004 330078
rect 112404 330076 113004 330078
rect 148404 330076 149004 330078
rect 184404 330076 185004 330078
rect 220404 330076 221004 330078
rect 256404 330076 257004 330078
rect 292404 330076 293004 330078
rect 328404 330076 329004 330078
rect 364404 330076 365004 330078
rect 400404 330076 401004 330078
rect 436404 330076 437004 330078
rect 472404 330076 473004 330078
rect 508404 330076 509004 330078
rect 544404 330076 545004 330078
rect 580404 330076 581004 330078
rect 587200 330076 587800 330078
rect -4816 330054 588740 330076
rect -4816 329818 -3694 330054
rect -3458 329818 4586 330054
rect 4822 329818 40586 330054
rect 40822 329818 76586 330054
rect 76822 329818 112586 330054
rect 112822 329818 148586 330054
rect 148822 329818 184586 330054
rect 184822 329818 220586 330054
rect 220822 329818 256586 330054
rect 256822 329818 292586 330054
rect 292822 329818 328586 330054
rect 328822 329818 364586 330054
rect 364822 329818 400586 330054
rect 400822 329818 436586 330054
rect 436822 329818 472586 330054
rect 472822 329818 508586 330054
rect 508822 329818 544586 330054
rect 544822 329818 580586 330054
rect 580822 329818 587382 330054
rect 587618 329818 588740 330054
rect -4816 329734 588740 329818
rect -4816 329498 -3694 329734
rect -3458 329498 4586 329734
rect 4822 329498 40586 329734
rect 40822 329498 76586 329734
rect 76822 329498 112586 329734
rect 112822 329498 148586 329734
rect 148822 329498 184586 329734
rect 184822 329498 220586 329734
rect 220822 329498 256586 329734
rect 256822 329498 292586 329734
rect 292822 329498 328586 329734
rect 328822 329498 364586 329734
rect 364822 329498 400586 329734
rect 400822 329498 436586 329734
rect 436822 329498 472586 329734
rect 472822 329498 508586 329734
rect 508822 329498 544586 329734
rect 544822 329498 580586 329734
rect 580822 329498 587382 329734
rect 587618 329498 588740 329734
rect -4816 329476 588740 329498
rect -3876 329474 -3276 329476
rect 4404 329474 5004 329476
rect 40404 329474 41004 329476
rect 76404 329474 77004 329476
rect 112404 329474 113004 329476
rect 148404 329474 149004 329476
rect 184404 329474 185004 329476
rect 220404 329474 221004 329476
rect 256404 329474 257004 329476
rect 292404 329474 293004 329476
rect 328404 329474 329004 329476
rect 364404 329474 365004 329476
rect 400404 329474 401004 329476
rect 436404 329474 437004 329476
rect 472404 329474 473004 329476
rect 508404 329474 509004 329476
rect 544404 329474 545004 329476
rect 580404 329474 581004 329476
rect 587200 329474 587800 329476
rect -1996 326476 -1396 326478
rect 804 326476 1404 326478
rect 36804 326476 37404 326478
rect 72804 326476 73404 326478
rect 108804 326476 109404 326478
rect 144804 326476 145404 326478
rect 180804 326476 181404 326478
rect 216804 326476 217404 326478
rect 252804 326476 253404 326478
rect 288804 326476 289404 326478
rect 324804 326476 325404 326478
rect 360804 326476 361404 326478
rect 396804 326476 397404 326478
rect 432804 326476 433404 326478
rect 468804 326476 469404 326478
rect 504804 326476 505404 326478
rect 540804 326476 541404 326478
rect 576804 326476 577404 326478
rect 585320 326476 585920 326478
rect -2936 326454 586860 326476
rect -2936 326218 -1814 326454
rect -1578 326218 986 326454
rect 1222 326218 36986 326454
rect 37222 326218 72986 326454
rect 73222 326218 108986 326454
rect 109222 326218 144986 326454
rect 145222 326218 180986 326454
rect 181222 326218 216986 326454
rect 217222 326218 252986 326454
rect 253222 326218 288986 326454
rect 289222 326218 324986 326454
rect 325222 326218 360986 326454
rect 361222 326218 396986 326454
rect 397222 326218 432986 326454
rect 433222 326218 468986 326454
rect 469222 326218 504986 326454
rect 505222 326218 540986 326454
rect 541222 326218 576986 326454
rect 577222 326218 585502 326454
rect 585738 326218 586860 326454
rect -2936 326134 586860 326218
rect -2936 325898 -1814 326134
rect -1578 325898 986 326134
rect 1222 325898 36986 326134
rect 37222 325898 72986 326134
rect 73222 325898 108986 326134
rect 109222 325898 144986 326134
rect 145222 325898 180986 326134
rect 181222 325898 216986 326134
rect 217222 325898 252986 326134
rect 253222 325898 288986 326134
rect 289222 325898 324986 326134
rect 325222 325898 360986 326134
rect 361222 325898 396986 326134
rect 397222 325898 432986 326134
rect 433222 325898 468986 326134
rect 469222 325898 504986 326134
rect 505222 325898 540986 326134
rect 541222 325898 576986 326134
rect 577222 325898 585502 326134
rect 585738 325898 586860 326134
rect -2936 325876 586860 325898
rect -1996 325874 -1396 325876
rect 804 325874 1404 325876
rect 36804 325874 37404 325876
rect 72804 325874 73404 325876
rect 108804 325874 109404 325876
rect 144804 325874 145404 325876
rect 180804 325874 181404 325876
rect 216804 325874 217404 325876
rect 252804 325874 253404 325876
rect 288804 325874 289404 325876
rect 324804 325874 325404 325876
rect 360804 325874 361404 325876
rect 396804 325874 397404 325876
rect 432804 325874 433404 325876
rect 468804 325874 469404 325876
rect 504804 325874 505404 325876
rect 540804 325874 541404 325876
rect 576804 325874 577404 325876
rect 585320 325874 585920 325876
rect -8576 319276 -7976 319278
rect 29604 319276 30204 319278
rect 65604 319276 66204 319278
rect 101604 319276 102204 319278
rect 137604 319276 138204 319278
rect 173604 319276 174204 319278
rect 209604 319276 210204 319278
rect 245604 319276 246204 319278
rect 281604 319276 282204 319278
rect 317604 319276 318204 319278
rect 353604 319276 354204 319278
rect 389604 319276 390204 319278
rect 425604 319276 426204 319278
rect 461604 319276 462204 319278
rect 497604 319276 498204 319278
rect 533604 319276 534204 319278
rect 569604 319276 570204 319278
rect 591900 319276 592500 319278
rect -8576 319254 592500 319276
rect -8576 319018 -8394 319254
rect -8158 319018 29786 319254
rect 30022 319018 65786 319254
rect 66022 319018 101786 319254
rect 102022 319018 137786 319254
rect 138022 319018 173786 319254
rect 174022 319018 209786 319254
rect 210022 319018 245786 319254
rect 246022 319018 281786 319254
rect 282022 319018 317786 319254
rect 318022 319018 353786 319254
rect 354022 319018 389786 319254
rect 390022 319018 425786 319254
rect 426022 319018 461786 319254
rect 462022 319018 497786 319254
rect 498022 319018 533786 319254
rect 534022 319018 569786 319254
rect 570022 319018 592082 319254
rect 592318 319018 592500 319254
rect -8576 318934 592500 319018
rect -8576 318698 -8394 318934
rect -8158 318698 29786 318934
rect 30022 318698 65786 318934
rect 66022 318698 101786 318934
rect 102022 318698 137786 318934
rect 138022 318698 173786 318934
rect 174022 318698 209786 318934
rect 210022 318698 245786 318934
rect 246022 318698 281786 318934
rect 282022 318698 317786 318934
rect 318022 318698 353786 318934
rect 354022 318698 389786 318934
rect 390022 318698 425786 318934
rect 426022 318698 461786 318934
rect 462022 318698 497786 318934
rect 498022 318698 533786 318934
rect 534022 318698 569786 318934
rect 570022 318698 592082 318934
rect 592318 318698 592500 318934
rect -8576 318676 592500 318698
rect -8576 318674 -7976 318676
rect 29604 318674 30204 318676
rect 65604 318674 66204 318676
rect 101604 318674 102204 318676
rect 137604 318674 138204 318676
rect 173604 318674 174204 318676
rect 209604 318674 210204 318676
rect 245604 318674 246204 318676
rect 281604 318674 282204 318676
rect 317604 318674 318204 318676
rect 353604 318674 354204 318676
rect 389604 318674 390204 318676
rect 425604 318674 426204 318676
rect 461604 318674 462204 318676
rect 497604 318674 498204 318676
rect 533604 318674 534204 318676
rect 569604 318674 570204 318676
rect 591900 318674 592500 318676
rect -6696 315676 -6096 315678
rect 26004 315676 26604 315678
rect 62004 315676 62604 315678
rect 98004 315676 98604 315678
rect 134004 315676 134604 315678
rect 170004 315676 170604 315678
rect 206004 315676 206604 315678
rect 242004 315676 242604 315678
rect 278004 315676 278604 315678
rect 314004 315676 314604 315678
rect 350004 315676 350604 315678
rect 386004 315676 386604 315678
rect 422004 315676 422604 315678
rect 458004 315676 458604 315678
rect 494004 315676 494604 315678
rect 530004 315676 530604 315678
rect 566004 315676 566604 315678
rect 590020 315676 590620 315678
rect -6696 315654 590620 315676
rect -6696 315418 -6514 315654
rect -6278 315418 26186 315654
rect 26422 315418 62186 315654
rect 62422 315418 98186 315654
rect 98422 315418 134186 315654
rect 134422 315418 170186 315654
rect 170422 315418 206186 315654
rect 206422 315418 242186 315654
rect 242422 315418 278186 315654
rect 278422 315418 314186 315654
rect 314422 315418 350186 315654
rect 350422 315418 386186 315654
rect 386422 315418 422186 315654
rect 422422 315418 458186 315654
rect 458422 315418 494186 315654
rect 494422 315418 530186 315654
rect 530422 315418 566186 315654
rect 566422 315418 590202 315654
rect 590438 315418 590620 315654
rect -6696 315334 590620 315418
rect -6696 315098 -6514 315334
rect -6278 315098 26186 315334
rect 26422 315098 62186 315334
rect 62422 315098 98186 315334
rect 98422 315098 134186 315334
rect 134422 315098 170186 315334
rect 170422 315098 206186 315334
rect 206422 315098 242186 315334
rect 242422 315098 278186 315334
rect 278422 315098 314186 315334
rect 314422 315098 350186 315334
rect 350422 315098 386186 315334
rect 386422 315098 422186 315334
rect 422422 315098 458186 315334
rect 458422 315098 494186 315334
rect 494422 315098 530186 315334
rect 530422 315098 566186 315334
rect 566422 315098 590202 315334
rect 590438 315098 590620 315334
rect -6696 315076 590620 315098
rect -6696 315074 -6096 315076
rect 26004 315074 26604 315076
rect 62004 315074 62604 315076
rect 98004 315074 98604 315076
rect 134004 315074 134604 315076
rect 170004 315074 170604 315076
rect 206004 315074 206604 315076
rect 242004 315074 242604 315076
rect 278004 315074 278604 315076
rect 314004 315074 314604 315076
rect 350004 315074 350604 315076
rect 386004 315074 386604 315076
rect 422004 315074 422604 315076
rect 458004 315074 458604 315076
rect 494004 315074 494604 315076
rect 530004 315074 530604 315076
rect 566004 315074 566604 315076
rect 590020 315074 590620 315076
rect -4816 312076 -4216 312078
rect 22404 312076 23004 312078
rect 58404 312076 59004 312078
rect 94404 312076 95004 312078
rect 130404 312076 131004 312078
rect 166404 312076 167004 312078
rect 202404 312076 203004 312078
rect 238404 312076 239004 312078
rect 274404 312076 275004 312078
rect 310404 312076 311004 312078
rect 346404 312076 347004 312078
rect 382404 312076 383004 312078
rect 418404 312076 419004 312078
rect 454404 312076 455004 312078
rect 490404 312076 491004 312078
rect 526404 312076 527004 312078
rect 562404 312076 563004 312078
rect 588140 312076 588740 312078
rect -4816 312054 588740 312076
rect -4816 311818 -4634 312054
rect -4398 311818 22586 312054
rect 22822 311818 58586 312054
rect 58822 311818 94586 312054
rect 94822 311818 130586 312054
rect 130822 311818 166586 312054
rect 166822 311818 202586 312054
rect 202822 311818 238586 312054
rect 238822 311818 274586 312054
rect 274822 311818 310586 312054
rect 310822 311818 346586 312054
rect 346822 311818 382586 312054
rect 382822 311818 418586 312054
rect 418822 311818 454586 312054
rect 454822 311818 490586 312054
rect 490822 311818 526586 312054
rect 526822 311818 562586 312054
rect 562822 311818 588322 312054
rect 588558 311818 588740 312054
rect -4816 311734 588740 311818
rect -4816 311498 -4634 311734
rect -4398 311498 22586 311734
rect 22822 311498 58586 311734
rect 58822 311498 94586 311734
rect 94822 311498 130586 311734
rect 130822 311498 166586 311734
rect 166822 311498 202586 311734
rect 202822 311498 238586 311734
rect 238822 311498 274586 311734
rect 274822 311498 310586 311734
rect 310822 311498 346586 311734
rect 346822 311498 382586 311734
rect 382822 311498 418586 311734
rect 418822 311498 454586 311734
rect 454822 311498 490586 311734
rect 490822 311498 526586 311734
rect 526822 311498 562586 311734
rect 562822 311498 588322 311734
rect 588558 311498 588740 311734
rect -4816 311476 588740 311498
rect -4816 311474 -4216 311476
rect 22404 311474 23004 311476
rect 58404 311474 59004 311476
rect 94404 311474 95004 311476
rect 130404 311474 131004 311476
rect 166404 311474 167004 311476
rect 202404 311474 203004 311476
rect 238404 311474 239004 311476
rect 274404 311474 275004 311476
rect 310404 311474 311004 311476
rect 346404 311474 347004 311476
rect 382404 311474 383004 311476
rect 418404 311474 419004 311476
rect 454404 311474 455004 311476
rect 490404 311474 491004 311476
rect 526404 311474 527004 311476
rect 562404 311474 563004 311476
rect 588140 311474 588740 311476
rect -2936 308476 -2336 308478
rect 18804 308476 19404 308478
rect 54804 308476 55404 308478
rect 90804 308476 91404 308478
rect 126804 308476 127404 308478
rect 162804 308476 163404 308478
rect 198804 308476 199404 308478
rect 234804 308476 235404 308478
rect 270804 308476 271404 308478
rect 306804 308476 307404 308478
rect 342804 308476 343404 308478
rect 378804 308476 379404 308478
rect 414804 308476 415404 308478
rect 450804 308476 451404 308478
rect 486804 308476 487404 308478
rect 522804 308476 523404 308478
rect 558804 308476 559404 308478
rect 586260 308476 586860 308478
rect -2936 308454 586860 308476
rect -2936 308218 -2754 308454
rect -2518 308218 18986 308454
rect 19222 308218 54986 308454
rect 55222 308218 90986 308454
rect 91222 308218 126986 308454
rect 127222 308218 162986 308454
rect 163222 308218 198986 308454
rect 199222 308218 234986 308454
rect 235222 308218 270986 308454
rect 271222 308218 306986 308454
rect 307222 308218 342986 308454
rect 343222 308218 378986 308454
rect 379222 308218 414986 308454
rect 415222 308218 450986 308454
rect 451222 308218 486986 308454
rect 487222 308218 522986 308454
rect 523222 308218 558986 308454
rect 559222 308218 586442 308454
rect 586678 308218 586860 308454
rect -2936 308134 586860 308218
rect -2936 307898 -2754 308134
rect -2518 307898 18986 308134
rect 19222 307898 54986 308134
rect 55222 307898 90986 308134
rect 91222 307898 126986 308134
rect 127222 307898 162986 308134
rect 163222 307898 198986 308134
rect 199222 307898 234986 308134
rect 235222 307898 270986 308134
rect 271222 307898 306986 308134
rect 307222 307898 342986 308134
rect 343222 307898 378986 308134
rect 379222 307898 414986 308134
rect 415222 307898 450986 308134
rect 451222 307898 486986 308134
rect 487222 307898 522986 308134
rect 523222 307898 558986 308134
rect 559222 307898 586442 308134
rect 586678 307898 586860 308134
rect -2936 307876 586860 307898
rect -2936 307874 -2336 307876
rect 18804 307874 19404 307876
rect 54804 307874 55404 307876
rect 90804 307874 91404 307876
rect 126804 307874 127404 307876
rect 162804 307874 163404 307876
rect 198804 307874 199404 307876
rect 234804 307874 235404 307876
rect 270804 307874 271404 307876
rect 306804 307874 307404 307876
rect 342804 307874 343404 307876
rect 378804 307874 379404 307876
rect 414804 307874 415404 307876
rect 450804 307874 451404 307876
rect 486804 307874 487404 307876
rect 522804 307874 523404 307876
rect 558804 307874 559404 307876
rect 586260 307874 586860 307876
rect -7636 301276 -7036 301278
rect 11604 301276 12204 301278
rect 47604 301276 48204 301278
rect 83604 301276 84204 301278
rect 119604 301276 120204 301278
rect 155604 301276 156204 301278
rect 191604 301276 192204 301278
rect 227604 301276 228204 301278
rect 263604 301276 264204 301278
rect 299604 301276 300204 301278
rect 335604 301276 336204 301278
rect 371604 301276 372204 301278
rect 407604 301276 408204 301278
rect 443604 301276 444204 301278
rect 479604 301276 480204 301278
rect 515604 301276 516204 301278
rect 551604 301276 552204 301278
rect 590960 301276 591560 301278
rect -8576 301254 592500 301276
rect -8576 301018 -7454 301254
rect -7218 301018 11786 301254
rect 12022 301018 47786 301254
rect 48022 301018 83786 301254
rect 84022 301018 119786 301254
rect 120022 301018 155786 301254
rect 156022 301018 191786 301254
rect 192022 301018 227786 301254
rect 228022 301018 263786 301254
rect 264022 301018 299786 301254
rect 300022 301018 335786 301254
rect 336022 301018 371786 301254
rect 372022 301018 407786 301254
rect 408022 301018 443786 301254
rect 444022 301018 479786 301254
rect 480022 301018 515786 301254
rect 516022 301018 551786 301254
rect 552022 301018 591142 301254
rect 591378 301018 592500 301254
rect -8576 300934 592500 301018
rect -8576 300698 -7454 300934
rect -7218 300698 11786 300934
rect 12022 300698 47786 300934
rect 48022 300698 83786 300934
rect 84022 300698 119786 300934
rect 120022 300698 155786 300934
rect 156022 300698 191786 300934
rect 192022 300698 227786 300934
rect 228022 300698 263786 300934
rect 264022 300698 299786 300934
rect 300022 300698 335786 300934
rect 336022 300698 371786 300934
rect 372022 300698 407786 300934
rect 408022 300698 443786 300934
rect 444022 300698 479786 300934
rect 480022 300698 515786 300934
rect 516022 300698 551786 300934
rect 552022 300698 591142 300934
rect 591378 300698 592500 300934
rect -8576 300676 592500 300698
rect -7636 300674 -7036 300676
rect 11604 300674 12204 300676
rect 47604 300674 48204 300676
rect 83604 300674 84204 300676
rect 119604 300674 120204 300676
rect 155604 300674 156204 300676
rect 191604 300674 192204 300676
rect 227604 300674 228204 300676
rect 263604 300674 264204 300676
rect 299604 300674 300204 300676
rect 335604 300674 336204 300676
rect 371604 300674 372204 300676
rect 407604 300674 408204 300676
rect 443604 300674 444204 300676
rect 479604 300674 480204 300676
rect 515604 300674 516204 300676
rect 551604 300674 552204 300676
rect 590960 300674 591560 300676
rect -5756 297676 -5156 297678
rect 8004 297676 8604 297678
rect 44004 297676 44604 297678
rect 80004 297676 80604 297678
rect 116004 297676 116604 297678
rect 152004 297676 152604 297678
rect 188004 297676 188604 297678
rect 224004 297676 224604 297678
rect 260004 297676 260604 297678
rect 296004 297676 296604 297678
rect 332004 297676 332604 297678
rect 368004 297676 368604 297678
rect 404004 297676 404604 297678
rect 440004 297676 440604 297678
rect 476004 297676 476604 297678
rect 512004 297676 512604 297678
rect 548004 297676 548604 297678
rect 589080 297676 589680 297678
rect -6696 297654 590620 297676
rect -6696 297418 -5574 297654
rect -5338 297418 8186 297654
rect 8422 297418 44186 297654
rect 44422 297418 80186 297654
rect 80422 297418 116186 297654
rect 116422 297418 152186 297654
rect 152422 297418 188186 297654
rect 188422 297418 224186 297654
rect 224422 297418 260186 297654
rect 260422 297418 296186 297654
rect 296422 297418 332186 297654
rect 332422 297418 368186 297654
rect 368422 297418 404186 297654
rect 404422 297418 440186 297654
rect 440422 297418 476186 297654
rect 476422 297418 512186 297654
rect 512422 297418 548186 297654
rect 548422 297418 589262 297654
rect 589498 297418 590620 297654
rect -6696 297334 590620 297418
rect -6696 297098 -5574 297334
rect -5338 297098 8186 297334
rect 8422 297098 44186 297334
rect 44422 297098 80186 297334
rect 80422 297098 116186 297334
rect 116422 297098 152186 297334
rect 152422 297098 188186 297334
rect 188422 297098 224186 297334
rect 224422 297098 260186 297334
rect 260422 297098 296186 297334
rect 296422 297098 332186 297334
rect 332422 297098 368186 297334
rect 368422 297098 404186 297334
rect 404422 297098 440186 297334
rect 440422 297098 476186 297334
rect 476422 297098 512186 297334
rect 512422 297098 548186 297334
rect 548422 297098 589262 297334
rect 589498 297098 590620 297334
rect -6696 297076 590620 297098
rect -5756 297074 -5156 297076
rect 8004 297074 8604 297076
rect 44004 297074 44604 297076
rect 80004 297074 80604 297076
rect 116004 297074 116604 297076
rect 152004 297074 152604 297076
rect 188004 297074 188604 297076
rect 224004 297074 224604 297076
rect 260004 297074 260604 297076
rect 296004 297074 296604 297076
rect 332004 297074 332604 297076
rect 368004 297074 368604 297076
rect 404004 297074 404604 297076
rect 440004 297074 440604 297076
rect 476004 297074 476604 297076
rect 512004 297074 512604 297076
rect 548004 297074 548604 297076
rect 589080 297074 589680 297076
rect -3876 294076 -3276 294078
rect 4404 294076 5004 294078
rect 40404 294076 41004 294078
rect 76404 294076 77004 294078
rect 112404 294076 113004 294078
rect 148404 294076 149004 294078
rect 184404 294076 185004 294078
rect 220404 294076 221004 294078
rect 256404 294076 257004 294078
rect 292404 294076 293004 294078
rect 328404 294076 329004 294078
rect 364404 294076 365004 294078
rect 400404 294076 401004 294078
rect 436404 294076 437004 294078
rect 472404 294076 473004 294078
rect 508404 294076 509004 294078
rect 544404 294076 545004 294078
rect 580404 294076 581004 294078
rect 587200 294076 587800 294078
rect -4816 294054 588740 294076
rect -4816 293818 -3694 294054
rect -3458 293818 4586 294054
rect 4822 293818 40586 294054
rect 40822 293818 76586 294054
rect 76822 293818 112586 294054
rect 112822 293818 148586 294054
rect 148822 293818 184586 294054
rect 184822 293818 220586 294054
rect 220822 293818 256586 294054
rect 256822 293818 292586 294054
rect 292822 293818 328586 294054
rect 328822 293818 364586 294054
rect 364822 293818 400586 294054
rect 400822 293818 436586 294054
rect 436822 293818 472586 294054
rect 472822 293818 508586 294054
rect 508822 293818 544586 294054
rect 544822 293818 580586 294054
rect 580822 293818 587382 294054
rect 587618 293818 588740 294054
rect -4816 293734 588740 293818
rect -4816 293498 -3694 293734
rect -3458 293498 4586 293734
rect 4822 293498 40586 293734
rect 40822 293498 76586 293734
rect 76822 293498 112586 293734
rect 112822 293498 148586 293734
rect 148822 293498 184586 293734
rect 184822 293498 220586 293734
rect 220822 293498 256586 293734
rect 256822 293498 292586 293734
rect 292822 293498 328586 293734
rect 328822 293498 364586 293734
rect 364822 293498 400586 293734
rect 400822 293498 436586 293734
rect 436822 293498 472586 293734
rect 472822 293498 508586 293734
rect 508822 293498 544586 293734
rect 544822 293498 580586 293734
rect 580822 293498 587382 293734
rect 587618 293498 588740 293734
rect -4816 293476 588740 293498
rect -3876 293474 -3276 293476
rect 4404 293474 5004 293476
rect 40404 293474 41004 293476
rect 76404 293474 77004 293476
rect 112404 293474 113004 293476
rect 148404 293474 149004 293476
rect 184404 293474 185004 293476
rect 220404 293474 221004 293476
rect 256404 293474 257004 293476
rect 292404 293474 293004 293476
rect 328404 293474 329004 293476
rect 364404 293474 365004 293476
rect 400404 293474 401004 293476
rect 436404 293474 437004 293476
rect 472404 293474 473004 293476
rect 508404 293474 509004 293476
rect 544404 293474 545004 293476
rect 580404 293474 581004 293476
rect 587200 293474 587800 293476
rect -1996 290476 -1396 290478
rect 804 290476 1404 290478
rect 36804 290476 37404 290478
rect 72804 290476 73404 290478
rect 108804 290476 109404 290478
rect 144804 290476 145404 290478
rect 180804 290476 181404 290478
rect 216804 290476 217404 290478
rect 252804 290476 253404 290478
rect 288804 290476 289404 290478
rect 324804 290476 325404 290478
rect 360804 290476 361404 290478
rect 396804 290476 397404 290478
rect 432804 290476 433404 290478
rect 468804 290476 469404 290478
rect 504804 290476 505404 290478
rect 540804 290476 541404 290478
rect 576804 290476 577404 290478
rect 585320 290476 585920 290478
rect -2936 290454 586860 290476
rect -2936 290218 -1814 290454
rect -1578 290218 986 290454
rect 1222 290218 36986 290454
rect 37222 290218 72986 290454
rect 73222 290218 108986 290454
rect 109222 290218 144986 290454
rect 145222 290218 180986 290454
rect 181222 290218 216986 290454
rect 217222 290218 252986 290454
rect 253222 290218 288986 290454
rect 289222 290218 324986 290454
rect 325222 290218 360986 290454
rect 361222 290218 396986 290454
rect 397222 290218 432986 290454
rect 433222 290218 468986 290454
rect 469222 290218 504986 290454
rect 505222 290218 540986 290454
rect 541222 290218 576986 290454
rect 577222 290218 585502 290454
rect 585738 290218 586860 290454
rect -2936 290134 586860 290218
rect -2936 289898 -1814 290134
rect -1578 289898 986 290134
rect 1222 289898 36986 290134
rect 37222 289898 72986 290134
rect 73222 289898 108986 290134
rect 109222 289898 144986 290134
rect 145222 289898 180986 290134
rect 181222 289898 216986 290134
rect 217222 289898 252986 290134
rect 253222 289898 288986 290134
rect 289222 289898 324986 290134
rect 325222 289898 360986 290134
rect 361222 289898 396986 290134
rect 397222 289898 432986 290134
rect 433222 289898 468986 290134
rect 469222 289898 504986 290134
rect 505222 289898 540986 290134
rect 541222 289898 576986 290134
rect 577222 289898 585502 290134
rect 585738 289898 586860 290134
rect -2936 289876 586860 289898
rect -1996 289874 -1396 289876
rect 804 289874 1404 289876
rect 36804 289874 37404 289876
rect 72804 289874 73404 289876
rect 108804 289874 109404 289876
rect 144804 289874 145404 289876
rect 180804 289874 181404 289876
rect 216804 289874 217404 289876
rect 252804 289874 253404 289876
rect 288804 289874 289404 289876
rect 324804 289874 325404 289876
rect 360804 289874 361404 289876
rect 396804 289874 397404 289876
rect 432804 289874 433404 289876
rect 468804 289874 469404 289876
rect 504804 289874 505404 289876
rect 540804 289874 541404 289876
rect 576804 289874 577404 289876
rect 585320 289874 585920 289876
rect -8576 283276 -7976 283278
rect 29604 283276 30204 283278
rect 65604 283276 66204 283278
rect 101604 283276 102204 283278
rect 137604 283276 138204 283278
rect 173604 283276 174204 283278
rect 209604 283276 210204 283278
rect 245604 283276 246204 283278
rect 281604 283276 282204 283278
rect 317604 283276 318204 283278
rect 353604 283276 354204 283278
rect 389604 283276 390204 283278
rect 425604 283276 426204 283278
rect 461604 283276 462204 283278
rect 497604 283276 498204 283278
rect 533604 283276 534204 283278
rect 569604 283276 570204 283278
rect 591900 283276 592500 283278
rect -8576 283254 592500 283276
rect -8576 283018 -8394 283254
rect -8158 283018 29786 283254
rect 30022 283018 65786 283254
rect 66022 283018 101786 283254
rect 102022 283018 137786 283254
rect 138022 283018 173786 283254
rect 174022 283018 209786 283254
rect 210022 283018 245786 283254
rect 246022 283018 281786 283254
rect 282022 283018 317786 283254
rect 318022 283018 353786 283254
rect 354022 283018 389786 283254
rect 390022 283018 425786 283254
rect 426022 283018 461786 283254
rect 462022 283018 497786 283254
rect 498022 283018 533786 283254
rect 534022 283018 569786 283254
rect 570022 283018 592082 283254
rect 592318 283018 592500 283254
rect -8576 282934 592500 283018
rect -8576 282698 -8394 282934
rect -8158 282698 29786 282934
rect 30022 282698 65786 282934
rect 66022 282698 101786 282934
rect 102022 282698 137786 282934
rect 138022 282698 173786 282934
rect 174022 282698 209786 282934
rect 210022 282698 245786 282934
rect 246022 282698 281786 282934
rect 282022 282698 317786 282934
rect 318022 282698 353786 282934
rect 354022 282698 389786 282934
rect 390022 282698 425786 282934
rect 426022 282698 461786 282934
rect 462022 282698 497786 282934
rect 498022 282698 533786 282934
rect 534022 282698 569786 282934
rect 570022 282698 592082 282934
rect 592318 282698 592500 282934
rect -8576 282676 592500 282698
rect -8576 282674 -7976 282676
rect 29604 282674 30204 282676
rect 65604 282674 66204 282676
rect 101604 282674 102204 282676
rect 137604 282674 138204 282676
rect 173604 282674 174204 282676
rect 209604 282674 210204 282676
rect 245604 282674 246204 282676
rect 281604 282674 282204 282676
rect 317604 282674 318204 282676
rect 353604 282674 354204 282676
rect 389604 282674 390204 282676
rect 425604 282674 426204 282676
rect 461604 282674 462204 282676
rect 497604 282674 498204 282676
rect 533604 282674 534204 282676
rect 569604 282674 570204 282676
rect 591900 282674 592500 282676
rect -6696 279676 -6096 279678
rect 26004 279676 26604 279678
rect 62004 279676 62604 279678
rect 98004 279676 98604 279678
rect 134004 279676 134604 279678
rect 170004 279676 170604 279678
rect 206004 279676 206604 279678
rect 242004 279676 242604 279678
rect 278004 279676 278604 279678
rect 314004 279676 314604 279678
rect 350004 279676 350604 279678
rect 386004 279676 386604 279678
rect 422004 279676 422604 279678
rect 458004 279676 458604 279678
rect 494004 279676 494604 279678
rect 530004 279676 530604 279678
rect 566004 279676 566604 279678
rect 590020 279676 590620 279678
rect -6696 279654 590620 279676
rect -6696 279418 -6514 279654
rect -6278 279418 26186 279654
rect 26422 279418 62186 279654
rect 62422 279418 98186 279654
rect 98422 279418 134186 279654
rect 134422 279418 170186 279654
rect 170422 279418 206186 279654
rect 206422 279418 242186 279654
rect 242422 279418 278186 279654
rect 278422 279418 314186 279654
rect 314422 279418 350186 279654
rect 350422 279418 386186 279654
rect 386422 279418 422186 279654
rect 422422 279418 458186 279654
rect 458422 279418 494186 279654
rect 494422 279418 530186 279654
rect 530422 279418 566186 279654
rect 566422 279418 590202 279654
rect 590438 279418 590620 279654
rect -6696 279334 590620 279418
rect -6696 279098 -6514 279334
rect -6278 279098 26186 279334
rect 26422 279098 62186 279334
rect 62422 279098 98186 279334
rect 98422 279098 134186 279334
rect 134422 279098 170186 279334
rect 170422 279098 206186 279334
rect 206422 279098 242186 279334
rect 242422 279098 278186 279334
rect 278422 279098 314186 279334
rect 314422 279098 350186 279334
rect 350422 279098 386186 279334
rect 386422 279098 422186 279334
rect 422422 279098 458186 279334
rect 458422 279098 494186 279334
rect 494422 279098 530186 279334
rect 530422 279098 566186 279334
rect 566422 279098 590202 279334
rect 590438 279098 590620 279334
rect -6696 279076 590620 279098
rect -6696 279074 -6096 279076
rect 26004 279074 26604 279076
rect 62004 279074 62604 279076
rect 98004 279074 98604 279076
rect 134004 279074 134604 279076
rect 170004 279074 170604 279076
rect 206004 279074 206604 279076
rect 242004 279074 242604 279076
rect 278004 279074 278604 279076
rect 314004 279074 314604 279076
rect 350004 279074 350604 279076
rect 386004 279074 386604 279076
rect 422004 279074 422604 279076
rect 458004 279074 458604 279076
rect 494004 279074 494604 279076
rect 530004 279074 530604 279076
rect 566004 279074 566604 279076
rect 590020 279074 590620 279076
rect -4816 276076 -4216 276078
rect 22404 276076 23004 276078
rect 58404 276076 59004 276078
rect 94404 276076 95004 276078
rect 130404 276076 131004 276078
rect 166404 276076 167004 276078
rect 202404 276076 203004 276078
rect 238404 276076 239004 276078
rect 274404 276076 275004 276078
rect 310404 276076 311004 276078
rect 346404 276076 347004 276078
rect 382404 276076 383004 276078
rect 418404 276076 419004 276078
rect 454404 276076 455004 276078
rect 490404 276076 491004 276078
rect 526404 276076 527004 276078
rect 562404 276076 563004 276078
rect 588140 276076 588740 276078
rect -4816 276054 588740 276076
rect -4816 275818 -4634 276054
rect -4398 275818 22586 276054
rect 22822 275818 58586 276054
rect 58822 275818 94586 276054
rect 94822 275818 130586 276054
rect 130822 275818 166586 276054
rect 166822 275818 202586 276054
rect 202822 275818 238586 276054
rect 238822 275818 274586 276054
rect 274822 275818 310586 276054
rect 310822 275818 346586 276054
rect 346822 275818 382586 276054
rect 382822 275818 418586 276054
rect 418822 275818 454586 276054
rect 454822 275818 490586 276054
rect 490822 275818 526586 276054
rect 526822 275818 562586 276054
rect 562822 275818 588322 276054
rect 588558 275818 588740 276054
rect -4816 275734 588740 275818
rect -4816 275498 -4634 275734
rect -4398 275498 22586 275734
rect 22822 275498 58586 275734
rect 58822 275498 94586 275734
rect 94822 275498 130586 275734
rect 130822 275498 166586 275734
rect 166822 275498 202586 275734
rect 202822 275498 238586 275734
rect 238822 275498 274586 275734
rect 274822 275498 310586 275734
rect 310822 275498 346586 275734
rect 346822 275498 382586 275734
rect 382822 275498 418586 275734
rect 418822 275498 454586 275734
rect 454822 275498 490586 275734
rect 490822 275498 526586 275734
rect 526822 275498 562586 275734
rect 562822 275498 588322 275734
rect 588558 275498 588740 275734
rect -4816 275476 588740 275498
rect -4816 275474 -4216 275476
rect 22404 275474 23004 275476
rect 58404 275474 59004 275476
rect 94404 275474 95004 275476
rect 130404 275474 131004 275476
rect 166404 275474 167004 275476
rect 202404 275474 203004 275476
rect 238404 275474 239004 275476
rect 274404 275474 275004 275476
rect 310404 275474 311004 275476
rect 346404 275474 347004 275476
rect 382404 275474 383004 275476
rect 418404 275474 419004 275476
rect 454404 275474 455004 275476
rect 490404 275474 491004 275476
rect 526404 275474 527004 275476
rect 562404 275474 563004 275476
rect 588140 275474 588740 275476
rect -2936 272476 -2336 272478
rect 18804 272476 19404 272478
rect 54804 272476 55404 272478
rect 90804 272476 91404 272478
rect 126804 272476 127404 272478
rect 162804 272476 163404 272478
rect 198804 272476 199404 272478
rect 234804 272476 235404 272478
rect 270804 272476 271404 272478
rect 306804 272476 307404 272478
rect 342804 272476 343404 272478
rect 378804 272476 379404 272478
rect 414804 272476 415404 272478
rect 450804 272476 451404 272478
rect 486804 272476 487404 272478
rect 522804 272476 523404 272478
rect 558804 272476 559404 272478
rect 586260 272476 586860 272478
rect -2936 272454 586860 272476
rect -2936 272218 -2754 272454
rect -2518 272218 18986 272454
rect 19222 272218 54986 272454
rect 55222 272218 90986 272454
rect 91222 272218 126986 272454
rect 127222 272218 162986 272454
rect 163222 272218 198986 272454
rect 199222 272218 234986 272454
rect 235222 272218 270986 272454
rect 271222 272218 306986 272454
rect 307222 272218 342986 272454
rect 343222 272218 378986 272454
rect 379222 272218 414986 272454
rect 415222 272218 450986 272454
rect 451222 272218 486986 272454
rect 487222 272218 522986 272454
rect 523222 272218 558986 272454
rect 559222 272218 586442 272454
rect 586678 272218 586860 272454
rect -2936 272134 586860 272218
rect -2936 271898 -2754 272134
rect -2518 271898 18986 272134
rect 19222 271898 54986 272134
rect 55222 271898 90986 272134
rect 91222 271898 126986 272134
rect 127222 271898 162986 272134
rect 163222 271898 198986 272134
rect 199222 271898 234986 272134
rect 235222 271898 270986 272134
rect 271222 271898 306986 272134
rect 307222 271898 342986 272134
rect 343222 271898 378986 272134
rect 379222 271898 414986 272134
rect 415222 271898 450986 272134
rect 451222 271898 486986 272134
rect 487222 271898 522986 272134
rect 523222 271898 558986 272134
rect 559222 271898 586442 272134
rect 586678 271898 586860 272134
rect -2936 271876 586860 271898
rect -2936 271874 -2336 271876
rect 18804 271874 19404 271876
rect 54804 271874 55404 271876
rect 90804 271874 91404 271876
rect 126804 271874 127404 271876
rect 162804 271874 163404 271876
rect 198804 271874 199404 271876
rect 234804 271874 235404 271876
rect 270804 271874 271404 271876
rect 306804 271874 307404 271876
rect 342804 271874 343404 271876
rect 378804 271874 379404 271876
rect 414804 271874 415404 271876
rect 450804 271874 451404 271876
rect 486804 271874 487404 271876
rect 522804 271874 523404 271876
rect 558804 271874 559404 271876
rect 586260 271874 586860 271876
rect -7636 265276 -7036 265278
rect 11604 265276 12204 265278
rect 47604 265276 48204 265278
rect 83604 265276 84204 265278
rect 119604 265276 120204 265278
rect 155604 265276 156204 265278
rect 191604 265276 192204 265278
rect 227604 265276 228204 265278
rect 263604 265276 264204 265278
rect 299604 265276 300204 265278
rect 335604 265276 336204 265278
rect 371604 265276 372204 265278
rect 407604 265276 408204 265278
rect 443604 265276 444204 265278
rect 479604 265276 480204 265278
rect 515604 265276 516204 265278
rect 551604 265276 552204 265278
rect 590960 265276 591560 265278
rect -8576 265254 592500 265276
rect -8576 265018 -7454 265254
rect -7218 265018 11786 265254
rect 12022 265018 47786 265254
rect 48022 265018 83786 265254
rect 84022 265018 119786 265254
rect 120022 265018 155786 265254
rect 156022 265018 191786 265254
rect 192022 265018 227786 265254
rect 228022 265018 263786 265254
rect 264022 265018 299786 265254
rect 300022 265018 335786 265254
rect 336022 265018 371786 265254
rect 372022 265018 407786 265254
rect 408022 265018 443786 265254
rect 444022 265018 479786 265254
rect 480022 265018 515786 265254
rect 516022 265018 551786 265254
rect 552022 265018 591142 265254
rect 591378 265018 592500 265254
rect -8576 264934 592500 265018
rect -8576 264698 -7454 264934
rect -7218 264698 11786 264934
rect 12022 264698 47786 264934
rect 48022 264698 83786 264934
rect 84022 264698 119786 264934
rect 120022 264698 155786 264934
rect 156022 264698 191786 264934
rect 192022 264698 227786 264934
rect 228022 264698 263786 264934
rect 264022 264698 299786 264934
rect 300022 264698 335786 264934
rect 336022 264698 371786 264934
rect 372022 264698 407786 264934
rect 408022 264698 443786 264934
rect 444022 264698 479786 264934
rect 480022 264698 515786 264934
rect 516022 264698 551786 264934
rect 552022 264698 591142 264934
rect 591378 264698 592500 264934
rect -8576 264676 592500 264698
rect -7636 264674 -7036 264676
rect 11604 264674 12204 264676
rect 47604 264674 48204 264676
rect 83604 264674 84204 264676
rect 119604 264674 120204 264676
rect 155604 264674 156204 264676
rect 191604 264674 192204 264676
rect 227604 264674 228204 264676
rect 263604 264674 264204 264676
rect 299604 264674 300204 264676
rect 335604 264674 336204 264676
rect 371604 264674 372204 264676
rect 407604 264674 408204 264676
rect 443604 264674 444204 264676
rect 479604 264674 480204 264676
rect 515604 264674 516204 264676
rect 551604 264674 552204 264676
rect 590960 264674 591560 264676
rect -5756 261676 -5156 261678
rect 8004 261676 8604 261678
rect 44004 261676 44604 261678
rect 80004 261676 80604 261678
rect 116004 261676 116604 261678
rect 152004 261676 152604 261678
rect 188004 261676 188604 261678
rect 224004 261676 224604 261678
rect 260004 261676 260604 261678
rect 296004 261676 296604 261678
rect 332004 261676 332604 261678
rect 368004 261676 368604 261678
rect 404004 261676 404604 261678
rect 440004 261676 440604 261678
rect 476004 261676 476604 261678
rect 512004 261676 512604 261678
rect 548004 261676 548604 261678
rect 589080 261676 589680 261678
rect -6696 261654 590620 261676
rect -6696 261418 -5574 261654
rect -5338 261418 8186 261654
rect 8422 261418 44186 261654
rect 44422 261418 80186 261654
rect 80422 261418 116186 261654
rect 116422 261418 152186 261654
rect 152422 261418 188186 261654
rect 188422 261418 224186 261654
rect 224422 261418 260186 261654
rect 260422 261418 296186 261654
rect 296422 261418 332186 261654
rect 332422 261418 368186 261654
rect 368422 261418 404186 261654
rect 404422 261418 440186 261654
rect 440422 261418 476186 261654
rect 476422 261418 512186 261654
rect 512422 261418 548186 261654
rect 548422 261418 589262 261654
rect 589498 261418 590620 261654
rect -6696 261334 590620 261418
rect -6696 261098 -5574 261334
rect -5338 261098 8186 261334
rect 8422 261098 44186 261334
rect 44422 261098 80186 261334
rect 80422 261098 116186 261334
rect 116422 261098 152186 261334
rect 152422 261098 188186 261334
rect 188422 261098 224186 261334
rect 224422 261098 260186 261334
rect 260422 261098 296186 261334
rect 296422 261098 332186 261334
rect 332422 261098 368186 261334
rect 368422 261098 404186 261334
rect 404422 261098 440186 261334
rect 440422 261098 476186 261334
rect 476422 261098 512186 261334
rect 512422 261098 548186 261334
rect 548422 261098 589262 261334
rect 589498 261098 590620 261334
rect -6696 261076 590620 261098
rect -5756 261074 -5156 261076
rect 8004 261074 8604 261076
rect 44004 261074 44604 261076
rect 80004 261074 80604 261076
rect 116004 261074 116604 261076
rect 152004 261074 152604 261076
rect 188004 261074 188604 261076
rect 224004 261074 224604 261076
rect 260004 261074 260604 261076
rect 296004 261074 296604 261076
rect 332004 261074 332604 261076
rect 368004 261074 368604 261076
rect 404004 261074 404604 261076
rect 440004 261074 440604 261076
rect 476004 261074 476604 261076
rect 512004 261074 512604 261076
rect 548004 261074 548604 261076
rect 589080 261074 589680 261076
rect -3876 258076 -3276 258078
rect 4404 258076 5004 258078
rect 40404 258076 41004 258078
rect 76404 258076 77004 258078
rect 112404 258076 113004 258078
rect 148404 258076 149004 258078
rect 184404 258076 185004 258078
rect 220404 258076 221004 258078
rect 256404 258076 257004 258078
rect 292404 258076 293004 258078
rect 328404 258076 329004 258078
rect 364404 258076 365004 258078
rect 400404 258076 401004 258078
rect 436404 258076 437004 258078
rect 472404 258076 473004 258078
rect 508404 258076 509004 258078
rect 544404 258076 545004 258078
rect 580404 258076 581004 258078
rect 587200 258076 587800 258078
rect -4816 258054 588740 258076
rect -4816 257818 -3694 258054
rect -3458 257818 4586 258054
rect 4822 257818 40586 258054
rect 40822 257818 76586 258054
rect 76822 257818 112586 258054
rect 112822 257818 148586 258054
rect 148822 257818 184586 258054
rect 184822 257818 220586 258054
rect 220822 257818 256586 258054
rect 256822 257818 292586 258054
rect 292822 257818 328586 258054
rect 328822 257818 364586 258054
rect 364822 257818 400586 258054
rect 400822 257818 436586 258054
rect 436822 257818 472586 258054
rect 472822 257818 508586 258054
rect 508822 257818 544586 258054
rect 544822 257818 580586 258054
rect 580822 257818 587382 258054
rect 587618 257818 588740 258054
rect -4816 257734 588740 257818
rect -4816 257498 -3694 257734
rect -3458 257498 4586 257734
rect 4822 257498 40586 257734
rect 40822 257498 76586 257734
rect 76822 257498 112586 257734
rect 112822 257498 148586 257734
rect 148822 257498 184586 257734
rect 184822 257498 220586 257734
rect 220822 257498 256586 257734
rect 256822 257498 292586 257734
rect 292822 257498 328586 257734
rect 328822 257498 364586 257734
rect 364822 257498 400586 257734
rect 400822 257498 436586 257734
rect 436822 257498 472586 257734
rect 472822 257498 508586 257734
rect 508822 257498 544586 257734
rect 544822 257498 580586 257734
rect 580822 257498 587382 257734
rect 587618 257498 588740 257734
rect -4816 257476 588740 257498
rect -3876 257474 -3276 257476
rect 4404 257474 5004 257476
rect 40404 257474 41004 257476
rect 76404 257474 77004 257476
rect 112404 257474 113004 257476
rect 148404 257474 149004 257476
rect 184404 257474 185004 257476
rect 220404 257474 221004 257476
rect 256404 257474 257004 257476
rect 292404 257474 293004 257476
rect 328404 257474 329004 257476
rect 364404 257474 365004 257476
rect 400404 257474 401004 257476
rect 436404 257474 437004 257476
rect 472404 257474 473004 257476
rect 508404 257474 509004 257476
rect 544404 257474 545004 257476
rect 580404 257474 581004 257476
rect 587200 257474 587800 257476
rect -1996 254476 -1396 254478
rect 804 254476 1404 254478
rect 36804 254476 37404 254478
rect 72804 254476 73404 254478
rect 108804 254476 109404 254478
rect 144804 254476 145404 254478
rect 180804 254476 181404 254478
rect 216804 254476 217404 254478
rect 252804 254476 253404 254478
rect 288804 254476 289404 254478
rect 324804 254476 325404 254478
rect 360804 254476 361404 254478
rect 396804 254476 397404 254478
rect 432804 254476 433404 254478
rect 468804 254476 469404 254478
rect 504804 254476 505404 254478
rect 540804 254476 541404 254478
rect 576804 254476 577404 254478
rect 585320 254476 585920 254478
rect -2936 254454 586860 254476
rect -2936 254218 -1814 254454
rect -1578 254218 986 254454
rect 1222 254218 36986 254454
rect 37222 254218 72986 254454
rect 73222 254218 108986 254454
rect 109222 254218 144986 254454
rect 145222 254218 180986 254454
rect 181222 254218 216986 254454
rect 217222 254218 252986 254454
rect 253222 254218 288986 254454
rect 289222 254218 324986 254454
rect 325222 254218 360986 254454
rect 361222 254218 396986 254454
rect 397222 254218 432986 254454
rect 433222 254218 468986 254454
rect 469222 254218 504986 254454
rect 505222 254218 540986 254454
rect 541222 254218 576986 254454
rect 577222 254218 585502 254454
rect 585738 254218 586860 254454
rect -2936 254134 586860 254218
rect -2936 253898 -1814 254134
rect -1578 253898 986 254134
rect 1222 253898 36986 254134
rect 37222 253898 72986 254134
rect 73222 253898 108986 254134
rect 109222 253898 144986 254134
rect 145222 253898 180986 254134
rect 181222 253898 216986 254134
rect 217222 253898 252986 254134
rect 253222 253898 288986 254134
rect 289222 253898 324986 254134
rect 325222 253898 360986 254134
rect 361222 253898 396986 254134
rect 397222 253898 432986 254134
rect 433222 253898 468986 254134
rect 469222 253898 504986 254134
rect 505222 253898 540986 254134
rect 541222 253898 576986 254134
rect 577222 253898 585502 254134
rect 585738 253898 586860 254134
rect -2936 253876 586860 253898
rect -1996 253874 -1396 253876
rect 804 253874 1404 253876
rect 36804 253874 37404 253876
rect 72804 253874 73404 253876
rect 108804 253874 109404 253876
rect 144804 253874 145404 253876
rect 180804 253874 181404 253876
rect 216804 253874 217404 253876
rect 252804 253874 253404 253876
rect 288804 253874 289404 253876
rect 324804 253874 325404 253876
rect 360804 253874 361404 253876
rect 396804 253874 397404 253876
rect 432804 253874 433404 253876
rect 468804 253874 469404 253876
rect 504804 253874 505404 253876
rect 540804 253874 541404 253876
rect 576804 253874 577404 253876
rect 585320 253874 585920 253876
rect -8576 247276 -7976 247278
rect 29604 247276 30204 247278
rect 65604 247276 66204 247278
rect 101604 247276 102204 247278
rect 137604 247276 138204 247278
rect 173604 247276 174204 247278
rect 209604 247276 210204 247278
rect 245604 247276 246204 247278
rect 281604 247276 282204 247278
rect 317604 247276 318204 247278
rect 353604 247276 354204 247278
rect 389604 247276 390204 247278
rect 425604 247276 426204 247278
rect 461604 247276 462204 247278
rect 497604 247276 498204 247278
rect 533604 247276 534204 247278
rect 569604 247276 570204 247278
rect 591900 247276 592500 247278
rect -8576 247254 592500 247276
rect -8576 247018 -8394 247254
rect -8158 247018 29786 247254
rect 30022 247018 65786 247254
rect 66022 247018 101786 247254
rect 102022 247018 137786 247254
rect 138022 247018 173786 247254
rect 174022 247018 209786 247254
rect 210022 247018 245786 247254
rect 246022 247018 281786 247254
rect 282022 247018 317786 247254
rect 318022 247018 353786 247254
rect 354022 247018 389786 247254
rect 390022 247018 425786 247254
rect 426022 247018 461786 247254
rect 462022 247018 497786 247254
rect 498022 247018 533786 247254
rect 534022 247018 569786 247254
rect 570022 247018 592082 247254
rect 592318 247018 592500 247254
rect -8576 246934 592500 247018
rect -8576 246698 -8394 246934
rect -8158 246698 29786 246934
rect 30022 246698 65786 246934
rect 66022 246698 101786 246934
rect 102022 246698 137786 246934
rect 138022 246698 173786 246934
rect 174022 246698 209786 246934
rect 210022 246698 245786 246934
rect 246022 246698 281786 246934
rect 282022 246698 317786 246934
rect 318022 246698 353786 246934
rect 354022 246698 389786 246934
rect 390022 246698 425786 246934
rect 426022 246698 461786 246934
rect 462022 246698 497786 246934
rect 498022 246698 533786 246934
rect 534022 246698 569786 246934
rect 570022 246698 592082 246934
rect 592318 246698 592500 246934
rect -8576 246676 592500 246698
rect -8576 246674 -7976 246676
rect 29604 246674 30204 246676
rect 65604 246674 66204 246676
rect 101604 246674 102204 246676
rect 137604 246674 138204 246676
rect 173604 246674 174204 246676
rect 209604 246674 210204 246676
rect 245604 246674 246204 246676
rect 281604 246674 282204 246676
rect 317604 246674 318204 246676
rect 353604 246674 354204 246676
rect 389604 246674 390204 246676
rect 425604 246674 426204 246676
rect 461604 246674 462204 246676
rect 497604 246674 498204 246676
rect 533604 246674 534204 246676
rect 569604 246674 570204 246676
rect 591900 246674 592500 246676
rect -6696 243676 -6096 243678
rect 26004 243676 26604 243678
rect 62004 243676 62604 243678
rect 98004 243676 98604 243678
rect 134004 243676 134604 243678
rect 170004 243676 170604 243678
rect 206004 243676 206604 243678
rect 242004 243676 242604 243678
rect 278004 243676 278604 243678
rect 314004 243676 314604 243678
rect 350004 243676 350604 243678
rect 386004 243676 386604 243678
rect 422004 243676 422604 243678
rect 458004 243676 458604 243678
rect 494004 243676 494604 243678
rect 530004 243676 530604 243678
rect 566004 243676 566604 243678
rect 590020 243676 590620 243678
rect -6696 243654 590620 243676
rect -6696 243418 -6514 243654
rect -6278 243418 26186 243654
rect 26422 243418 62186 243654
rect 62422 243418 98186 243654
rect 98422 243418 134186 243654
rect 134422 243418 170186 243654
rect 170422 243418 206186 243654
rect 206422 243418 242186 243654
rect 242422 243418 278186 243654
rect 278422 243418 314186 243654
rect 314422 243418 350186 243654
rect 350422 243418 386186 243654
rect 386422 243418 422186 243654
rect 422422 243418 458186 243654
rect 458422 243418 494186 243654
rect 494422 243418 530186 243654
rect 530422 243418 566186 243654
rect 566422 243418 590202 243654
rect 590438 243418 590620 243654
rect -6696 243334 590620 243418
rect -6696 243098 -6514 243334
rect -6278 243098 26186 243334
rect 26422 243098 62186 243334
rect 62422 243098 98186 243334
rect 98422 243098 134186 243334
rect 134422 243098 170186 243334
rect 170422 243098 206186 243334
rect 206422 243098 242186 243334
rect 242422 243098 278186 243334
rect 278422 243098 314186 243334
rect 314422 243098 350186 243334
rect 350422 243098 386186 243334
rect 386422 243098 422186 243334
rect 422422 243098 458186 243334
rect 458422 243098 494186 243334
rect 494422 243098 530186 243334
rect 530422 243098 566186 243334
rect 566422 243098 590202 243334
rect 590438 243098 590620 243334
rect -6696 243076 590620 243098
rect -6696 243074 -6096 243076
rect 26004 243074 26604 243076
rect 62004 243074 62604 243076
rect 98004 243074 98604 243076
rect 134004 243074 134604 243076
rect 170004 243074 170604 243076
rect 206004 243074 206604 243076
rect 242004 243074 242604 243076
rect 278004 243074 278604 243076
rect 314004 243074 314604 243076
rect 350004 243074 350604 243076
rect 386004 243074 386604 243076
rect 422004 243074 422604 243076
rect 458004 243074 458604 243076
rect 494004 243074 494604 243076
rect 530004 243074 530604 243076
rect 566004 243074 566604 243076
rect 590020 243074 590620 243076
rect -4816 240076 -4216 240078
rect 22404 240076 23004 240078
rect 58404 240076 59004 240078
rect 94404 240076 95004 240078
rect 130404 240076 131004 240078
rect 166404 240076 167004 240078
rect 202404 240076 203004 240078
rect 238404 240076 239004 240078
rect 274404 240076 275004 240078
rect 310404 240076 311004 240078
rect 346404 240076 347004 240078
rect 382404 240076 383004 240078
rect 418404 240076 419004 240078
rect 454404 240076 455004 240078
rect 490404 240076 491004 240078
rect 526404 240076 527004 240078
rect 562404 240076 563004 240078
rect 588140 240076 588740 240078
rect -4816 240054 588740 240076
rect -4816 239818 -4634 240054
rect -4398 239818 22586 240054
rect 22822 239818 58586 240054
rect 58822 239818 94586 240054
rect 94822 239818 130586 240054
rect 130822 239818 166586 240054
rect 166822 239818 202586 240054
rect 202822 239818 238586 240054
rect 238822 239818 274586 240054
rect 274822 239818 310586 240054
rect 310822 239818 346586 240054
rect 346822 239818 382586 240054
rect 382822 239818 418586 240054
rect 418822 239818 454586 240054
rect 454822 239818 490586 240054
rect 490822 239818 526586 240054
rect 526822 239818 562586 240054
rect 562822 239818 588322 240054
rect 588558 239818 588740 240054
rect -4816 239734 588740 239818
rect -4816 239498 -4634 239734
rect -4398 239498 22586 239734
rect 22822 239498 58586 239734
rect 58822 239498 94586 239734
rect 94822 239498 130586 239734
rect 130822 239498 166586 239734
rect 166822 239498 202586 239734
rect 202822 239498 238586 239734
rect 238822 239498 274586 239734
rect 274822 239498 310586 239734
rect 310822 239498 346586 239734
rect 346822 239498 382586 239734
rect 382822 239498 418586 239734
rect 418822 239498 454586 239734
rect 454822 239498 490586 239734
rect 490822 239498 526586 239734
rect 526822 239498 562586 239734
rect 562822 239498 588322 239734
rect 588558 239498 588740 239734
rect -4816 239476 588740 239498
rect -4816 239474 -4216 239476
rect 22404 239474 23004 239476
rect 58404 239474 59004 239476
rect 94404 239474 95004 239476
rect 130404 239474 131004 239476
rect 166404 239474 167004 239476
rect 202404 239474 203004 239476
rect 238404 239474 239004 239476
rect 274404 239474 275004 239476
rect 310404 239474 311004 239476
rect 346404 239474 347004 239476
rect 382404 239474 383004 239476
rect 418404 239474 419004 239476
rect 454404 239474 455004 239476
rect 490404 239474 491004 239476
rect 526404 239474 527004 239476
rect 562404 239474 563004 239476
rect 588140 239474 588740 239476
rect -2936 236476 -2336 236478
rect 18804 236476 19404 236478
rect 54804 236476 55404 236478
rect 90804 236476 91404 236478
rect 126804 236476 127404 236478
rect 162804 236476 163404 236478
rect 198804 236476 199404 236478
rect 234804 236476 235404 236478
rect 270804 236476 271404 236478
rect 306804 236476 307404 236478
rect 342804 236476 343404 236478
rect 378804 236476 379404 236478
rect 414804 236476 415404 236478
rect 450804 236476 451404 236478
rect 486804 236476 487404 236478
rect 522804 236476 523404 236478
rect 558804 236476 559404 236478
rect 586260 236476 586860 236478
rect -2936 236454 586860 236476
rect -2936 236218 -2754 236454
rect -2518 236218 18986 236454
rect 19222 236218 54986 236454
rect 55222 236218 90986 236454
rect 91222 236218 126986 236454
rect 127222 236218 162986 236454
rect 163222 236218 198986 236454
rect 199222 236218 234986 236454
rect 235222 236218 270986 236454
rect 271222 236218 306986 236454
rect 307222 236218 342986 236454
rect 343222 236218 378986 236454
rect 379222 236218 414986 236454
rect 415222 236218 450986 236454
rect 451222 236218 486986 236454
rect 487222 236218 522986 236454
rect 523222 236218 558986 236454
rect 559222 236218 586442 236454
rect 586678 236218 586860 236454
rect -2936 236134 586860 236218
rect -2936 235898 -2754 236134
rect -2518 235898 18986 236134
rect 19222 235898 54986 236134
rect 55222 235898 90986 236134
rect 91222 235898 126986 236134
rect 127222 235898 162986 236134
rect 163222 235898 198986 236134
rect 199222 235898 234986 236134
rect 235222 235898 270986 236134
rect 271222 235898 306986 236134
rect 307222 235898 342986 236134
rect 343222 235898 378986 236134
rect 379222 235898 414986 236134
rect 415222 235898 450986 236134
rect 451222 235898 486986 236134
rect 487222 235898 522986 236134
rect 523222 235898 558986 236134
rect 559222 235898 586442 236134
rect 586678 235898 586860 236134
rect -2936 235876 586860 235898
rect -2936 235874 -2336 235876
rect 18804 235874 19404 235876
rect 54804 235874 55404 235876
rect 90804 235874 91404 235876
rect 126804 235874 127404 235876
rect 162804 235874 163404 235876
rect 198804 235874 199404 235876
rect 234804 235874 235404 235876
rect 270804 235874 271404 235876
rect 306804 235874 307404 235876
rect 342804 235874 343404 235876
rect 378804 235874 379404 235876
rect 414804 235874 415404 235876
rect 450804 235874 451404 235876
rect 486804 235874 487404 235876
rect 522804 235874 523404 235876
rect 558804 235874 559404 235876
rect 586260 235874 586860 235876
rect -7636 229276 -7036 229278
rect 11604 229276 12204 229278
rect 47604 229276 48204 229278
rect 83604 229276 84204 229278
rect 119604 229276 120204 229278
rect 155604 229276 156204 229278
rect 191604 229276 192204 229278
rect 227604 229276 228204 229278
rect 263604 229276 264204 229278
rect 299604 229276 300204 229278
rect 335604 229276 336204 229278
rect 371604 229276 372204 229278
rect 407604 229276 408204 229278
rect 443604 229276 444204 229278
rect 479604 229276 480204 229278
rect 515604 229276 516204 229278
rect 551604 229276 552204 229278
rect 590960 229276 591560 229278
rect -8576 229254 592500 229276
rect -8576 229018 -7454 229254
rect -7218 229018 11786 229254
rect 12022 229018 47786 229254
rect 48022 229018 83786 229254
rect 84022 229018 119786 229254
rect 120022 229018 155786 229254
rect 156022 229018 191786 229254
rect 192022 229018 227786 229254
rect 228022 229018 263786 229254
rect 264022 229018 299786 229254
rect 300022 229018 335786 229254
rect 336022 229018 371786 229254
rect 372022 229018 407786 229254
rect 408022 229018 443786 229254
rect 444022 229018 479786 229254
rect 480022 229018 515786 229254
rect 516022 229018 551786 229254
rect 552022 229018 591142 229254
rect 591378 229018 592500 229254
rect -8576 228934 592500 229018
rect -8576 228698 -7454 228934
rect -7218 228698 11786 228934
rect 12022 228698 47786 228934
rect 48022 228698 83786 228934
rect 84022 228698 119786 228934
rect 120022 228698 155786 228934
rect 156022 228698 191786 228934
rect 192022 228698 227786 228934
rect 228022 228698 263786 228934
rect 264022 228698 299786 228934
rect 300022 228698 335786 228934
rect 336022 228698 371786 228934
rect 372022 228698 407786 228934
rect 408022 228698 443786 228934
rect 444022 228698 479786 228934
rect 480022 228698 515786 228934
rect 516022 228698 551786 228934
rect 552022 228698 591142 228934
rect 591378 228698 592500 228934
rect -8576 228676 592500 228698
rect -7636 228674 -7036 228676
rect 11604 228674 12204 228676
rect 47604 228674 48204 228676
rect 83604 228674 84204 228676
rect 119604 228674 120204 228676
rect 155604 228674 156204 228676
rect 191604 228674 192204 228676
rect 227604 228674 228204 228676
rect 263604 228674 264204 228676
rect 299604 228674 300204 228676
rect 335604 228674 336204 228676
rect 371604 228674 372204 228676
rect 407604 228674 408204 228676
rect 443604 228674 444204 228676
rect 479604 228674 480204 228676
rect 515604 228674 516204 228676
rect 551604 228674 552204 228676
rect 590960 228674 591560 228676
rect -5756 225676 -5156 225678
rect 8004 225676 8604 225678
rect 44004 225676 44604 225678
rect 80004 225676 80604 225678
rect 116004 225676 116604 225678
rect 152004 225676 152604 225678
rect 188004 225676 188604 225678
rect 224004 225676 224604 225678
rect 260004 225676 260604 225678
rect 296004 225676 296604 225678
rect 332004 225676 332604 225678
rect 368004 225676 368604 225678
rect 404004 225676 404604 225678
rect 440004 225676 440604 225678
rect 476004 225676 476604 225678
rect 512004 225676 512604 225678
rect 548004 225676 548604 225678
rect 589080 225676 589680 225678
rect -6696 225654 590620 225676
rect -6696 225418 -5574 225654
rect -5338 225418 8186 225654
rect 8422 225418 44186 225654
rect 44422 225418 80186 225654
rect 80422 225418 116186 225654
rect 116422 225418 152186 225654
rect 152422 225418 188186 225654
rect 188422 225418 224186 225654
rect 224422 225418 260186 225654
rect 260422 225418 296186 225654
rect 296422 225418 332186 225654
rect 332422 225418 368186 225654
rect 368422 225418 404186 225654
rect 404422 225418 440186 225654
rect 440422 225418 476186 225654
rect 476422 225418 512186 225654
rect 512422 225418 548186 225654
rect 548422 225418 589262 225654
rect 589498 225418 590620 225654
rect -6696 225334 590620 225418
rect -6696 225098 -5574 225334
rect -5338 225098 8186 225334
rect 8422 225098 44186 225334
rect 44422 225098 80186 225334
rect 80422 225098 116186 225334
rect 116422 225098 152186 225334
rect 152422 225098 188186 225334
rect 188422 225098 224186 225334
rect 224422 225098 260186 225334
rect 260422 225098 296186 225334
rect 296422 225098 332186 225334
rect 332422 225098 368186 225334
rect 368422 225098 404186 225334
rect 404422 225098 440186 225334
rect 440422 225098 476186 225334
rect 476422 225098 512186 225334
rect 512422 225098 548186 225334
rect 548422 225098 589262 225334
rect 589498 225098 590620 225334
rect -6696 225076 590620 225098
rect -5756 225074 -5156 225076
rect 8004 225074 8604 225076
rect 44004 225074 44604 225076
rect 80004 225074 80604 225076
rect 116004 225074 116604 225076
rect 152004 225074 152604 225076
rect 188004 225074 188604 225076
rect 224004 225074 224604 225076
rect 260004 225074 260604 225076
rect 296004 225074 296604 225076
rect 332004 225074 332604 225076
rect 368004 225074 368604 225076
rect 404004 225074 404604 225076
rect 440004 225074 440604 225076
rect 476004 225074 476604 225076
rect 512004 225074 512604 225076
rect 548004 225074 548604 225076
rect 589080 225074 589680 225076
rect -3876 222076 -3276 222078
rect 4404 222076 5004 222078
rect 40404 222076 41004 222078
rect 76404 222076 77004 222078
rect 112404 222076 113004 222078
rect 148404 222076 149004 222078
rect 184404 222076 185004 222078
rect 220404 222076 221004 222078
rect 256404 222076 257004 222078
rect 292404 222076 293004 222078
rect 328404 222076 329004 222078
rect 364404 222076 365004 222078
rect 400404 222076 401004 222078
rect 436404 222076 437004 222078
rect 472404 222076 473004 222078
rect 508404 222076 509004 222078
rect 544404 222076 545004 222078
rect 580404 222076 581004 222078
rect 587200 222076 587800 222078
rect -4816 222054 588740 222076
rect -4816 221818 -3694 222054
rect -3458 221818 4586 222054
rect 4822 221818 40586 222054
rect 40822 221818 76586 222054
rect 76822 221818 112586 222054
rect 112822 221818 148586 222054
rect 148822 221818 184586 222054
rect 184822 221818 220586 222054
rect 220822 221818 256586 222054
rect 256822 221818 292586 222054
rect 292822 221818 328586 222054
rect 328822 221818 364586 222054
rect 364822 221818 400586 222054
rect 400822 221818 436586 222054
rect 436822 221818 472586 222054
rect 472822 221818 508586 222054
rect 508822 221818 544586 222054
rect 544822 221818 580586 222054
rect 580822 221818 587382 222054
rect 587618 221818 588740 222054
rect -4816 221734 588740 221818
rect -4816 221498 -3694 221734
rect -3458 221498 4586 221734
rect 4822 221498 40586 221734
rect 40822 221498 76586 221734
rect 76822 221498 112586 221734
rect 112822 221498 148586 221734
rect 148822 221498 184586 221734
rect 184822 221498 220586 221734
rect 220822 221498 256586 221734
rect 256822 221498 292586 221734
rect 292822 221498 328586 221734
rect 328822 221498 364586 221734
rect 364822 221498 400586 221734
rect 400822 221498 436586 221734
rect 436822 221498 472586 221734
rect 472822 221498 508586 221734
rect 508822 221498 544586 221734
rect 544822 221498 580586 221734
rect 580822 221498 587382 221734
rect 587618 221498 588740 221734
rect -4816 221476 588740 221498
rect -3876 221474 -3276 221476
rect 4404 221474 5004 221476
rect 40404 221474 41004 221476
rect 76404 221474 77004 221476
rect 112404 221474 113004 221476
rect 148404 221474 149004 221476
rect 184404 221474 185004 221476
rect 220404 221474 221004 221476
rect 256404 221474 257004 221476
rect 292404 221474 293004 221476
rect 328404 221474 329004 221476
rect 364404 221474 365004 221476
rect 400404 221474 401004 221476
rect 436404 221474 437004 221476
rect 472404 221474 473004 221476
rect 508404 221474 509004 221476
rect 544404 221474 545004 221476
rect 580404 221474 581004 221476
rect 587200 221474 587800 221476
rect -1996 218476 -1396 218478
rect 804 218476 1404 218478
rect 36804 218476 37404 218478
rect 72804 218476 73404 218478
rect 108804 218476 109404 218478
rect 144804 218476 145404 218478
rect 180804 218476 181404 218478
rect 216804 218476 217404 218478
rect 252804 218476 253404 218478
rect 288804 218476 289404 218478
rect 324804 218476 325404 218478
rect 360804 218476 361404 218478
rect 396804 218476 397404 218478
rect 432804 218476 433404 218478
rect 468804 218476 469404 218478
rect 504804 218476 505404 218478
rect 540804 218476 541404 218478
rect 576804 218476 577404 218478
rect 585320 218476 585920 218478
rect -2936 218454 586860 218476
rect -2936 218218 -1814 218454
rect -1578 218218 986 218454
rect 1222 218218 36986 218454
rect 37222 218218 72986 218454
rect 73222 218218 108986 218454
rect 109222 218218 144986 218454
rect 145222 218218 180986 218454
rect 181222 218218 216986 218454
rect 217222 218218 252986 218454
rect 253222 218218 288986 218454
rect 289222 218218 324986 218454
rect 325222 218218 360986 218454
rect 361222 218218 396986 218454
rect 397222 218218 432986 218454
rect 433222 218218 468986 218454
rect 469222 218218 504986 218454
rect 505222 218218 540986 218454
rect 541222 218218 576986 218454
rect 577222 218218 585502 218454
rect 585738 218218 586860 218454
rect -2936 218134 586860 218218
rect -2936 217898 -1814 218134
rect -1578 217898 986 218134
rect 1222 217898 36986 218134
rect 37222 217898 72986 218134
rect 73222 217898 108986 218134
rect 109222 217898 144986 218134
rect 145222 217898 180986 218134
rect 181222 217898 216986 218134
rect 217222 217898 252986 218134
rect 253222 217898 288986 218134
rect 289222 217898 324986 218134
rect 325222 217898 360986 218134
rect 361222 217898 396986 218134
rect 397222 217898 432986 218134
rect 433222 217898 468986 218134
rect 469222 217898 504986 218134
rect 505222 217898 540986 218134
rect 541222 217898 576986 218134
rect 577222 217898 585502 218134
rect 585738 217898 586860 218134
rect -2936 217876 586860 217898
rect -1996 217874 -1396 217876
rect 804 217874 1404 217876
rect 36804 217874 37404 217876
rect 72804 217874 73404 217876
rect 108804 217874 109404 217876
rect 144804 217874 145404 217876
rect 180804 217874 181404 217876
rect 216804 217874 217404 217876
rect 252804 217874 253404 217876
rect 288804 217874 289404 217876
rect 324804 217874 325404 217876
rect 360804 217874 361404 217876
rect 396804 217874 397404 217876
rect 432804 217874 433404 217876
rect 468804 217874 469404 217876
rect 504804 217874 505404 217876
rect 540804 217874 541404 217876
rect 576804 217874 577404 217876
rect 585320 217874 585920 217876
rect -8576 211276 -7976 211278
rect 29604 211276 30204 211278
rect 65604 211276 66204 211278
rect 101604 211276 102204 211278
rect 137604 211276 138204 211278
rect 173604 211276 174204 211278
rect 209604 211276 210204 211278
rect 245604 211276 246204 211278
rect 281604 211276 282204 211278
rect 317604 211276 318204 211278
rect 353604 211276 354204 211278
rect 389604 211276 390204 211278
rect 425604 211276 426204 211278
rect 461604 211276 462204 211278
rect 497604 211276 498204 211278
rect 533604 211276 534204 211278
rect 569604 211276 570204 211278
rect 591900 211276 592500 211278
rect -8576 211254 592500 211276
rect -8576 211018 -8394 211254
rect -8158 211018 29786 211254
rect 30022 211018 65786 211254
rect 66022 211018 101786 211254
rect 102022 211018 137786 211254
rect 138022 211018 173786 211254
rect 174022 211018 209786 211254
rect 210022 211018 245786 211254
rect 246022 211018 281786 211254
rect 282022 211018 317786 211254
rect 318022 211018 353786 211254
rect 354022 211018 389786 211254
rect 390022 211018 425786 211254
rect 426022 211018 461786 211254
rect 462022 211018 497786 211254
rect 498022 211018 533786 211254
rect 534022 211018 569786 211254
rect 570022 211018 592082 211254
rect 592318 211018 592500 211254
rect -8576 210934 592500 211018
rect -8576 210698 -8394 210934
rect -8158 210698 29786 210934
rect 30022 210698 65786 210934
rect 66022 210698 101786 210934
rect 102022 210698 137786 210934
rect 138022 210698 173786 210934
rect 174022 210698 209786 210934
rect 210022 210698 245786 210934
rect 246022 210698 281786 210934
rect 282022 210698 317786 210934
rect 318022 210698 353786 210934
rect 354022 210698 389786 210934
rect 390022 210698 425786 210934
rect 426022 210698 461786 210934
rect 462022 210698 497786 210934
rect 498022 210698 533786 210934
rect 534022 210698 569786 210934
rect 570022 210698 592082 210934
rect 592318 210698 592500 210934
rect -8576 210676 592500 210698
rect -8576 210674 -7976 210676
rect 29604 210674 30204 210676
rect 65604 210674 66204 210676
rect 101604 210674 102204 210676
rect 137604 210674 138204 210676
rect 173604 210674 174204 210676
rect 209604 210674 210204 210676
rect 245604 210674 246204 210676
rect 281604 210674 282204 210676
rect 317604 210674 318204 210676
rect 353604 210674 354204 210676
rect 389604 210674 390204 210676
rect 425604 210674 426204 210676
rect 461604 210674 462204 210676
rect 497604 210674 498204 210676
rect 533604 210674 534204 210676
rect 569604 210674 570204 210676
rect 591900 210674 592500 210676
rect -6696 207676 -6096 207678
rect 26004 207676 26604 207678
rect 62004 207676 62604 207678
rect 98004 207676 98604 207678
rect 134004 207676 134604 207678
rect 170004 207676 170604 207678
rect 206004 207676 206604 207678
rect 242004 207676 242604 207678
rect 278004 207676 278604 207678
rect 314004 207676 314604 207678
rect 350004 207676 350604 207678
rect 386004 207676 386604 207678
rect 422004 207676 422604 207678
rect 458004 207676 458604 207678
rect 494004 207676 494604 207678
rect 530004 207676 530604 207678
rect 566004 207676 566604 207678
rect 590020 207676 590620 207678
rect -6696 207654 590620 207676
rect -6696 207418 -6514 207654
rect -6278 207418 26186 207654
rect 26422 207418 62186 207654
rect 62422 207418 98186 207654
rect 98422 207418 134186 207654
rect 134422 207418 170186 207654
rect 170422 207418 206186 207654
rect 206422 207418 242186 207654
rect 242422 207418 278186 207654
rect 278422 207418 314186 207654
rect 314422 207418 350186 207654
rect 350422 207418 386186 207654
rect 386422 207418 422186 207654
rect 422422 207418 458186 207654
rect 458422 207418 494186 207654
rect 494422 207418 530186 207654
rect 530422 207418 566186 207654
rect 566422 207418 590202 207654
rect 590438 207418 590620 207654
rect -6696 207334 590620 207418
rect -6696 207098 -6514 207334
rect -6278 207098 26186 207334
rect 26422 207098 62186 207334
rect 62422 207098 98186 207334
rect 98422 207098 134186 207334
rect 134422 207098 170186 207334
rect 170422 207098 206186 207334
rect 206422 207098 242186 207334
rect 242422 207098 278186 207334
rect 278422 207098 314186 207334
rect 314422 207098 350186 207334
rect 350422 207098 386186 207334
rect 386422 207098 422186 207334
rect 422422 207098 458186 207334
rect 458422 207098 494186 207334
rect 494422 207098 530186 207334
rect 530422 207098 566186 207334
rect 566422 207098 590202 207334
rect 590438 207098 590620 207334
rect -6696 207076 590620 207098
rect -6696 207074 -6096 207076
rect 26004 207074 26604 207076
rect 62004 207074 62604 207076
rect 98004 207074 98604 207076
rect 134004 207074 134604 207076
rect 170004 207074 170604 207076
rect 206004 207074 206604 207076
rect 242004 207074 242604 207076
rect 278004 207074 278604 207076
rect 314004 207074 314604 207076
rect 350004 207074 350604 207076
rect 386004 207074 386604 207076
rect 422004 207074 422604 207076
rect 458004 207074 458604 207076
rect 494004 207074 494604 207076
rect 530004 207074 530604 207076
rect 566004 207074 566604 207076
rect 590020 207074 590620 207076
rect -4816 204076 -4216 204078
rect 22404 204076 23004 204078
rect 58404 204076 59004 204078
rect 94404 204076 95004 204078
rect 130404 204076 131004 204078
rect 166404 204076 167004 204078
rect 202404 204076 203004 204078
rect 238404 204076 239004 204078
rect 274404 204076 275004 204078
rect 310404 204076 311004 204078
rect 346404 204076 347004 204078
rect 382404 204076 383004 204078
rect 418404 204076 419004 204078
rect 454404 204076 455004 204078
rect 490404 204076 491004 204078
rect 526404 204076 527004 204078
rect 562404 204076 563004 204078
rect 588140 204076 588740 204078
rect -4816 204054 588740 204076
rect -4816 203818 -4634 204054
rect -4398 203818 22586 204054
rect 22822 203818 58586 204054
rect 58822 203818 94586 204054
rect 94822 203818 130586 204054
rect 130822 203818 166586 204054
rect 166822 203818 202586 204054
rect 202822 203818 238586 204054
rect 238822 203818 274586 204054
rect 274822 203818 310586 204054
rect 310822 203818 346586 204054
rect 346822 203818 382586 204054
rect 382822 203818 418586 204054
rect 418822 203818 454586 204054
rect 454822 203818 490586 204054
rect 490822 203818 526586 204054
rect 526822 203818 562586 204054
rect 562822 203818 588322 204054
rect 588558 203818 588740 204054
rect -4816 203734 588740 203818
rect -4816 203498 -4634 203734
rect -4398 203498 22586 203734
rect 22822 203498 58586 203734
rect 58822 203498 94586 203734
rect 94822 203498 130586 203734
rect 130822 203498 166586 203734
rect 166822 203498 202586 203734
rect 202822 203498 238586 203734
rect 238822 203498 274586 203734
rect 274822 203498 310586 203734
rect 310822 203498 346586 203734
rect 346822 203498 382586 203734
rect 382822 203498 418586 203734
rect 418822 203498 454586 203734
rect 454822 203498 490586 203734
rect 490822 203498 526586 203734
rect 526822 203498 562586 203734
rect 562822 203498 588322 203734
rect 588558 203498 588740 203734
rect -4816 203476 588740 203498
rect -4816 203474 -4216 203476
rect 22404 203474 23004 203476
rect 58404 203474 59004 203476
rect 94404 203474 95004 203476
rect 130404 203474 131004 203476
rect 166404 203474 167004 203476
rect 202404 203474 203004 203476
rect 238404 203474 239004 203476
rect 274404 203474 275004 203476
rect 310404 203474 311004 203476
rect 346404 203474 347004 203476
rect 382404 203474 383004 203476
rect 418404 203474 419004 203476
rect 454404 203474 455004 203476
rect 490404 203474 491004 203476
rect 526404 203474 527004 203476
rect 562404 203474 563004 203476
rect 588140 203474 588740 203476
rect -2936 200476 -2336 200478
rect 18804 200476 19404 200478
rect 54804 200476 55404 200478
rect 90804 200476 91404 200478
rect 126804 200476 127404 200478
rect 162804 200476 163404 200478
rect 198804 200476 199404 200478
rect 234804 200476 235404 200478
rect 270804 200476 271404 200478
rect 306804 200476 307404 200478
rect 342804 200476 343404 200478
rect 378804 200476 379404 200478
rect 414804 200476 415404 200478
rect 450804 200476 451404 200478
rect 486804 200476 487404 200478
rect 522804 200476 523404 200478
rect 558804 200476 559404 200478
rect 586260 200476 586860 200478
rect -2936 200454 586860 200476
rect -2936 200218 -2754 200454
rect -2518 200218 18986 200454
rect 19222 200218 54986 200454
rect 55222 200218 90986 200454
rect 91222 200218 126986 200454
rect 127222 200218 162986 200454
rect 163222 200218 198986 200454
rect 199222 200218 234986 200454
rect 235222 200218 270986 200454
rect 271222 200218 306986 200454
rect 307222 200218 342986 200454
rect 343222 200218 378986 200454
rect 379222 200218 414986 200454
rect 415222 200218 450986 200454
rect 451222 200218 486986 200454
rect 487222 200218 522986 200454
rect 523222 200218 558986 200454
rect 559222 200218 586442 200454
rect 586678 200218 586860 200454
rect -2936 200134 586860 200218
rect -2936 199898 -2754 200134
rect -2518 199898 18986 200134
rect 19222 199898 54986 200134
rect 55222 199898 90986 200134
rect 91222 199898 126986 200134
rect 127222 199898 162986 200134
rect 163222 199898 198986 200134
rect 199222 199898 234986 200134
rect 235222 199898 270986 200134
rect 271222 199898 306986 200134
rect 307222 199898 342986 200134
rect 343222 199898 378986 200134
rect 379222 199898 414986 200134
rect 415222 199898 450986 200134
rect 451222 199898 486986 200134
rect 487222 199898 522986 200134
rect 523222 199898 558986 200134
rect 559222 199898 586442 200134
rect 586678 199898 586860 200134
rect -2936 199876 586860 199898
rect -2936 199874 -2336 199876
rect 18804 199874 19404 199876
rect 54804 199874 55404 199876
rect 90804 199874 91404 199876
rect 126804 199874 127404 199876
rect 162804 199874 163404 199876
rect 198804 199874 199404 199876
rect 234804 199874 235404 199876
rect 270804 199874 271404 199876
rect 306804 199874 307404 199876
rect 342804 199874 343404 199876
rect 378804 199874 379404 199876
rect 414804 199874 415404 199876
rect 450804 199874 451404 199876
rect 486804 199874 487404 199876
rect 522804 199874 523404 199876
rect 558804 199874 559404 199876
rect 586260 199874 586860 199876
rect -7636 193276 -7036 193278
rect 11604 193276 12204 193278
rect 47604 193276 48204 193278
rect 83604 193276 84204 193278
rect 119604 193276 120204 193278
rect 155604 193276 156204 193278
rect 191604 193276 192204 193278
rect 227604 193276 228204 193278
rect 263604 193276 264204 193278
rect 299604 193276 300204 193278
rect 335604 193276 336204 193278
rect 371604 193276 372204 193278
rect 407604 193276 408204 193278
rect 443604 193276 444204 193278
rect 479604 193276 480204 193278
rect 515604 193276 516204 193278
rect 551604 193276 552204 193278
rect 590960 193276 591560 193278
rect -8576 193254 592500 193276
rect -8576 193018 -7454 193254
rect -7218 193018 11786 193254
rect 12022 193018 47786 193254
rect 48022 193018 83786 193254
rect 84022 193018 119786 193254
rect 120022 193018 155786 193254
rect 156022 193018 191786 193254
rect 192022 193018 227786 193254
rect 228022 193018 263786 193254
rect 264022 193018 299786 193254
rect 300022 193018 335786 193254
rect 336022 193018 371786 193254
rect 372022 193018 407786 193254
rect 408022 193018 443786 193254
rect 444022 193018 479786 193254
rect 480022 193018 515786 193254
rect 516022 193018 551786 193254
rect 552022 193018 591142 193254
rect 591378 193018 592500 193254
rect -8576 192934 592500 193018
rect -8576 192698 -7454 192934
rect -7218 192698 11786 192934
rect 12022 192698 47786 192934
rect 48022 192698 83786 192934
rect 84022 192698 119786 192934
rect 120022 192698 155786 192934
rect 156022 192698 191786 192934
rect 192022 192698 227786 192934
rect 228022 192698 263786 192934
rect 264022 192698 299786 192934
rect 300022 192698 335786 192934
rect 336022 192698 371786 192934
rect 372022 192698 407786 192934
rect 408022 192698 443786 192934
rect 444022 192698 479786 192934
rect 480022 192698 515786 192934
rect 516022 192698 551786 192934
rect 552022 192698 591142 192934
rect 591378 192698 592500 192934
rect -8576 192676 592500 192698
rect -7636 192674 -7036 192676
rect 11604 192674 12204 192676
rect 47604 192674 48204 192676
rect 83604 192674 84204 192676
rect 119604 192674 120204 192676
rect 155604 192674 156204 192676
rect 191604 192674 192204 192676
rect 227604 192674 228204 192676
rect 263604 192674 264204 192676
rect 299604 192674 300204 192676
rect 335604 192674 336204 192676
rect 371604 192674 372204 192676
rect 407604 192674 408204 192676
rect 443604 192674 444204 192676
rect 479604 192674 480204 192676
rect 515604 192674 516204 192676
rect 551604 192674 552204 192676
rect 590960 192674 591560 192676
rect -5756 189676 -5156 189678
rect 8004 189676 8604 189678
rect 44004 189676 44604 189678
rect 80004 189676 80604 189678
rect 116004 189676 116604 189678
rect 152004 189676 152604 189678
rect 188004 189676 188604 189678
rect 224004 189676 224604 189678
rect 260004 189676 260604 189678
rect 296004 189676 296604 189678
rect 332004 189676 332604 189678
rect 368004 189676 368604 189678
rect 404004 189676 404604 189678
rect 440004 189676 440604 189678
rect 476004 189676 476604 189678
rect 512004 189676 512604 189678
rect 548004 189676 548604 189678
rect 589080 189676 589680 189678
rect -6696 189654 590620 189676
rect -6696 189418 -5574 189654
rect -5338 189418 8186 189654
rect 8422 189418 44186 189654
rect 44422 189418 80186 189654
rect 80422 189418 116186 189654
rect 116422 189418 152186 189654
rect 152422 189418 188186 189654
rect 188422 189418 224186 189654
rect 224422 189418 260186 189654
rect 260422 189418 296186 189654
rect 296422 189418 332186 189654
rect 332422 189418 368186 189654
rect 368422 189418 404186 189654
rect 404422 189418 440186 189654
rect 440422 189418 476186 189654
rect 476422 189418 512186 189654
rect 512422 189418 548186 189654
rect 548422 189418 589262 189654
rect 589498 189418 590620 189654
rect -6696 189334 590620 189418
rect -6696 189098 -5574 189334
rect -5338 189098 8186 189334
rect 8422 189098 44186 189334
rect 44422 189098 80186 189334
rect 80422 189098 116186 189334
rect 116422 189098 152186 189334
rect 152422 189098 188186 189334
rect 188422 189098 224186 189334
rect 224422 189098 260186 189334
rect 260422 189098 296186 189334
rect 296422 189098 332186 189334
rect 332422 189098 368186 189334
rect 368422 189098 404186 189334
rect 404422 189098 440186 189334
rect 440422 189098 476186 189334
rect 476422 189098 512186 189334
rect 512422 189098 548186 189334
rect 548422 189098 589262 189334
rect 589498 189098 590620 189334
rect -6696 189076 590620 189098
rect -5756 189074 -5156 189076
rect 8004 189074 8604 189076
rect 44004 189074 44604 189076
rect 80004 189074 80604 189076
rect 116004 189074 116604 189076
rect 152004 189074 152604 189076
rect 188004 189074 188604 189076
rect 224004 189074 224604 189076
rect 260004 189074 260604 189076
rect 296004 189074 296604 189076
rect 332004 189074 332604 189076
rect 368004 189074 368604 189076
rect 404004 189074 404604 189076
rect 440004 189074 440604 189076
rect 476004 189074 476604 189076
rect 512004 189074 512604 189076
rect 548004 189074 548604 189076
rect 589080 189074 589680 189076
rect -3876 186076 -3276 186078
rect 4404 186076 5004 186078
rect 40404 186076 41004 186078
rect 76404 186076 77004 186078
rect 112404 186076 113004 186078
rect 148404 186076 149004 186078
rect 184404 186076 185004 186078
rect 220404 186076 221004 186078
rect 256404 186076 257004 186078
rect 292404 186076 293004 186078
rect 328404 186076 329004 186078
rect 364404 186076 365004 186078
rect 400404 186076 401004 186078
rect 436404 186076 437004 186078
rect 472404 186076 473004 186078
rect 508404 186076 509004 186078
rect 544404 186076 545004 186078
rect 580404 186076 581004 186078
rect 587200 186076 587800 186078
rect -4816 186054 588740 186076
rect -4816 185818 -3694 186054
rect -3458 185818 4586 186054
rect 4822 185818 40586 186054
rect 40822 185818 76586 186054
rect 76822 185818 112586 186054
rect 112822 185818 148586 186054
rect 148822 185818 184586 186054
rect 184822 185818 220586 186054
rect 220822 185818 256586 186054
rect 256822 185818 292586 186054
rect 292822 185818 328586 186054
rect 328822 185818 364586 186054
rect 364822 185818 400586 186054
rect 400822 185818 436586 186054
rect 436822 185818 472586 186054
rect 472822 185818 508586 186054
rect 508822 185818 544586 186054
rect 544822 185818 580586 186054
rect 580822 185818 587382 186054
rect 587618 185818 588740 186054
rect -4816 185734 588740 185818
rect -4816 185498 -3694 185734
rect -3458 185498 4586 185734
rect 4822 185498 40586 185734
rect 40822 185498 76586 185734
rect 76822 185498 112586 185734
rect 112822 185498 148586 185734
rect 148822 185498 184586 185734
rect 184822 185498 220586 185734
rect 220822 185498 256586 185734
rect 256822 185498 292586 185734
rect 292822 185498 328586 185734
rect 328822 185498 364586 185734
rect 364822 185498 400586 185734
rect 400822 185498 436586 185734
rect 436822 185498 472586 185734
rect 472822 185498 508586 185734
rect 508822 185498 544586 185734
rect 544822 185498 580586 185734
rect 580822 185498 587382 185734
rect 587618 185498 588740 185734
rect -4816 185476 588740 185498
rect -3876 185474 -3276 185476
rect 4404 185474 5004 185476
rect 40404 185474 41004 185476
rect 76404 185474 77004 185476
rect 112404 185474 113004 185476
rect 148404 185474 149004 185476
rect 184404 185474 185004 185476
rect 220404 185474 221004 185476
rect 256404 185474 257004 185476
rect 292404 185474 293004 185476
rect 328404 185474 329004 185476
rect 364404 185474 365004 185476
rect 400404 185474 401004 185476
rect 436404 185474 437004 185476
rect 472404 185474 473004 185476
rect 508404 185474 509004 185476
rect 544404 185474 545004 185476
rect 580404 185474 581004 185476
rect 587200 185474 587800 185476
rect -1996 182476 -1396 182478
rect 804 182476 1404 182478
rect 36804 182476 37404 182478
rect 72804 182476 73404 182478
rect 108804 182476 109404 182478
rect 144804 182476 145404 182478
rect 180804 182476 181404 182478
rect 216804 182476 217404 182478
rect 252804 182476 253404 182478
rect 288804 182476 289404 182478
rect 324804 182476 325404 182478
rect 360804 182476 361404 182478
rect 396804 182476 397404 182478
rect 432804 182476 433404 182478
rect 468804 182476 469404 182478
rect 504804 182476 505404 182478
rect 540804 182476 541404 182478
rect 576804 182476 577404 182478
rect 585320 182476 585920 182478
rect -2936 182454 586860 182476
rect -2936 182218 -1814 182454
rect -1578 182218 986 182454
rect 1222 182218 36986 182454
rect 37222 182218 72986 182454
rect 73222 182218 108986 182454
rect 109222 182218 144986 182454
rect 145222 182218 180986 182454
rect 181222 182218 216986 182454
rect 217222 182218 252986 182454
rect 253222 182218 288986 182454
rect 289222 182218 324986 182454
rect 325222 182218 360986 182454
rect 361222 182218 396986 182454
rect 397222 182218 432986 182454
rect 433222 182218 468986 182454
rect 469222 182218 504986 182454
rect 505222 182218 540986 182454
rect 541222 182218 576986 182454
rect 577222 182218 585502 182454
rect 585738 182218 586860 182454
rect -2936 182134 586860 182218
rect -2936 181898 -1814 182134
rect -1578 181898 986 182134
rect 1222 181898 36986 182134
rect 37222 181898 72986 182134
rect 73222 181898 108986 182134
rect 109222 181898 144986 182134
rect 145222 181898 180986 182134
rect 181222 181898 216986 182134
rect 217222 181898 252986 182134
rect 253222 181898 288986 182134
rect 289222 181898 324986 182134
rect 325222 181898 360986 182134
rect 361222 181898 396986 182134
rect 397222 181898 432986 182134
rect 433222 181898 468986 182134
rect 469222 181898 504986 182134
rect 505222 181898 540986 182134
rect 541222 181898 576986 182134
rect 577222 181898 585502 182134
rect 585738 181898 586860 182134
rect -2936 181876 586860 181898
rect -1996 181874 -1396 181876
rect 804 181874 1404 181876
rect 36804 181874 37404 181876
rect 72804 181874 73404 181876
rect 108804 181874 109404 181876
rect 144804 181874 145404 181876
rect 180804 181874 181404 181876
rect 216804 181874 217404 181876
rect 252804 181874 253404 181876
rect 288804 181874 289404 181876
rect 324804 181874 325404 181876
rect 360804 181874 361404 181876
rect 396804 181874 397404 181876
rect 432804 181874 433404 181876
rect 468804 181874 469404 181876
rect 504804 181874 505404 181876
rect 540804 181874 541404 181876
rect 576804 181874 577404 181876
rect 585320 181874 585920 181876
rect -8576 175276 -7976 175278
rect 29604 175276 30204 175278
rect 65604 175276 66204 175278
rect 101604 175276 102204 175278
rect 137604 175276 138204 175278
rect 173604 175276 174204 175278
rect 209604 175276 210204 175278
rect 245604 175276 246204 175278
rect 281604 175276 282204 175278
rect 317604 175276 318204 175278
rect 353604 175276 354204 175278
rect 389604 175276 390204 175278
rect 425604 175276 426204 175278
rect 461604 175276 462204 175278
rect 497604 175276 498204 175278
rect 533604 175276 534204 175278
rect 569604 175276 570204 175278
rect 591900 175276 592500 175278
rect -8576 175254 592500 175276
rect -8576 175018 -8394 175254
rect -8158 175018 29786 175254
rect 30022 175018 65786 175254
rect 66022 175018 101786 175254
rect 102022 175018 137786 175254
rect 138022 175018 173786 175254
rect 174022 175018 209786 175254
rect 210022 175018 245786 175254
rect 246022 175018 281786 175254
rect 282022 175018 317786 175254
rect 318022 175018 353786 175254
rect 354022 175018 389786 175254
rect 390022 175018 425786 175254
rect 426022 175018 461786 175254
rect 462022 175018 497786 175254
rect 498022 175018 533786 175254
rect 534022 175018 569786 175254
rect 570022 175018 592082 175254
rect 592318 175018 592500 175254
rect -8576 174934 592500 175018
rect -8576 174698 -8394 174934
rect -8158 174698 29786 174934
rect 30022 174698 65786 174934
rect 66022 174698 101786 174934
rect 102022 174698 137786 174934
rect 138022 174698 173786 174934
rect 174022 174698 209786 174934
rect 210022 174698 245786 174934
rect 246022 174698 281786 174934
rect 282022 174698 317786 174934
rect 318022 174698 353786 174934
rect 354022 174698 389786 174934
rect 390022 174698 425786 174934
rect 426022 174698 461786 174934
rect 462022 174698 497786 174934
rect 498022 174698 533786 174934
rect 534022 174698 569786 174934
rect 570022 174698 592082 174934
rect 592318 174698 592500 174934
rect -8576 174676 592500 174698
rect -8576 174674 -7976 174676
rect 29604 174674 30204 174676
rect 65604 174674 66204 174676
rect 101604 174674 102204 174676
rect 137604 174674 138204 174676
rect 173604 174674 174204 174676
rect 209604 174674 210204 174676
rect 245604 174674 246204 174676
rect 281604 174674 282204 174676
rect 317604 174674 318204 174676
rect 353604 174674 354204 174676
rect 389604 174674 390204 174676
rect 425604 174674 426204 174676
rect 461604 174674 462204 174676
rect 497604 174674 498204 174676
rect 533604 174674 534204 174676
rect 569604 174674 570204 174676
rect 591900 174674 592500 174676
rect -6696 171676 -6096 171678
rect 26004 171676 26604 171678
rect 62004 171676 62604 171678
rect 98004 171676 98604 171678
rect 134004 171676 134604 171678
rect 170004 171676 170604 171678
rect 206004 171676 206604 171678
rect 242004 171676 242604 171678
rect 278004 171676 278604 171678
rect 314004 171676 314604 171678
rect 350004 171676 350604 171678
rect 386004 171676 386604 171678
rect 422004 171676 422604 171678
rect 458004 171676 458604 171678
rect 494004 171676 494604 171678
rect 530004 171676 530604 171678
rect 566004 171676 566604 171678
rect 590020 171676 590620 171678
rect -6696 171654 590620 171676
rect -6696 171418 -6514 171654
rect -6278 171418 26186 171654
rect 26422 171418 62186 171654
rect 62422 171418 98186 171654
rect 98422 171418 134186 171654
rect 134422 171418 170186 171654
rect 170422 171418 206186 171654
rect 206422 171418 242186 171654
rect 242422 171418 278186 171654
rect 278422 171418 314186 171654
rect 314422 171418 350186 171654
rect 350422 171418 386186 171654
rect 386422 171418 422186 171654
rect 422422 171418 458186 171654
rect 458422 171418 494186 171654
rect 494422 171418 530186 171654
rect 530422 171418 566186 171654
rect 566422 171418 590202 171654
rect 590438 171418 590620 171654
rect -6696 171334 590620 171418
rect -6696 171098 -6514 171334
rect -6278 171098 26186 171334
rect 26422 171098 62186 171334
rect 62422 171098 98186 171334
rect 98422 171098 134186 171334
rect 134422 171098 170186 171334
rect 170422 171098 206186 171334
rect 206422 171098 242186 171334
rect 242422 171098 278186 171334
rect 278422 171098 314186 171334
rect 314422 171098 350186 171334
rect 350422 171098 386186 171334
rect 386422 171098 422186 171334
rect 422422 171098 458186 171334
rect 458422 171098 494186 171334
rect 494422 171098 530186 171334
rect 530422 171098 566186 171334
rect 566422 171098 590202 171334
rect 590438 171098 590620 171334
rect -6696 171076 590620 171098
rect -6696 171074 -6096 171076
rect 26004 171074 26604 171076
rect 62004 171074 62604 171076
rect 98004 171074 98604 171076
rect 134004 171074 134604 171076
rect 170004 171074 170604 171076
rect 206004 171074 206604 171076
rect 242004 171074 242604 171076
rect 278004 171074 278604 171076
rect 314004 171074 314604 171076
rect 350004 171074 350604 171076
rect 386004 171074 386604 171076
rect 422004 171074 422604 171076
rect 458004 171074 458604 171076
rect 494004 171074 494604 171076
rect 530004 171074 530604 171076
rect 566004 171074 566604 171076
rect 590020 171074 590620 171076
rect -4816 168076 -4216 168078
rect 22404 168076 23004 168078
rect 58404 168076 59004 168078
rect 94404 168076 95004 168078
rect 130404 168076 131004 168078
rect 166404 168076 167004 168078
rect 202404 168076 203004 168078
rect 238404 168076 239004 168078
rect 274404 168076 275004 168078
rect 310404 168076 311004 168078
rect 346404 168076 347004 168078
rect 382404 168076 383004 168078
rect 418404 168076 419004 168078
rect 454404 168076 455004 168078
rect 490404 168076 491004 168078
rect 526404 168076 527004 168078
rect 562404 168076 563004 168078
rect 588140 168076 588740 168078
rect -4816 168054 588740 168076
rect -4816 167818 -4634 168054
rect -4398 167818 22586 168054
rect 22822 167818 58586 168054
rect 58822 167818 94586 168054
rect 94822 167818 130586 168054
rect 130822 167818 166586 168054
rect 166822 167818 202586 168054
rect 202822 167818 238586 168054
rect 238822 167818 274586 168054
rect 274822 167818 310586 168054
rect 310822 167818 346586 168054
rect 346822 167818 382586 168054
rect 382822 167818 418586 168054
rect 418822 167818 454586 168054
rect 454822 167818 490586 168054
rect 490822 167818 526586 168054
rect 526822 167818 562586 168054
rect 562822 167818 588322 168054
rect 588558 167818 588740 168054
rect -4816 167734 588740 167818
rect -4816 167498 -4634 167734
rect -4398 167498 22586 167734
rect 22822 167498 58586 167734
rect 58822 167498 94586 167734
rect 94822 167498 130586 167734
rect 130822 167498 166586 167734
rect 166822 167498 202586 167734
rect 202822 167498 238586 167734
rect 238822 167498 274586 167734
rect 274822 167498 310586 167734
rect 310822 167498 346586 167734
rect 346822 167498 382586 167734
rect 382822 167498 418586 167734
rect 418822 167498 454586 167734
rect 454822 167498 490586 167734
rect 490822 167498 526586 167734
rect 526822 167498 562586 167734
rect 562822 167498 588322 167734
rect 588558 167498 588740 167734
rect -4816 167476 588740 167498
rect -4816 167474 -4216 167476
rect 22404 167474 23004 167476
rect 58404 167474 59004 167476
rect 94404 167474 95004 167476
rect 130404 167474 131004 167476
rect 166404 167474 167004 167476
rect 202404 167474 203004 167476
rect 238404 167474 239004 167476
rect 274404 167474 275004 167476
rect 310404 167474 311004 167476
rect 346404 167474 347004 167476
rect 382404 167474 383004 167476
rect 418404 167474 419004 167476
rect 454404 167474 455004 167476
rect 490404 167474 491004 167476
rect 526404 167474 527004 167476
rect 562404 167474 563004 167476
rect 588140 167474 588740 167476
rect -2936 164476 -2336 164478
rect 18804 164476 19404 164478
rect 54804 164476 55404 164478
rect 90804 164476 91404 164478
rect 126804 164476 127404 164478
rect 162804 164476 163404 164478
rect 198804 164476 199404 164478
rect 234804 164476 235404 164478
rect 270804 164476 271404 164478
rect 306804 164476 307404 164478
rect 342804 164476 343404 164478
rect 378804 164476 379404 164478
rect 414804 164476 415404 164478
rect 450804 164476 451404 164478
rect 486804 164476 487404 164478
rect 522804 164476 523404 164478
rect 558804 164476 559404 164478
rect 586260 164476 586860 164478
rect -2936 164454 586860 164476
rect -2936 164218 -2754 164454
rect -2518 164218 18986 164454
rect 19222 164218 54986 164454
rect 55222 164218 90986 164454
rect 91222 164218 126986 164454
rect 127222 164218 162986 164454
rect 163222 164218 198986 164454
rect 199222 164218 234986 164454
rect 235222 164218 270986 164454
rect 271222 164218 306986 164454
rect 307222 164218 342986 164454
rect 343222 164218 378986 164454
rect 379222 164218 414986 164454
rect 415222 164218 450986 164454
rect 451222 164218 486986 164454
rect 487222 164218 522986 164454
rect 523222 164218 558986 164454
rect 559222 164218 586442 164454
rect 586678 164218 586860 164454
rect -2936 164134 586860 164218
rect -2936 163898 -2754 164134
rect -2518 163898 18986 164134
rect 19222 163898 54986 164134
rect 55222 163898 90986 164134
rect 91222 163898 126986 164134
rect 127222 163898 162986 164134
rect 163222 163898 198986 164134
rect 199222 163898 234986 164134
rect 235222 163898 270986 164134
rect 271222 163898 306986 164134
rect 307222 163898 342986 164134
rect 343222 163898 378986 164134
rect 379222 163898 414986 164134
rect 415222 163898 450986 164134
rect 451222 163898 486986 164134
rect 487222 163898 522986 164134
rect 523222 163898 558986 164134
rect 559222 163898 586442 164134
rect 586678 163898 586860 164134
rect -2936 163876 586860 163898
rect -2936 163874 -2336 163876
rect 18804 163874 19404 163876
rect 54804 163874 55404 163876
rect 90804 163874 91404 163876
rect 126804 163874 127404 163876
rect 162804 163874 163404 163876
rect 198804 163874 199404 163876
rect 234804 163874 235404 163876
rect 270804 163874 271404 163876
rect 306804 163874 307404 163876
rect 342804 163874 343404 163876
rect 378804 163874 379404 163876
rect 414804 163874 415404 163876
rect 450804 163874 451404 163876
rect 486804 163874 487404 163876
rect 522804 163874 523404 163876
rect 558804 163874 559404 163876
rect 586260 163874 586860 163876
rect -7636 157276 -7036 157278
rect 11604 157276 12204 157278
rect 47604 157276 48204 157278
rect 83604 157276 84204 157278
rect 119604 157276 120204 157278
rect 155604 157276 156204 157278
rect 191604 157276 192204 157278
rect 227604 157276 228204 157278
rect 263604 157276 264204 157278
rect 299604 157276 300204 157278
rect 335604 157276 336204 157278
rect 371604 157276 372204 157278
rect 407604 157276 408204 157278
rect 443604 157276 444204 157278
rect 479604 157276 480204 157278
rect 515604 157276 516204 157278
rect 551604 157276 552204 157278
rect 590960 157276 591560 157278
rect -8576 157254 592500 157276
rect -8576 157018 -7454 157254
rect -7218 157018 11786 157254
rect 12022 157018 47786 157254
rect 48022 157018 83786 157254
rect 84022 157018 119786 157254
rect 120022 157018 155786 157254
rect 156022 157018 191786 157254
rect 192022 157018 227786 157254
rect 228022 157018 263786 157254
rect 264022 157018 299786 157254
rect 300022 157018 335786 157254
rect 336022 157018 371786 157254
rect 372022 157018 407786 157254
rect 408022 157018 443786 157254
rect 444022 157018 479786 157254
rect 480022 157018 515786 157254
rect 516022 157018 551786 157254
rect 552022 157018 591142 157254
rect 591378 157018 592500 157254
rect -8576 156934 592500 157018
rect -8576 156698 -7454 156934
rect -7218 156698 11786 156934
rect 12022 156698 47786 156934
rect 48022 156698 83786 156934
rect 84022 156698 119786 156934
rect 120022 156698 155786 156934
rect 156022 156698 191786 156934
rect 192022 156698 227786 156934
rect 228022 156698 263786 156934
rect 264022 156698 299786 156934
rect 300022 156698 335786 156934
rect 336022 156698 371786 156934
rect 372022 156698 407786 156934
rect 408022 156698 443786 156934
rect 444022 156698 479786 156934
rect 480022 156698 515786 156934
rect 516022 156698 551786 156934
rect 552022 156698 591142 156934
rect 591378 156698 592500 156934
rect -8576 156676 592500 156698
rect -7636 156674 -7036 156676
rect 11604 156674 12204 156676
rect 47604 156674 48204 156676
rect 83604 156674 84204 156676
rect 119604 156674 120204 156676
rect 155604 156674 156204 156676
rect 191604 156674 192204 156676
rect 227604 156674 228204 156676
rect 263604 156674 264204 156676
rect 299604 156674 300204 156676
rect 335604 156674 336204 156676
rect 371604 156674 372204 156676
rect 407604 156674 408204 156676
rect 443604 156674 444204 156676
rect 479604 156674 480204 156676
rect 515604 156674 516204 156676
rect 551604 156674 552204 156676
rect 590960 156674 591560 156676
rect -5756 153676 -5156 153678
rect 8004 153676 8604 153678
rect 44004 153676 44604 153678
rect 80004 153676 80604 153678
rect 116004 153676 116604 153678
rect 152004 153676 152604 153678
rect 188004 153676 188604 153678
rect 224004 153676 224604 153678
rect 260004 153676 260604 153678
rect 296004 153676 296604 153678
rect 332004 153676 332604 153678
rect 368004 153676 368604 153678
rect 404004 153676 404604 153678
rect 440004 153676 440604 153678
rect 476004 153676 476604 153678
rect 512004 153676 512604 153678
rect 548004 153676 548604 153678
rect 589080 153676 589680 153678
rect -6696 153654 590620 153676
rect -6696 153418 -5574 153654
rect -5338 153418 8186 153654
rect 8422 153418 44186 153654
rect 44422 153418 80186 153654
rect 80422 153418 116186 153654
rect 116422 153418 152186 153654
rect 152422 153418 188186 153654
rect 188422 153418 224186 153654
rect 224422 153418 260186 153654
rect 260422 153418 296186 153654
rect 296422 153418 332186 153654
rect 332422 153418 368186 153654
rect 368422 153418 404186 153654
rect 404422 153418 440186 153654
rect 440422 153418 476186 153654
rect 476422 153418 512186 153654
rect 512422 153418 548186 153654
rect 548422 153418 589262 153654
rect 589498 153418 590620 153654
rect -6696 153334 590620 153418
rect -6696 153098 -5574 153334
rect -5338 153098 8186 153334
rect 8422 153098 44186 153334
rect 44422 153098 80186 153334
rect 80422 153098 116186 153334
rect 116422 153098 152186 153334
rect 152422 153098 188186 153334
rect 188422 153098 224186 153334
rect 224422 153098 260186 153334
rect 260422 153098 296186 153334
rect 296422 153098 332186 153334
rect 332422 153098 368186 153334
rect 368422 153098 404186 153334
rect 404422 153098 440186 153334
rect 440422 153098 476186 153334
rect 476422 153098 512186 153334
rect 512422 153098 548186 153334
rect 548422 153098 589262 153334
rect 589498 153098 590620 153334
rect -6696 153076 590620 153098
rect -5756 153074 -5156 153076
rect 8004 153074 8604 153076
rect 44004 153074 44604 153076
rect 80004 153074 80604 153076
rect 116004 153074 116604 153076
rect 152004 153074 152604 153076
rect 188004 153074 188604 153076
rect 224004 153074 224604 153076
rect 260004 153074 260604 153076
rect 296004 153074 296604 153076
rect 332004 153074 332604 153076
rect 368004 153074 368604 153076
rect 404004 153074 404604 153076
rect 440004 153074 440604 153076
rect 476004 153074 476604 153076
rect 512004 153074 512604 153076
rect 548004 153074 548604 153076
rect 589080 153074 589680 153076
rect -3876 150076 -3276 150078
rect 4404 150076 5004 150078
rect 40404 150076 41004 150078
rect 76404 150076 77004 150078
rect 112404 150076 113004 150078
rect 148404 150076 149004 150078
rect 184404 150076 185004 150078
rect 220404 150076 221004 150078
rect 256404 150076 257004 150078
rect 292404 150076 293004 150078
rect 328404 150076 329004 150078
rect 364404 150076 365004 150078
rect 400404 150076 401004 150078
rect 436404 150076 437004 150078
rect 472404 150076 473004 150078
rect 508404 150076 509004 150078
rect 544404 150076 545004 150078
rect 580404 150076 581004 150078
rect 587200 150076 587800 150078
rect -4816 150054 588740 150076
rect -4816 149818 -3694 150054
rect -3458 149818 4586 150054
rect 4822 149818 40586 150054
rect 40822 149818 76586 150054
rect 76822 149818 112586 150054
rect 112822 149818 148586 150054
rect 148822 149818 184586 150054
rect 184822 149818 220586 150054
rect 220822 149818 256586 150054
rect 256822 149818 292586 150054
rect 292822 149818 328586 150054
rect 328822 149818 364586 150054
rect 364822 149818 400586 150054
rect 400822 149818 436586 150054
rect 436822 149818 472586 150054
rect 472822 149818 508586 150054
rect 508822 149818 544586 150054
rect 544822 149818 580586 150054
rect 580822 149818 587382 150054
rect 587618 149818 588740 150054
rect -4816 149734 588740 149818
rect -4816 149498 -3694 149734
rect -3458 149498 4586 149734
rect 4822 149498 40586 149734
rect 40822 149498 76586 149734
rect 76822 149498 112586 149734
rect 112822 149498 148586 149734
rect 148822 149498 184586 149734
rect 184822 149498 220586 149734
rect 220822 149498 256586 149734
rect 256822 149498 292586 149734
rect 292822 149498 328586 149734
rect 328822 149498 364586 149734
rect 364822 149498 400586 149734
rect 400822 149498 436586 149734
rect 436822 149498 472586 149734
rect 472822 149498 508586 149734
rect 508822 149498 544586 149734
rect 544822 149498 580586 149734
rect 580822 149498 587382 149734
rect 587618 149498 588740 149734
rect -4816 149476 588740 149498
rect -3876 149474 -3276 149476
rect 4404 149474 5004 149476
rect 40404 149474 41004 149476
rect 76404 149474 77004 149476
rect 112404 149474 113004 149476
rect 148404 149474 149004 149476
rect 184404 149474 185004 149476
rect 220404 149474 221004 149476
rect 256404 149474 257004 149476
rect 292404 149474 293004 149476
rect 328404 149474 329004 149476
rect 364404 149474 365004 149476
rect 400404 149474 401004 149476
rect 436404 149474 437004 149476
rect 472404 149474 473004 149476
rect 508404 149474 509004 149476
rect 544404 149474 545004 149476
rect 580404 149474 581004 149476
rect 587200 149474 587800 149476
rect -1996 146476 -1396 146478
rect 804 146476 1404 146478
rect 36804 146476 37404 146478
rect 72804 146476 73404 146478
rect 108804 146476 109404 146478
rect 144804 146476 145404 146478
rect 180804 146476 181404 146478
rect 216804 146476 217404 146478
rect 252804 146476 253404 146478
rect 288804 146476 289404 146478
rect 324804 146476 325404 146478
rect 360804 146476 361404 146478
rect 396804 146476 397404 146478
rect 432804 146476 433404 146478
rect 468804 146476 469404 146478
rect 504804 146476 505404 146478
rect 540804 146476 541404 146478
rect 576804 146476 577404 146478
rect 585320 146476 585920 146478
rect -2936 146454 586860 146476
rect -2936 146218 -1814 146454
rect -1578 146218 986 146454
rect 1222 146218 36986 146454
rect 37222 146218 72986 146454
rect 73222 146218 108986 146454
rect 109222 146218 144986 146454
rect 145222 146218 180986 146454
rect 181222 146218 216986 146454
rect 217222 146218 252986 146454
rect 253222 146218 288986 146454
rect 289222 146218 324986 146454
rect 325222 146218 360986 146454
rect 361222 146218 396986 146454
rect 397222 146218 432986 146454
rect 433222 146218 468986 146454
rect 469222 146218 504986 146454
rect 505222 146218 540986 146454
rect 541222 146218 576986 146454
rect 577222 146218 585502 146454
rect 585738 146218 586860 146454
rect -2936 146134 586860 146218
rect -2936 145898 -1814 146134
rect -1578 145898 986 146134
rect 1222 145898 36986 146134
rect 37222 145898 72986 146134
rect 73222 145898 108986 146134
rect 109222 145898 144986 146134
rect 145222 145898 180986 146134
rect 181222 145898 216986 146134
rect 217222 145898 252986 146134
rect 253222 145898 288986 146134
rect 289222 145898 324986 146134
rect 325222 145898 360986 146134
rect 361222 145898 396986 146134
rect 397222 145898 432986 146134
rect 433222 145898 468986 146134
rect 469222 145898 504986 146134
rect 505222 145898 540986 146134
rect 541222 145898 576986 146134
rect 577222 145898 585502 146134
rect 585738 145898 586860 146134
rect -2936 145876 586860 145898
rect -1996 145874 -1396 145876
rect 804 145874 1404 145876
rect 36804 145874 37404 145876
rect 72804 145874 73404 145876
rect 108804 145874 109404 145876
rect 144804 145874 145404 145876
rect 180804 145874 181404 145876
rect 216804 145874 217404 145876
rect 252804 145874 253404 145876
rect 288804 145874 289404 145876
rect 324804 145874 325404 145876
rect 360804 145874 361404 145876
rect 396804 145874 397404 145876
rect 432804 145874 433404 145876
rect 468804 145874 469404 145876
rect 504804 145874 505404 145876
rect 540804 145874 541404 145876
rect 576804 145874 577404 145876
rect 585320 145874 585920 145876
rect -8576 139276 -7976 139278
rect 29604 139276 30204 139278
rect 65604 139276 66204 139278
rect 101604 139276 102204 139278
rect 137604 139276 138204 139278
rect 173604 139276 174204 139278
rect 209604 139276 210204 139278
rect 245604 139276 246204 139278
rect 281604 139276 282204 139278
rect 317604 139276 318204 139278
rect 353604 139276 354204 139278
rect 389604 139276 390204 139278
rect 425604 139276 426204 139278
rect 461604 139276 462204 139278
rect 497604 139276 498204 139278
rect 533604 139276 534204 139278
rect 569604 139276 570204 139278
rect 591900 139276 592500 139278
rect -8576 139254 592500 139276
rect -8576 139018 -8394 139254
rect -8158 139018 29786 139254
rect 30022 139018 65786 139254
rect 66022 139018 101786 139254
rect 102022 139018 137786 139254
rect 138022 139018 173786 139254
rect 174022 139018 209786 139254
rect 210022 139018 245786 139254
rect 246022 139018 281786 139254
rect 282022 139018 317786 139254
rect 318022 139018 353786 139254
rect 354022 139018 389786 139254
rect 390022 139018 425786 139254
rect 426022 139018 461786 139254
rect 462022 139018 497786 139254
rect 498022 139018 533786 139254
rect 534022 139018 569786 139254
rect 570022 139018 592082 139254
rect 592318 139018 592500 139254
rect -8576 138934 592500 139018
rect -8576 138698 -8394 138934
rect -8158 138698 29786 138934
rect 30022 138698 65786 138934
rect 66022 138698 101786 138934
rect 102022 138698 137786 138934
rect 138022 138698 173786 138934
rect 174022 138698 209786 138934
rect 210022 138698 245786 138934
rect 246022 138698 281786 138934
rect 282022 138698 317786 138934
rect 318022 138698 353786 138934
rect 354022 138698 389786 138934
rect 390022 138698 425786 138934
rect 426022 138698 461786 138934
rect 462022 138698 497786 138934
rect 498022 138698 533786 138934
rect 534022 138698 569786 138934
rect 570022 138698 592082 138934
rect 592318 138698 592500 138934
rect -8576 138676 592500 138698
rect -8576 138674 -7976 138676
rect 29604 138674 30204 138676
rect 65604 138674 66204 138676
rect 101604 138674 102204 138676
rect 137604 138674 138204 138676
rect 173604 138674 174204 138676
rect 209604 138674 210204 138676
rect 245604 138674 246204 138676
rect 281604 138674 282204 138676
rect 317604 138674 318204 138676
rect 353604 138674 354204 138676
rect 389604 138674 390204 138676
rect 425604 138674 426204 138676
rect 461604 138674 462204 138676
rect 497604 138674 498204 138676
rect 533604 138674 534204 138676
rect 569604 138674 570204 138676
rect 591900 138674 592500 138676
rect -6696 135676 -6096 135678
rect 26004 135676 26604 135678
rect 62004 135676 62604 135678
rect 98004 135676 98604 135678
rect 134004 135676 134604 135678
rect 170004 135676 170604 135678
rect 206004 135676 206604 135678
rect 242004 135676 242604 135678
rect 278004 135676 278604 135678
rect 314004 135676 314604 135678
rect 350004 135676 350604 135678
rect 386004 135676 386604 135678
rect 422004 135676 422604 135678
rect 458004 135676 458604 135678
rect 494004 135676 494604 135678
rect 530004 135676 530604 135678
rect 566004 135676 566604 135678
rect 590020 135676 590620 135678
rect -6696 135654 590620 135676
rect -6696 135418 -6514 135654
rect -6278 135418 26186 135654
rect 26422 135418 62186 135654
rect 62422 135418 98186 135654
rect 98422 135418 134186 135654
rect 134422 135418 170186 135654
rect 170422 135418 206186 135654
rect 206422 135418 242186 135654
rect 242422 135418 278186 135654
rect 278422 135418 314186 135654
rect 314422 135418 350186 135654
rect 350422 135418 386186 135654
rect 386422 135418 422186 135654
rect 422422 135418 458186 135654
rect 458422 135418 494186 135654
rect 494422 135418 530186 135654
rect 530422 135418 566186 135654
rect 566422 135418 590202 135654
rect 590438 135418 590620 135654
rect -6696 135334 590620 135418
rect -6696 135098 -6514 135334
rect -6278 135098 26186 135334
rect 26422 135098 62186 135334
rect 62422 135098 98186 135334
rect 98422 135098 134186 135334
rect 134422 135098 170186 135334
rect 170422 135098 206186 135334
rect 206422 135098 242186 135334
rect 242422 135098 278186 135334
rect 278422 135098 314186 135334
rect 314422 135098 350186 135334
rect 350422 135098 386186 135334
rect 386422 135098 422186 135334
rect 422422 135098 458186 135334
rect 458422 135098 494186 135334
rect 494422 135098 530186 135334
rect 530422 135098 566186 135334
rect 566422 135098 590202 135334
rect 590438 135098 590620 135334
rect -6696 135076 590620 135098
rect -6696 135074 -6096 135076
rect 26004 135074 26604 135076
rect 62004 135074 62604 135076
rect 98004 135074 98604 135076
rect 134004 135074 134604 135076
rect 170004 135074 170604 135076
rect 206004 135074 206604 135076
rect 242004 135074 242604 135076
rect 278004 135074 278604 135076
rect 314004 135074 314604 135076
rect 350004 135074 350604 135076
rect 386004 135074 386604 135076
rect 422004 135074 422604 135076
rect 458004 135074 458604 135076
rect 494004 135074 494604 135076
rect 530004 135074 530604 135076
rect 566004 135074 566604 135076
rect 590020 135074 590620 135076
rect -4816 132076 -4216 132078
rect 22404 132076 23004 132078
rect 58404 132076 59004 132078
rect 94404 132076 95004 132078
rect 130404 132076 131004 132078
rect 166404 132076 167004 132078
rect 202404 132076 203004 132078
rect 238404 132076 239004 132078
rect 274404 132076 275004 132078
rect 310404 132076 311004 132078
rect 346404 132076 347004 132078
rect 382404 132076 383004 132078
rect 418404 132076 419004 132078
rect 454404 132076 455004 132078
rect 490404 132076 491004 132078
rect 526404 132076 527004 132078
rect 562404 132076 563004 132078
rect 588140 132076 588740 132078
rect -4816 132054 588740 132076
rect -4816 131818 -4634 132054
rect -4398 131818 22586 132054
rect 22822 131818 58586 132054
rect 58822 131818 94586 132054
rect 94822 131818 130586 132054
rect 130822 131818 166586 132054
rect 166822 131818 202586 132054
rect 202822 131818 238586 132054
rect 238822 131818 274586 132054
rect 274822 131818 310586 132054
rect 310822 131818 346586 132054
rect 346822 131818 382586 132054
rect 382822 131818 418586 132054
rect 418822 131818 454586 132054
rect 454822 131818 490586 132054
rect 490822 131818 526586 132054
rect 526822 131818 562586 132054
rect 562822 131818 588322 132054
rect 588558 131818 588740 132054
rect -4816 131734 588740 131818
rect -4816 131498 -4634 131734
rect -4398 131498 22586 131734
rect 22822 131498 58586 131734
rect 58822 131498 94586 131734
rect 94822 131498 130586 131734
rect 130822 131498 166586 131734
rect 166822 131498 202586 131734
rect 202822 131498 238586 131734
rect 238822 131498 274586 131734
rect 274822 131498 310586 131734
rect 310822 131498 346586 131734
rect 346822 131498 382586 131734
rect 382822 131498 418586 131734
rect 418822 131498 454586 131734
rect 454822 131498 490586 131734
rect 490822 131498 526586 131734
rect 526822 131498 562586 131734
rect 562822 131498 588322 131734
rect 588558 131498 588740 131734
rect -4816 131476 588740 131498
rect -4816 131474 -4216 131476
rect 22404 131474 23004 131476
rect 58404 131474 59004 131476
rect 94404 131474 95004 131476
rect 130404 131474 131004 131476
rect 166404 131474 167004 131476
rect 202404 131474 203004 131476
rect 238404 131474 239004 131476
rect 274404 131474 275004 131476
rect 310404 131474 311004 131476
rect 346404 131474 347004 131476
rect 382404 131474 383004 131476
rect 418404 131474 419004 131476
rect 454404 131474 455004 131476
rect 490404 131474 491004 131476
rect 526404 131474 527004 131476
rect 562404 131474 563004 131476
rect 588140 131474 588740 131476
rect -2936 128476 -2336 128478
rect 18804 128476 19404 128478
rect 54804 128476 55404 128478
rect 90804 128476 91404 128478
rect 126804 128476 127404 128478
rect 162804 128476 163404 128478
rect 198804 128476 199404 128478
rect 234804 128476 235404 128478
rect 270804 128476 271404 128478
rect 306804 128476 307404 128478
rect 342804 128476 343404 128478
rect 378804 128476 379404 128478
rect 414804 128476 415404 128478
rect 450804 128476 451404 128478
rect 486804 128476 487404 128478
rect 522804 128476 523404 128478
rect 558804 128476 559404 128478
rect 586260 128476 586860 128478
rect -2936 128454 586860 128476
rect -2936 128218 -2754 128454
rect -2518 128218 18986 128454
rect 19222 128218 54986 128454
rect 55222 128218 90986 128454
rect 91222 128218 126986 128454
rect 127222 128218 162986 128454
rect 163222 128218 198986 128454
rect 199222 128218 234986 128454
rect 235222 128218 270986 128454
rect 271222 128218 306986 128454
rect 307222 128218 342986 128454
rect 343222 128218 378986 128454
rect 379222 128218 414986 128454
rect 415222 128218 450986 128454
rect 451222 128218 486986 128454
rect 487222 128218 522986 128454
rect 523222 128218 558986 128454
rect 559222 128218 586442 128454
rect 586678 128218 586860 128454
rect -2936 128134 586860 128218
rect -2936 127898 -2754 128134
rect -2518 127898 18986 128134
rect 19222 127898 54986 128134
rect 55222 127898 90986 128134
rect 91222 127898 126986 128134
rect 127222 127898 162986 128134
rect 163222 127898 198986 128134
rect 199222 127898 234986 128134
rect 235222 127898 270986 128134
rect 271222 127898 306986 128134
rect 307222 127898 342986 128134
rect 343222 127898 378986 128134
rect 379222 127898 414986 128134
rect 415222 127898 450986 128134
rect 451222 127898 486986 128134
rect 487222 127898 522986 128134
rect 523222 127898 558986 128134
rect 559222 127898 586442 128134
rect 586678 127898 586860 128134
rect -2936 127876 586860 127898
rect -2936 127874 -2336 127876
rect 18804 127874 19404 127876
rect 54804 127874 55404 127876
rect 90804 127874 91404 127876
rect 126804 127874 127404 127876
rect 162804 127874 163404 127876
rect 198804 127874 199404 127876
rect 234804 127874 235404 127876
rect 270804 127874 271404 127876
rect 306804 127874 307404 127876
rect 342804 127874 343404 127876
rect 378804 127874 379404 127876
rect 414804 127874 415404 127876
rect 450804 127874 451404 127876
rect 486804 127874 487404 127876
rect 522804 127874 523404 127876
rect 558804 127874 559404 127876
rect 586260 127874 586860 127876
rect -7636 121276 -7036 121278
rect 11604 121276 12204 121278
rect 47604 121276 48204 121278
rect 83604 121276 84204 121278
rect 119604 121276 120204 121278
rect 155604 121276 156204 121278
rect 191604 121276 192204 121278
rect 227604 121276 228204 121278
rect 263604 121276 264204 121278
rect 299604 121276 300204 121278
rect 335604 121276 336204 121278
rect 371604 121276 372204 121278
rect 407604 121276 408204 121278
rect 443604 121276 444204 121278
rect 479604 121276 480204 121278
rect 515604 121276 516204 121278
rect 551604 121276 552204 121278
rect 590960 121276 591560 121278
rect -8576 121254 592500 121276
rect -8576 121018 -7454 121254
rect -7218 121018 11786 121254
rect 12022 121018 47786 121254
rect 48022 121018 83786 121254
rect 84022 121018 119786 121254
rect 120022 121018 155786 121254
rect 156022 121018 191786 121254
rect 192022 121018 227786 121254
rect 228022 121018 263786 121254
rect 264022 121018 299786 121254
rect 300022 121018 335786 121254
rect 336022 121018 371786 121254
rect 372022 121018 407786 121254
rect 408022 121018 443786 121254
rect 444022 121018 479786 121254
rect 480022 121018 515786 121254
rect 516022 121018 551786 121254
rect 552022 121018 591142 121254
rect 591378 121018 592500 121254
rect -8576 120934 592500 121018
rect -8576 120698 -7454 120934
rect -7218 120698 11786 120934
rect 12022 120698 47786 120934
rect 48022 120698 83786 120934
rect 84022 120698 119786 120934
rect 120022 120698 155786 120934
rect 156022 120698 191786 120934
rect 192022 120698 227786 120934
rect 228022 120698 263786 120934
rect 264022 120698 299786 120934
rect 300022 120698 335786 120934
rect 336022 120698 371786 120934
rect 372022 120698 407786 120934
rect 408022 120698 443786 120934
rect 444022 120698 479786 120934
rect 480022 120698 515786 120934
rect 516022 120698 551786 120934
rect 552022 120698 591142 120934
rect 591378 120698 592500 120934
rect -8576 120676 592500 120698
rect -7636 120674 -7036 120676
rect 11604 120674 12204 120676
rect 47604 120674 48204 120676
rect 83604 120674 84204 120676
rect 119604 120674 120204 120676
rect 155604 120674 156204 120676
rect 191604 120674 192204 120676
rect 227604 120674 228204 120676
rect 263604 120674 264204 120676
rect 299604 120674 300204 120676
rect 335604 120674 336204 120676
rect 371604 120674 372204 120676
rect 407604 120674 408204 120676
rect 443604 120674 444204 120676
rect 479604 120674 480204 120676
rect 515604 120674 516204 120676
rect 551604 120674 552204 120676
rect 590960 120674 591560 120676
rect -5756 117676 -5156 117678
rect 8004 117676 8604 117678
rect 44004 117676 44604 117678
rect 80004 117676 80604 117678
rect 116004 117676 116604 117678
rect 152004 117676 152604 117678
rect 188004 117676 188604 117678
rect 224004 117676 224604 117678
rect 260004 117676 260604 117678
rect 296004 117676 296604 117678
rect 332004 117676 332604 117678
rect 368004 117676 368604 117678
rect 404004 117676 404604 117678
rect 440004 117676 440604 117678
rect 476004 117676 476604 117678
rect 512004 117676 512604 117678
rect 548004 117676 548604 117678
rect 589080 117676 589680 117678
rect -6696 117654 590620 117676
rect -6696 117418 -5574 117654
rect -5338 117418 8186 117654
rect 8422 117418 44186 117654
rect 44422 117418 80186 117654
rect 80422 117418 116186 117654
rect 116422 117418 152186 117654
rect 152422 117418 188186 117654
rect 188422 117418 224186 117654
rect 224422 117418 260186 117654
rect 260422 117418 296186 117654
rect 296422 117418 332186 117654
rect 332422 117418 368186 117654
rect 368422 117418 404186 117654
rect 404422 117418 440186 117654
rect 440422 117418 476186 117654
rect 476422 117418 512186 117654
rect 512422 117418 548186 117654
rect 548422 117418 589262 117654
rect 589498 117418 590620 117654
rect -6696 117334 590620 117418
rect -6696 117098 -5574 117334
rect -5338 117098 8186 117334
rect 8422 117098 44186 117334
rect 44422 117098 80186 117334
rect 80422 117098 116186 117334
rect 116422 117098 152186 117334
rect 152422 117098 188186 117334
rect 188422 117098 224186 117334
rect 224422 117098 260186 117334
rect 260422 117098 296186 117334
rect 296422 117098 332186 117334
rect 332422 117098 368186 117334
rect 368422 117098 404186 117334
rect 404422 117098 440186 117334
rect 440422 117098 476186 117334
rect 476422 117098 512186 117334
rect 512422 117098 548186 117334
rect 548422 117098 589262 117334
rect 589498 117098 590620 117334
rect -6696 117076 590620 117098
rect -5756 117074 -5156 117076
rect 8004 117074 8604 117076
rect 44004 117074 44604 117076
rect 80004 117074 80604 117076
rect 116004 117074 116604 117076
rect 152004 117074 152604 117076
rect 188004 117074 188604 117076
rect 224004 117074 224604 117076
rect 260004 117074 260604 117076
rect 296004 117074 296604 117076
rect 332004 117074 332604 117076
rect 368004 117074 368604 117076
rect 404004 117074 404604 117076
rect 440004 117074 440604 117076
rect 476004 117074 476604 117076
rect 512004 117074 512604 117076
rect 548004 117074 548604 117076
rect 589080 117074 589680 117076
rect -3876 114076 -3276 114078
rect 4404 114076 5004 114078
rect 40404 114076 41004 114078
rect 76404 114076 77004 114078
rect 112404 114076 113004 114078
rect 148404 114076 149004 114078
rect 184404 114076 185004 114078
rect 220404 114076 221004 114078
rect 256404 114076 257004 114078
rect 292404 114076 293004 114078
rect 328404 114076 329004 114078
rect 364404 114076 365004 114078
rect 400404 114076 401004 114078
rect 436404 114076 437004 114078
rect 472404 114076 473004 114078
rect 508404 114076 509004 114078
rect 544404 114076 545004 114078
rect 580404 114076 581004 114078
rect 587200 114076 587800 114078
rect -4816 114054 588740 114076
rect -4816 113818 -3694 114054
rect -3458 113818 4586 114054
rect 4822 113818 40586 114054
rect 40822 113818 76586 114054
rect 76822 113818 112586 114054
rect 112822 113818 148586 114054
rect 148822 113818 184586 114054
rect 184822 113818 220586 114054
rect 220822 113818 256586 114054
rect 256822 113818 292586 114054
rect 292822 113818 328586 114054
rect 328822 113818 364586 114054
rect 364822 113818 400586 114054
rect 400822 113818 436586 114054
rect 436822 113818 472586 114054
rect 472822 113818 508586 114054
rect 508822 113818 544586 114054
rect 544822 113818 580586 114054
rect 580822 113818 587382 114054
rect 587618 113818 588740 114054
rect -4816 113734 588740 113818
rect -4816 113498 -3694 113734
rect -3458 113498 4586 113734
rect 4822 113498 40586 113734
rect 40822 113498 76586 113734
rect 76822 113498 112586 113734
rect 112822 113498 148586 113734
rect 148822 113498 184586 113734
rect 184822 113498 220586 113734
rect 220822 113498 256586 113734
rect 256822 113498 292586 113734
rect 292822 113498 328586 113734
rect 328822 113498 364586 113734
rect 364822 113498 400586 113734
rect 400822 113498 436586 113734
rect 436822 113498 472586 113734
rect 472822 113498 508586 113734
rect 508822 113498 544586 113734
rect 544822 113498 580586 113734
rect 580822 113498 587382 113734
rect 587618 113498 588740 113734
rect -4816 113476 588740 113498
rect -3876 113474 -3276 113476
rect 4404 113474 5004 113476
rect 40404 113474 41004 113476
rect 76404 113474 77004 113476
rect 112404 113474 113004 113476
rect 148404 113474 149004 113476
rect 184404 113474 185004 113476
rect 220404 113474 221004 113476
rect 256404 113474 257004 113476
rect 292404 113474 293004 113476
rect 328404 113474 329004 113476
rect 364404 113474 365004 113476
rect 400404 113474 401004 113476
rect 436404 113474 437004 113476
rect 472404 113474 473004 113476
rect 508404 113474 509004 113476
rect 544404 113474 545004 113476
rect 580404 113474 581004 113476
rect 587200 113474 587800 113476
rect -1996 110476 -1396 110478
rect 804 110476 1404 110478
rect 36804 110476 37404 110478
rect 72804 110476 73404 110478
rect 108804 110476 109404 110478
rect 144804 110476 145404 110478
rect 180804 110476 181404 110478
rect 216804 110476 217404 110478
rect 252804 110476 253404 110478
rect 288804 110476 289404 110478
rect 324804 110476 325404 110478
rect 360804 110476 361404 110478
rect 396804 110476 397404 110478
rect 432804 110476 433404 110478
rect 468804 110476 469404 110478
rect 504804 110476 505404 110478
rect 540804 110476 541404 110478
rect 576804 110476 577404 110478
rect 585320 110476 585920 110478
rect -2936 110454 586860 110476
rect -2936 110218 -1814 110454
rect -1578 110218 986 110454
rect 1222 110218 36986 110454
rect 37222 110218 72986 110454
rect 73222 110218 108986 110454
rect 109222 110218 144986 110454
rect 145222 110218 180986 110454
rect 181222 110218 216986 110454
rect 217222 110218 252986 110454
rect 253222 110218 288986 110454
rect 289222 110218 324986 110454
rect 325222 110218 360986 110454
rect 361222 110218 396986 110454
rect 397222 110218 432986 110454
rect 433222 110218 468986 110454
rect 469222 110218 504986 110454
rect 505222 110218 540986 110454
rect 541222 110218 576986 110454
rect 577222 110218 585502 110454
rect 585738 110218 586860 110454
rect -2936 110134 586860 110218
rect -2936 109898 -1814 110134
rect -1578 109898 986 110134
rect 1222 109898 36986 110134
rect 37222 109898 72986 110134
rect 73222 109898 108986 110134
rect 109222 109898 144986 110134
rect 145222 109898 180986 110134
rect 181222 109898 216986 110134
rect 217222 109898 252986 110134
rect 253222 109898 288986 110134
rect 289222 109898 324986 110134
rect 325222 109898 360986 110134
rect 361222 109898 396986 110134
rect 397222 109898 432986 110134
rect 433222 109898 468986 110134
rect 469222 109898 504986 110134
rect 505222 109898 540986 110134
rect 541222 109898 576986 110134
rect 577222 109898 585502 110134
rect 585738 109898 586860 110134
rect -2936 109876 586860 109898
rect -1996 109874 -1396 109876
rect 804 109874 1404 109876
rect 36804 109874 37404 109876
rect 72804 109874 73404 109876
rect 108804 109874 109404 109876
rect 144804 109874 145404 109876
rect 180804 109874 181404 109876
rect 216804 109874 217404 109876
rect 252804 109874 253404 109876
rect 288804 109874 289404 109876
rect 324804 109874 325404 109876
rect 360804 109874 361404 109876
rect 396804 109874 397404 109876
rect 432804 109874 433404 109876
rect 468804 109874 469404 109876
rect 504804 109874 505404 109876
rect 540804 109874 541404 109876
rect 576804 109874 577404 109876
rect 585320 109874 585920 109876
rect -8576 103276 -7976 103278
rect 29604 103276 30204 103278
rect 65604 103276 66204 103278
rect 101604 103276 102204 103278
rect 137604 103276 138204 103278
rect 173604 103276 174204 103278
rect 209604 103276 210204 103278
rect 245604 103276 246204 103278
rect 281604 103276 282204 103278
rect 317604 103276 318204 103278
rect 353604 103276 354204 103278
rect 389604 103276 390204 103278
rect 425604 103276 426204 103278
rect 461604 103276 462204 103278
rect 497604 103276 498204 103278
rect 533604 103276 534204 103278
rect 569604 103276 570204 103278
rect 591900 103276 592500 103278
rect -8576 103254 592500 103276
rect -8576 103018 -8394 103254
rect -8158 103018 29786 103254
rect 30022 103018 65786 103254
rect 66022 103018 101786 103254
rect 102022 103018 137786 103254
rect 138022 103018 173786 103254
rect 174022 103018 209786 103254
rect 210022 103018 245786 103254
rect 246022 103018 281786 103254
rect 282022 103018 317786 103254
rect 318022 103018 353786 103254
rect 354022 103018 389786 103254
rect 390022 103018 425786 103254
rect 426022 103018 461786 103254
rect 462022 103018 497786 103254
rect 498022 103018 533786 103254
rect 534022 103018 569786 103254
rect 570022 103018 592082 103254
rect 592318 103018 592500 103254
rect -8576 102934 592500 103018
rect -8576 102698 -8394 102934
rect -8158 102698 29786 102934
rect 30022 102698 65786 102934
rect 66022 102698 101786 102934
rect 102022 102698 137786 102934
rect 138022 102698 173786 102934
rect 174022 102698 209786 102934
rect 210022 102698 245786 102934
rect 246022 102698 281786 102934
rect 282022 102698 317786 102934
rect 318022 102698 353786 102934
rect 354022 102698 389786 102934
rect 390022 102698 425786 102934
rect 426022 102698 461786 102934
rect 462022 102698 497786 102934
rect 498022 102698 533786 102934
rect 534022 102698 569786 102934
rect 570022 102698 592082 102934
rect 592318 102698 592500 102934
rect -8576 102676 592500 102698
rect -8576 102674 -7976 102676
rect 29604 102674 30204 102676
rect 65604 102674 66204 102676
rect 101604 102674 102204 102676
rect 137604 102674 138204 102676
rect 173604 102674 174204 102676
rect 209604 102674 210204 102676
rect 245604 102674 246204 102676
rect 281604 102674 282204 102676
rect 317604 102674 318204 102676
rect 353604 102674 354204 102676
rect 389604 102674 390204 102676
rect 425604 102674 426204 102676
rect 461604 102674 462204 102676
rect 497604 102674 498204 102676
rect 533604 102674 534204 102676
rect 569604 102674 570204 102676
rect 591900 102674 592500 102676
rect -6696 99676 -6096 99678
rect 26004 99676 26604 99678
rect 62004 99676 62604 99678
rect 98004 99676 98604 99678
rect 134004 99676 134604 99678
rect 170004 99676 170604 99678
rect 206004 99676 206604 99678
rect 242004 99676 242604 99678
rect 278004 99676 278604 99678
rect 314004 99676 314604 99678
rect 350004 99676 350604 99678
rect 386004 99676 386604 99678
rect 422004 99676 422604 99678
rect 458004 99676 458604 99678
rect 494004 99676 494604 99678
rect 530004 99676 530604 99678
rect 566004 99676 566604 99678
rect 590020 99676 590620 99678
rect -6696 99654 590620 99676
rect -6696 99418 -6514 99654
rect -6278 99418 26186 99654
rect 26422 99418 62186 99654
rect 62422 99418 98186 99654
rect 98422 99418 134186 99654
rect 134422 99418 170186 99654
rect 170422 99418 206186 99654
rect 206422 99418 242186 99654
rect 242422 99418 278186 99654
rect 278422 99418 314186 99654
rect 314422 99418 350186 99654
rect 350422 99418 386186 99654
rect 386422 99418 422186 99654
rect 422422 99418 458186 99654
rect 458422 99418 494186 99654
rect 494422 99418 530186 99654
rect 530422 99418 566186 99654
rect 566422 99418 590202 99654
rect 590438 99418 590620 99654
rect -6696 99334 590620 99418
rect -6696 99098 -6514 99334
rect -6278 99098 26186 99334
rect 26422 99098 62186 99334
rect 62422 99098 98186 99334
rect 98422 99098 134186 99334
rect 134422 99098 170186 99334
rect 170422 99098 206186 99334
rect 206422 99098 242186 99334
rect 242422 99098 278186 99334
rect 278422 99098 314186 99334
rect 314422 99098 350186 99334
rect 350422 99098 386186 99334
rect 386422 99098 422186 99334
rect 422422 99098 458186 99334
rect 458422 99098 494186 99334
rect 494422 99098 530186 99334
rect 530422 99098 566186 99334
rect 566422 99098 590202 99334
rect 590438 99098 590620 99334
rect -6696 99076 590620 99098
rect -6696 99074 -6096 99076
rect 26004 99074 26604 99076
rect 62004 99074 62604 99076
rect 98004 99074 98604 99076
rect 134004 99074 134604 99076
rect 170004 99074 170604 99076
rect 206004 99074 206604 99076
rect 242004 99074 242604 99076
rect 278004 99074 278604 99076
rect 314004 99074 314604 99076
rect 350004 99074 350604 99076
rect 386004 99074 386604 99076
rect 422004 99074 422604 99076
rect 458004 99074 458604 99076
rect 494004 99074 494604 99076
rect 530004 99074 530604 99076
rect 566004 99074 566604 99076
rect 590020 99074 590620 99076
rect -4816 96076 -4216 96078
rect 22404 96076 23004 96078
rect 58404 96076 59004 96078
rect 94404 96076 95004 96078
rect 130404 96076 131004 96078
rect 166404 96076 167004 96078
rect 202404 96076 203004 96078
rect 238404 96076 239004 96078
rect 274404 96076 275004 96078
rect 310404 96076 311004 96078
rect 346404 96076 347004 96078
rect 382404 96076 383004 96078
rect 418404 96076 419004 96078
rect 454404 96076 455004 96078
rect 490404 96076 491004 96078
rect 526404 96076 527004 96078
rect 562404 96076 563004 96078
rect 588140 96076 588740 96078
rect -4816 96054 588740 96076
rect -4816 95818 -4634 96054
rect -4398 95818 22586 96054
rect 22822 95818 58586 96054
rect 58822 95818 94586 96054
rect 94822 95818 130586 96054
rect 130822 95818 166586 96054
rect 166822 95818 202586 96054
rect 202822 95818 238586 96054
rect 238822 95818 274586 96054
rect 274822 95818 310586 96054
rect 310822 95818 346586 96054
rect 346822 95818 382586 96054
rect 382822 95818 418586 96054
rect 418822 95818 454586 96054
rect 454822 95818 490586 96054
rect 490822 95818 526586 96054
rect 526822 95818 562586 96054
rect 562822 95818 588322 96054
rect 588558 95818 588740 96054
rect -4816 95734 588740 95818
rect -4816 95498 -4634 95734
rect -4398 95498 22586 95734
rect 22822 95498 58586 95734
rect 58822 95498 94586 95734
rect 94822 95498 130586 95734
rect 130822 95498 166586 95734
rect 166822 95498 202586 95734
rect 202822 95498 238586 95734
rect 238822 95498 274586 95734
rect 274822 95498 310586 95734
rect 310822 95498 346586 95734
rect 346822 95498 382586 95734
rect 382822 95498 418586 95734
rect 418822 95498 454586 95734
rect 454822 95498 490586 95734
rect 490822 95498 526586 95734
rect 526822 95498 562586 95734
rect 562822 95498 588322 95734
rect 588558 95498 588740 95734
rect -4816 95476 588740 95498
rect -4816 95474 -4216 95476
rect 22404 95474 23004 95476
rect 58404 95474 59004 95476
rect 94404 95474 95004 95476
rect 130404 95474 131004 95476
rect 166404 95474 167004 95476
rect 202404 95474 203004 95476
rect 238404 95474 239004 95476
rect 274404 95474 275004 95476
rect 310404 95474 311004 95476
rect 346404 95474 347004 95476
rect 382404 95474 383004 95476
rect 418404 95474 419004 95476
rect 454404 95474 455004 95476
rect 490404 95474 491004 95476
rect 526404 95474 527004 95476
rect 562404 95474 563004 95476
rect 588140 95474 588740 95476
rect -2936 92476 -2336 92478
rect 18804 92476 19404 92478
rect 54804 92476 55404 92478
rect 90804 92476 91404 92478
rect 126804 92476 127404 92478
rect 162804 92476 163404 92478
rect 198804 92476 199404 92478
rect 234804 92476 235404 92478
rect 270804 92476 271404 92478
rect 306804 92476 307404 92478
rect 342804 92476 343404 92478
rect 378804 92476 379404 92478
rect 414804 92476 415404 92478
rect 450804 92476 451404 92478
rect 486804 92476 487404 92478
rect 522804 92476 523404 92478
rect 558804 92476 559404 92478
rect 586260 92476 586860 92478
rect -2936 92454 586860 92476
rect -2936 92218 -2754 92454
rect -2518 92218 18986 92454
rect 19222 92218 54986 92454
rect 55222 92218 90986 92454
rect 91222 92218 126986 92454
rect 127222 92218 162986 92454
rect 163222 92218 198986 92454
rect 199222 92218 234986 92454
rect 235222 92218 270986 92454
rect 271222 92218 306986 92454
rect 307222 92218 342986 92454
rect 343222 92218 378986 92454
rect 379222 92218 414986 92454
rect 415222 92218 450986 92454
rect 451222 92218 486986 92454
rect 487222 92218 522986 92454
rect 523222 92218 558986 92454
rect 559222 92218 586442 92454
rect 586678 92218 586860 92454
rect -2936 92134 586860 92218
rect -2936 91898 -2754 92134
rect -2518 91898 18986 92134
rect 19222 91898 54986 92134
rect 55222 91898 90986 92134
rect 91222 91898 126986 92134
rect 127222 91898 162986 92134
rect 163222 91898 198986 92134
rect 199222 91898 234986 92134
rect 235222 91898 270986 92134
rect 271222 91898 306986 92134
rect 307222 91898 342986 92134
rect 343222 91898 378986 92134
rect 379222 91898 414986 92134
rect 415222 91898 450986 92134
rect 451222 91898 486986 92134
rect 487222 91898 522986 92134
rect 523222 91898 558986 92134
rect 559222 91898 586442 92134
rect 586678 91898 586860 92134
rect -2936 91876 586860 91898
rect -2936 91874 -2336 91876
rect 18804 91874 19404 91876
rect 54804 91874 55404 91876
rect 90804 91874 91404 91876
rect 126804 91874 127404 91876
rect 162804 91874 163404 91876
rect 198804 91874 199404 91876
rect 234804 91874 235404 91876
rect 270804 91874 271404 91876
rect 306804 91874 307404 91876
rect 342804 91874 343404 91876
rect 378804 91874 379404 91876
rect 414804 91874 415404 91876
rect 450804 91874 451404 91876
rect 486804 91874 487404 91876
rect 522804 91874 523404 91876
rect 558804 91874 559404 91876
rect 586260 91874 586860 91876
rect -7636 85276 -7036 85278
rect 11604 85276 12204 85278
rect 47604 85276 48204 85278
rect 83604 85276 84204 85278
rect 119604 85276 120204 85278
rect 155604 85276 156204 85278
rect 191604 85276 192204 85278
rect 227604 85276 228204 85278
rect 263604 85276 264204 85278
rect 299604 85276 300204 85278
rect 335604 85276 336204 85278
rect 371604 85276 372204 85278
rect 407604 85276 408204 85278
rect 443604 85276 444204 85278
rect 479604 85276 480204 85278
rect 515604 85276 516204 85278
rect 551604 85276 552204 85278
rect 590960 85276 591560 85278
rect -8576 85254 592500 85276
rect -8576 85018 -7454 85254
rect -7218 85018 11786 85254
rect 12022 85018 47786 85254
rect 48022 85018 83786 85254
rect 84022 85018 119786 85254
rect 120022 85018 155786 85254
rect 156022 85018 191786 85254
rect 192022 85018 227786 85254
rect 228022 85018 263786 85254
rect 264022 85018 299786 85254
rect 300022 85018 335786 85254
rect 336022 85018 371786 85254
rect 372022 85018 407786 85254
rect 408022 85018 443786 85254
rect 444022 85018 479786 85254
rect 480022 85018 515786 85254
rect 516022 85018 551786 85254
rect 552022 85018 591142 85254
rect 591378 85018 592500 85254
rect -8576 84934 592500 85018
rect -8576 84698 -7454 84934
rect -7218 84698 11786 84934
rect 12022 84698 47786 84934
rect 48022 84698 83786 84934
rect 84022 84698 119786 84934
rect 120022 84698 155786 84934
rect 156022 84698 191786 84934
rect 192022 84698 227786 84934
rect 228022 84698 263786 84934
rect 264022 84698 299786 84934
rect 300022 84698 335786 84934
rect 336022 84698 371786 84934
rect 372022 84698 407786 84934
rect 408022 84698 443786 84934
rect 444022 84698 479786 84934
rect 480022 84698 515786 84934
rect 516022 84698 551786 84934
rect 552022 84698 591142 84934
rect 591378 84698 592500 84934
rect -8576 84676 592500 84698
rect -7636 84674 -7036 84676
rect 11604 84674 12204 84676
rect 47604 84674 48204 84676
rect 83604 84674 84204 84676
rect 119604 84674 120204 84676
rect 155604 84674 156204 84676
rect 191604 84674 192204 84676
rect 227604 84674 228204 84676
rect 263604 84674 264204 84676
rect 299604 84674 300204 84676
rect 335604 84674 336204 84676
rect 371604 84674 372204 84676
rect 407604 84674 408204 84676
rect 443604 84674 444204 84676
rect 479604 84674 480204 84676
rect 515604 84674 516204 84676
rect 551604 84674 552204 84676
rect 590960 84674 591560 84676
rect -5756 81676 -5156 81678
rect 8004 81676 8604 81678
rect 44004 81676 44604 81678
rect 80004 81676 80604 81678
rect 116004 81676 116604 81678
rect 152004 81676 152604 81678
rect 188004 81676 188604 81678
rect 224004 81676 224604 81678
rect 260004 81676 260604 81678
rect 296004 81676 296604 81678
rect 332004 81676 332604 81678
rect 368004 81676 368604 81678
rect 404004 81676 404604 81678
rect 440004 81676 440604 81678
rect 476004 81676 476604 81678
rect 512004 81676 512604 81678
rect 548004 81676 548604 81678
rect 589080 81676 589680 81678
rect -6696 81654 590620 81676
rect -6696 81418 -5574 81654
rect -5338 81418 8186 81654
rect 8422 81418 44186 81654
rect 44422 81418 80186 81654
rect 80422 81418 116186 81654
rect 116422 81418 152186 81654
rect 152422 81418 188186 81654
rect 188422 81418 224186 81654
rect 224422 81418 260186 81654
rect 260422 81418 296186 81654
rect 296422 81418 332186 81654
rect 332422 81418 368186 81654
rect 368422 81418 404186 81654
rect 404422 81418 440186 81654
rect 440422 81418 476186 81654
rect 476422 81418 512186 81654
rect 512422 81418 548186 81654
rect 548422 81418 589262 81654
rect 589498 81418 590620 81654
rect -6696 81334 590620 81418
rect -6696 81098 -5574 81334
rect -5338 81098 8186 81334
rect 8422 81098 44186 81334
rect 44422 81098 80186 81334
rect 80422 81098 116186 81334
rect 116422 81098 152186 81334
rect 152422 81098 188186 81334
rect 188422 81098 224186 81334
rect 224422 81098 260186 81334
rect 260422 81098 296186 81334
rect 296422 81098 332186 81334
rect 332422 81098 368186 81334
rect 368422 81098 404186 81334
rect 404422 81098 440186 81334
rect 440422 81098 476186 81334
rect 476422 81098 512186 81334
rect 512422 81098 548186 81334
rect 548422 81098 589262 81334
rect 589498 81098 590620 81334
rect -6696 81076 590620 81098
rect -5756 81074 -5156 81076
rect 8004 81074 8604 81076
rect 44004 81074 44604 81076
rect 80004 81074 80604 81076
rect 116004 81074 116604 81076
rect 152004 81074 152604 81076
rect 188004 81074 188604 81076
rect 224004 81074 224604 81076
rect 260004 81074 260604 81076
rect 296004 81074 296604 81076
rect 332004 81074 332604 81076
rect 368004 81074 368604 81076
rect 404004 81074 404604 81076
rect 440004 81074 440604 81076
rect 476004 81074 476604 81076
rect 512004 81074 512604 81076
rect 548004 81074 548604 81076
rect 589080 81074 589680 81076
rect -3876 78076 -3276 78078
rect 4404 78076 5004 78078
rect 40404 78076 41004 78078
rect 76404 78076 77004 78078
rect 112404 78076 113004 78078
rect 148404 78076 149004 78078
rect 184404 78076 185004 78078
rect 220404 78076 221004 78078
rect 256404 78076 257004 78078
rect 292404 78076 293004 78078
rect 328404 78076 329004 78078
rect 364404 78076 365004 78078
rect 400404 78076 401004 78078
rect 436404 78076 437004 78078
rect 472404 78076 473004 78078
rect 508404 78076 509004 78078
rect 544404 78076 545004 78078
rect 580404 78076 581004 78078
rect 587200 78076 587800 78078
rect -4816 78054 588740 78076
rect -4816 77818 -3694 78054
rect -3458 77818 4586 78054
rect 4822 77818 40586 78054
rect 40822 77818 76586 78054
rect 76822 77818 112586 78054
rect 112822 77818 148586 78054
rect 148822 77818 184586 78054
rect 184822 77818 220586 78054
rect 220822 77818 256586 78054
rect 256822 77818 292586 78054
rect 292822 77818 328586 78054
rect 328822 77818 364586 78054
rect 364822 77818 400586 78054
rect 400822 77818 436586 78054
rect 436822 77818 472586 78054
rect 472822 77818 508586 78054
rect 508822 77818 544586 78054
rect 544822 77818 580586 78054
rect 580822 77818 587382 78054
rect 587618 77818 588740 78054
rect -4816 77734 588740 77818
rect -4816 77498 -3694 77734
rect -3458 77498 4586 77734
rect 4822 77498 40586 77734
rect 40822 77498 76586 77734
rect 76822 77498 112586 77734
rect 112822 77498 148586 77734
rect 148822 77498 184586 77734
rect 184822 77498 220586 77734
rect 220822 77498 256586 77734
rect 256822 77498 292586 77734
rect 292822 77498 328586 77734
rect 328822 77498 364586 77734
rect 364822 77498 400586 77734
rect 400822 77498 436586 77734
rect 436822 77498 472586 77734
rect 472822 77498 508586 77734
rect 508822 77498 544586 77734
rect 544822 77498 580586 77734
rect 580822 77498 587382 77734
rect 587618 77498 588740 77734
rect -4816 77476 588740 77498
rect -3876 77474 -3276 77476
rect 4404 77474 5004 77476
rect 40404 77474 41004 77476
rect 76404 77474 77004 77476
rect 112404 77474 113004 77476
rect 148404 77474 149004 77476
rect 184404 77474 185004 77476
rect 220404 77474 221004 77476
rect 256404 77474 257004 77476
rect 292404 77474 293004 77476
rect 328404 77474 329004 77476
rect 364404 77474 365004 77476
rect 400404 77474 401004 77476
rect 436404 77474 437004 77476
rect 472404 77474 473004 77476
rect 508404 77474 509004 77476
rect 544404 77474 545004 77476
rect 580404 77474 581004 77476
rect 587200 77474 587800 77476
rect -1996 74476 -1396 74478
rect 804 74476 1404 74478
rect 36804 74476 37404 74478
rect 72804 74476 73404 74478
rect 108804 74476 109404 74478
rect 144804 74476 145404 74478
rect 180804 74476 181404 74478
rect 216804 74476 217404 74478
rect 252804 74476 253404 74478
rect 288804 74476 289404 74478
rect 324804 74476 325404 74478
rect 360804 74476 361404 74478
rect 396804 74476 397404 74478
rect 432804 74476 433404 74478
rect 468804 74476 469404 74478
rect 504804 74476 505404 74478
rect 540804 74476 541404 74478
rect 576804 74476 577404 74478
rect 585320 74476 585920 74478
rect -2936 74454 586860 74476
rect -2936 74218 -1814 74454
rect -1578 74218 986 74454
rect 1222 74218 36986 74454
rect 37222 74218 72986 74454
rect 73222 74218 108986 74454
rect 109222 74218 144986 74454
rect 145222 74218 180986 74454
rect 181222 74218 216986 74454
rect 217222 74218 252986 74454
rect 253222 74218 288986 74454
rect 289222 74218 324986 74454
rect 325222 74218 360986 74454
rect 361222 74218 396986 74454
rect 397222 74218 432986 74454
rect 433222 74218 468986 74454
rect 469222 74218 504986 74454
rect 505222 74218 540986 74454
rect 541222 74218 576986 74454
rect 577222 74218 585502 74454
rect 585738 74218 586860 74454
rect -2936 74134 586860 74218
rect -2936 73898 -1814 74134
rect -1578 73898 986 74134
rect 1222 73898 36986 74134
rect 37222 73898 72986 74134
rect 73222 73898 108986 74134
rect 109222 73898 144986 74134
rect 145222 73898 180986 74134
rect 181222 73898 216986 74134
rect 217222 73898 252986 74134
rect 253222 73898 288986 74134
rect 289222 73898 324986 74134
rect 325222 73898 360986 74134
rect 361222 73898 396986 74134
rect 397222 73898 432986 74134
rect 433222 73898 468986 74134
rect 469222 73898 504986 74134
rect 505222 73898 540986 74134
rect 541222 73898 576986 74134
rect 577222 73898 585502 74134
rect 585738 73898 586860 74134
rect -2936 73876 586860 73898
rect -1996 73874 -1396 73876
rect 804 73874 1404 73876
rect 36804 73874 37404 73876
rect 72804 73874 73404 73876
rect 108804 73874 109404 73876
rect 144804 73874 145404 73876
rect 180804 73874 181404 73876
rect 216804 73874 217404 73876
rect 252804 73874 253404 73876
rect 288804 73874 289404 73876
rect 324804 73874 325404 73876
rect 360804 73874 361404 73876
rect 396804 73874 397404 73876
rect 432804 73874 433404 73876
rect 468804 73874 469404 73876
rect 504804 73874 505404 73876
rect 540804 73874 541404 73876
rect 576804 73874 577404 73876
rect 585320 73874 585920 73876
rect -8576 67276 -7976 67278
rect 29604 67276 30204 67278
rect 65604 67276 66204 67278
rect 101604 67276 102204 67278
rect 137604 67276 138204 67278
rect 173604 67276 174204 67278
rect 209604 67276 210204 67278
rect 245604 67276 246204 67278
rect 281604 67276 282204 67278
rect 317604 67276 318204 67278
rect 353604 67276 354204 67278
rect 389604 67276 390204 67278
rect 425604 67276 426204 67278
rect 461604 67276 462204 67278
rect 497604 67276 498204 67278
rect 533604 67276 534204 67278
rect 569604 67276 570204 67278
rect 591900 67276 592500 67278
rect -8576 67254 592500 67276
rect -8576 67018 -8394 67254
rect -8158 67018 29786 67254
rect 30022 67018 65786 67254
rect 66022 67018 101786 67254
rect 102022 67018 137786 67254
rect 138022 67018 173786 67254
rect 174022 67018 209786 67254
rect 210022 67018 245786 67254
rect 246022 67018 281786 67254
rect 282022 67018 317786 67254
rect 318022 67018 353786 67254
rect 354022 67018 389786 67254
rect 390022 67018 425786 67254
rect 426022 67018 461786 67254
rect 462022 67018 497786 67254
rect 498022 67018 533786 67254
rect 534022 67018 569786 67254
rect 570022 67018 592082 67254
rect 592318 67018 592500 67254
rect -8576 66934 592500 67018
rect -8576 66698 -8394 66934
rect -8158 66698 29786 66934
rect 30022 66698 65786 66934
rect 66022 66698 101786 66934
rect 102022 66698 137786 66934
rect 138022 66698 173786 66934
rect 174022 66698 209786 66934
rect 210022 66698 245786 66934
rect 246022 66698 281786 66934
rect 282022 66698 317786 66934
rect 318022 66698 353786 66934
rect 354022 66698 389786 66934
rect 390022 66698 425786 66934
rect 426022 66698 461786 66934
rect 462022 66698 497786 66934
rect 498022 66698 533786 66934
rect 534022 66698 569786 66934
rect 570022 66698 592082 66934
rect 592318 66698 592500 66934
rect -8576 66676 592500 66698
rect -8576 66674 -7976 66676
rect 29604 66674 30204 66676
rect 65604 66674 66204 66676
rect 101604 66674 102204 66676
rect 137604 66674 138204 66676
rect 173604 66674 174204 66676
rect 209604 66674 210204 66676
rect 245604 66674 246204 66676
rect 281604 66674 282204 66676
rect 317604 66674 318204 66676
rect 353604 66674 354204 66676
rect 389604 66674 390204 66676
rect 425604 66674 426204 66676
rect 461604 66674 462204 66676
rect 497604 66674 498204 66676
rect 533604 66674 534204 66676
rect 569604 66674 570204 66676
rect 591900 66674 592500 66676
rect -6696 63676 -6096 63678
rect 26004 63676 26604 63678
rect 62004 63676 62604 63678
rect 98004 63676 98604 63678
rect 134004 63676 134604 63678
rect 170004 63676 170604 63678
rect 206004 63676 206604 63678
rect 242004 63676 242604 63678
rect 278004 63676 278604 63678
rect 314004 63676 314604 63678
rect 350004 63676 350604 63678
rect 386004 63676 386604 63678
rect 422004 63676 422604 63678
rect 458004 63676 458604 63678
rect 494004 63676 494604 63678
rect 530004 63676 530604 63678
rect 566004 63676 566604 63678
rect 590020 63676 590620 63678
rect -6696 63654 590620 63676
rect -6696 63418 -6514 63654
rect -6278 63418 26186 63654
rect 26422 63418 62186 63654
rect 62422 63418 98186 63654
rect 98422 63418 134186 63654
rect 134422 63418 170186 63654
rect 170422 63418 206186 63654
rect 206422 63418 242186 63654
rect 242422 63418 278186 63654
rect 278422 63418 314186 63654
rect 314422 63418 350186 63654
rect 350422 63418 386186 63654
rect 386422 63418 422186 63654
rect 422422 63418 458186 63654
rect 458422 63418 494186 63654
rect 494422 63418 530186 63654
rect 530422 63418 566186 63654
rect 566422 63418 590202 63654
rect 590438 63418 590620 63654
rect -6696 63334 590620 63418
rect -6696 63098 -6514 63334
rect -6278 63098 26186 63334
rect 26422 63098 62186 63334
rect 62422 63098 98186 63334
rect 98422 63098 134186 63334
rect 134422 63098 170186 63334
rect 170422 63098 206186 63334
rect 206422 63098 242186 63334
rect 242422 63098 278186 63334
rect 278422 63098 314186 63334
rect 314422 63098 350186 63334
rect 350422 63098 386186 63334
rect 386422 63098 422186 63334
rect 422422 63098 458186 63334
rect 458422 63098 494186 63334
rect 494422 63098 530186 63334
rect 530422 63098 566186 63334
rect 566422 63098 590202 63334
rect 590438 63098 590620 63334
rect -6696 63076 590620 63098
rect -6696 63074 -6096 63076
rect 26004 63074 26604 63076
rect 62004 63074 62604 63076
rect 98004 63074 98604 63076
rect 134004 63074 134604 63076
rect 170004 63074 170604 63076
rect 206004 63074 206604 63076
rect 242004 63074 242604 63076
rect 278004 63074 278604 63076
rect 314004 63074 314604 63076
rect 350004 63074 350604 63076
rect 386004 63074 386604 63076
rect 422004 63074 422604 63076
rect 458004 63074 458604 63076
rect 494004 63074 494604 63076
rect 530004 63074 530604 63076
rect 566004 63074 566604 63076
rect 590020 63074 590620 63076
rect -4816 60076 -4216 60078
rect 22404 60076 23004 60078
rect 58404 60076 59004 60078
rect 94404 60076 95004 60078
rect 130404 60076 131004 60078
rect 166404 60076 167004 60078
rect 202404 60076 203004 60078
rect 238404 60076 239004 60078
rect 274404 60076 275004 60078
rect 310404 60076 311004 60078
rect 346404 60076 347004 60078
rect 382404 60076 383004 60078
rect 418404 60076 419004 60078
rect 454404 60076 455004 60078
rect 490404 60076 491004 60078
rect 526404 60076 527004 60078
rect 562404 60076 563004 60078
rect 588140 60076 588740 60078
rect -4816 60054 588740 60076
rect -4816 59818 -4634 60054
rect -4398 59818 22586 60054
rect 22822 59818 58586 60054
rect 58822 59818 94586 60054
rect 94822 59818 130586 60054
rect 130822 59818 166586 60054
rect 166822 59818 202586 60054
rect 202822 59818 238586 60054
rect 238822 59818 274586 60054
rect 274822 59818 310586 60054
rect 310822 59818 346586 60054
rect 346822 59818 382586 60054
rect 382822 59818 418586 60054
rect 418822 59818 454586 60054
rect 454822 59818 490586 60054
rect 490822 59818 526586 60054
rect 526822 59818 562586 60054
rect 562822 59818 588322 60054
rect 588558 59818 588740 60054
rect -4816 59734 588740 59818
rect -4816 59498 -4634 59734
rect -4398 59498 22586 59734
rect 22822 59498 58586 59734
rect 58822 59498 94586 59734
rect 94822 59498 130586 59734
rect 130822 59498 166586 59734
rect 166822 59498 202586 59734
rect 202822 59498 238586 59734
rect 238822 59498 274586 59734
rect 274822 59498 310586 59734
rect 310822 59498 346586 59734
rect 346822 59498 382586 59734
rect 382822 59498 418586 59734
rect 418822 59498 454586 59734
rect 454822 59498 490586 59734
rect 490822 59498 526586 59734
rect 526822 59498 562586 59734
rect 562822 59498 588322 59734
rect 588558 59498 588740 59734
rect -4816 59476 588740 59498
rect -4816 59474 -4216 59476
rect 22404 59474 23004 59476
rect 58404 59474 59004 59476
rect 94404 59474 95004 59476
rect 130404 59474 131004 59476
rect 166404 59474 167004 59476
rect 202404 59474 203004 59476
rect 238404 59474 239004 59476
rect 274404 59474 275004 59476
rect 310404 59474 311004 59476
rect 346404 59474 347004 59476
rect 382404 59474 383004 59476
rect 418404 59474 419004 59476
rect 454404 59474 455004 59476
rect 490404 59474 491004 59476
rect 526404 59474 527004 59476
rect 562404 59474 563004 59476
rect 588140 59474 588740 59476
rect -2936 56476 -2336 56478
rect 18804 56476 19404 56478
rect 54804 56476 55404 56478
rect 90804 56476 91404 56478
rect 126804 56476 127404 56478
rect 162804 56476 163404 56478
rect 198804 56476 199404 56478
rect 234804 56476 235404 56478
rect 270804 56476 271404 56478
rect 306804 56476 307404 56478
rect 342804 56476 343404 56478
rect 378804 56476 379404 56478
rect 414804 56476 415404 56478
rect 450804 56476 451404 56478
rect 486804 56476 487404 56478
rect 522804 56476 523404 56478
rect 558804 56476 559404 56478
rect 586260 56476 586860 56478
rect -2936 56454 586860 56476
rect -2936 56218 -2754 56454
rect -2518 56218 18986 56454
rect 19222 56218 54986 56454
rect 55222 56218 90986 56454
rect 91222 56218 126986 56454
rect 127222 56218 162986 56454
rect 163222 56218 198986 56454
rect 199222 56218 234986 56454
rect 235222 56218 270986 56454
rect 271222 56218 306986 56454
rect 307222 56218 342986 56454
rect 343222 56218 378986 56454
rect 379222 56218 414986 56454
rect 415222 56218 450986 56454
rect 451222 56218 486986 56454
rect 487222 56218 522986 56454
rect 523222 56218 558986 56454
rect 559222 56218 586442 56454
rect 586678 56218 586860 56454
rect -2936 56134 586860 56218
rect -2936 55898 -2754 56134
rect -2518 55898 18986 56134
rect 19222 55898 54986 56134
rect 55222 55898 90986 56134
rect 91222 55898 126986 56134
rect 127222 55898 162986 56134
rect 163222 55898 198986 56134
rect 199222 55898 234986 56134
rect 235222 55898 270986 56134
rect 271222 55898 306986 56134
rect 307222 55898 342986 56134
rect 343222 55898 378986 56134
rect 379222 55898 414986 56134
rect 415222 55898 450986 56134
rect 451222 55898 486986 56134
rect 487222 55898 522986 56134
rect 523222 55898 558986 56134
rect 559222 55898 586442 56134
rect 586678 55898 586860 56134
rect -2936 55876 586860 55898
rect -2936 55874 -2336 55876
rect 18804 55874 19404 55876
rect 54804 55874 55404 55876
rect 90804 55874 91404 55876
rect 126804 55874 127404 55876
rect 162804 55874 163404 55876
rect 198804 55874 199404 55876
rect 234804 55874 235404 55876
rect 270804 55874 271404 55876
rect 306804 55874 307404 55876
rect 342804 55874 343404 55876
rect 378804 55874 379404 55876
rect 414804 55874 415404 55876
rect 450804 55874 451404 55876
rect 486804 55874 487404 55876
rect 522804 55874 523404 55876
rect 558804 55874 559404 55876
rect 586260 55874 586860 55876
rect -7636 49276 -7036 49278
rect 11604 49276 12204 49278
rect 47604 49276 48204 49278
rect 83604 49276 84204 49278
rect 119604 49276 120204 49278
rect 155604 49276 156204 49278
rect 191604 49276 192204 49278
rect 227604 49276 228204 49278
rect 263604 49276 264204 49278
rect 299604 49276 300204 49278
rect 335604 49276 336204 49278
rect 371604 49276 372204 49278
rect 407604 49276 408204 49278
rect 443604 49276 444204 49278
rect 479604 49276 480204 49278
rect 515604 49276 516204 49278
rect 551604 49276 552204 49278
rect 590960 49276 591560 49278
rect -8576 49254 592500 49276
rect -8576 49018 -7454 49254
rect -7218 49018 11786 49254
rect 12022 49018 47786 49254
rect 48022 49018 83786 49254
rect 84022 49018 119786 49254
rect 120022 49018 155786 49254
rect 156022 49018 191786 49254
rect 192022 49018 227786 49254
rect 228022 49018 263786 49254
rect 264022 49018 299786 49254
rect 300022 49018 335786 49254
rect 336022 49018 371786 49254
rect 372022 49018 407786 49254
rect 408022 49018 443786 49254
rect 444022 49018 479786 49254
rect 480022 49018 515786 49254
rect 516022 49018 551786 49254
rect 552022 49018 591142 49254
rect 591378 49018 592500 49254
rect -8576 48934 592500 49018
rect -8576 48698 -7454 48934
rect -7218 48698 11786 48934
rect 12022 48698 47786 48934
rect 48022 48698 83786 48934
rect 84022 48698 119786 48934
rect 120022 48698 155786 48934
rect 156022 48698 191786 48934
rect 192022 48698 227786 48934
rect 228022 48698 263786 48934
rect 264022 48698 299786 48934
rect 300022 48698 335786 48934
rect 336022 48698 371786 48934
rect 372022 48698 407786 48934
rect 408022 48698 443786 48934
rect 444022 48698 479786 48934
rect 480022 48698 515786 48934
rect 516022 48698 551786 48934
rect 552022 48698 591142 48934
rect 591378 48698 592500 48934
rect -8576 48676 592500 48698
rect -7636 48674 -7036 48676
rect 11604 48674 12204 48676
rect 47604 48674 48204 48676
rect 83604 48674 84204 48676
rect 119604 48674 120204 48676
rect 155604 48674 156204 48676
rect 191604 48674 192204 48676
rect 227604 48674 228204 48676
rect 263604 48674 264204 48676
rect 299604 48674 300204 48676
rect 335604 48674 336204 48676
rect 371604 48674 372204 48676
rect 407604 48674 408204 48676
rect 443604 48674 444204 48676
rect 479604 48674 480204 48676
rect 515604 48674 516204 48676
rect 551604 48674 552204 48676
rect 590960 48674 591560 48676
rect -5756 45676 -5156 45678
rect 8004 45676 8604 45678
rect 44004 45676 44604 45678
rect 80004 45676 80604 45678
rect 116004 45676 116604 45678
rect 152004 45676 152604 45678
rect 188004 45676 188604 45678
rect 224004 45676 224604 45678
rect 260004 45676 260604 45678
rect 296004 45676 296604 45678
rect 332004 45676 332604 45678
rect 368004 45676 368604 45678
rect 404004 45676 404604 45678
rect 440004 45676 440604 45678
rect 476004 45676 476604 45678
rect 512004 45676 512604 45678
rect 548004 45676 548604 45678
rect 589080 45676 589680 45678
rect -6696 45654 590620 45676
rect -6696 45418 -5574 45654
rect -5338 45418 8186 45654
rect 8422 45418 44186 45654
rect 44422 45418 80186 45654
rect 80422 45418 116186 45654
rect 116422 45418 152186 45654
rect 152422 45418 188186 45654
rect 188422 45418 224186 45654
rect 224422 45418 260186 45654
rect 260422 45418 296186 45654
rect 296422 45418 332186 45654
rect 332422 45418 368186 45654
rect 368422 45418 404186 45654
rect 404422 45418 440186 45654
rect 440422 45418 476186 45654
rect 476422 45418 512186 45654
rect 512422 45418 548186 45654
rect 548422 45418 589262 45654
rect 589498 45418 590620 45654
rect -6696 45334 590620 45418
rect -6696 45098 -5574 45334
rect -5338 45098 8186 45334
rect 8422 45098 44186 45334
rect 44422 45098 80186 45334
rect 80422 45098 116186 45334
rect 116422 45098 152186 45334
rect 152422 45098 188186 45334
rect 188422 45098 224186 45334
rect 224422 45098 260186 45334
rect 260422 45098 296186 45334
rect 296422 45098 332186 45334
rect 332422 45098 368186 45334
rect 368422 45098 404186 45334
rect 404422 45098 440186 45334
rect 440422 45098 476186 45334
rect 476422 45098 512186 45334
rect 512422 45098 548186 45334
rect 548422 45098 589262 45334
rect 589498 45098 590620 45334
rect -6696 45076 590620 45098
rect -5756 45074 -5156 45076
rect 8004 45074 8604 45076
rect 44004 45074 44604 45076
rect 80004 45074 80604 45076
rect 116004 45074 116604 45076
rect 152004 45074 152604 45076
rect 188004 45074 188604 45076
rect 224004 45074 224604 45076
rect 260004 45074 260604 45076
rect 296004 45074 296604 45076
rect 332004 45074 332604 45076
rect 368004 45074 368604 45076
rect 404004 45074 404604 45076
rect 440004 45074 440604 45076
rect 476004 45074 476604 45076
rect 512004 45074 512604 45076
rect 548004 45074 548604 45076
rect 589080 45074 589680 45076
rect -3876 42076 -3276 42078
rect 4404 42076 5004 42078
rect 40404 42076 41004 42078
rect 76404 42076 77004 42078
rect 112404 42076 113004 42078
rect 148404 42076 149004 42078
rect 184404 42076 185004 42078
rect 220404 42076 221004 42078
rect 256404 42076 257004 42078
rect 292404 42076 293004 42078
rect 328404 42076 329004 42078
rect 364404 42076 365004 42078
rect 400404 42076 401004 42078
rect 436404 42076 437004 42078
rect 472404 42076 473004 42078
rect 508404 42076 509004 42078
rect 544404 42076 545004 42078
rect 580404 42076 581004 42078
rect 587200 42076 587800 42078
rect -4816 42054 588740 42076
rect -4816 41818 -3694 42054
rect -3458 41818 4586 42054
rect 4822 41818 40586 42054
rect 40822 41818 76586 42054
rect 76822 41818 112586 42054
rect 112822 41818 148586 42054
rect 148822 41818 184586 42054
rect 184822 41818 220586 42054
rect 220822 41818 256586 42054
rect 256822 41818 292586 42054
rect 292822 41818 328586 42054
rect 328822 41818 364586 42054
rect 364822 41818 400586 42054
rect 400822 41818 436586 42054
rect 436822 41818 472586 42054
rect 472822 41818 508586 42054
rect 508822 41818 544586 42054
rect 544822 41818 580586 42054
rect 580822 41818 587382 42054
rect 587618 41818 588740 42054
rect -4816 41734 588740 41818
rect -4816 41498 -3694 41734
rect -3458 41498 4586 41734
rect 4822 41498 40586 41734
rect 40822 41498 76586 41734
rect 76822 41498 112586 41734
rect 112822 41498 148586 41734
rect 148822 41498 184586 41734
rect 184822 41498 220586 41734
rect 220822 41498 256586 41734
rect 256822 41498 292586 41734
rect 292822 41498 328586 41734
rect 328822 41498 364586 41734
rect 364822 41498 400586 41734
rect 400822 41498 436586 41734
rect 436822 41498 472586 41734
rect 472822 41498 508586 41734
rect 508822 41498 544586 41734
rect 544822 41498 580586 41734
rect 580822 41498 587382 41734
rect 587618 41498 588740 41734
rect -4816 41476 588740 41498
rect -3876 41474 -3276 41476
rect 4404 41474 5004 41476
rect 40404 41474 41004 41476
rect 76404 41474 77004 41476
rect 112404 41474 113004 41476
rect 148404 41474 149004 41476
rect 184404 41474 185004 41476
rect 220404 41474 221004 41476
rect 256404 41474 257004 41476
rect 292404 41474 293004 41476
rect 328404 41474 329004 41476
rect 364404 41474 365004 41476
rect 400404 41474 401004 41476
rect 436404 41474 437004 41476
rect 472404 41474 473004 41476
rect 508404 41474 509004 41476
rect 544404 41474 545004 41476
rect 580404 41474 581004 41476
rect 587200 41474 587800 41476
rect -1996 38476 -1396 38478
rect 804 38476 1404 38478
rect 36804 38476 37404 38478
rect 72804 38476 73404 38478
rect 108804 38476 109404 38478
rect 144804 38476 145404 38478
rect 180804 38476 181404 38478
rect 216804 38476 217404 38478
rect 252804 38476 253404 38478
rect 288804 38476 289404 38478
rect 324804 38476 325404 38478
rect 360804 38476 361404 38478
rect 396804 38476 397404 38478
rect 432804 38476 433404 38478
rect 468804 38476 469404 38478
rect 504804 38476 505404 38478
rect 540804 38476 541404 38478
rect 576804 38476 577404 38478
rect 585320 38476 585920 38478
rect -2936 38454 586860 38476
rect -2936 38218 -1814 38454
rect -1578 38218 986 38454
rect 1222 38218 36986 38454
rect 37222 38218 72986 38454
rect 73222 38218 108986 38454
rect 109222 38218 144986 38454
rect 145222 38218 180986 38454
rect 181222 38218 216986 38454
rect 217222 38218 252986 38454
rect 253222 38218 288986 38454
rect 289222 38218 324986 38454
rect 325222 38218 360986 38454
rect 361222 38218 396986 38454
rect 397222 38218 432986 38454
rect 433222 38218 468986 38454
rect 469222 38218 504986 38454
rect 505222 38218 540986 38454
rect 541222 38218 576986 38454
rect 577222 38218 585502 38454
rect 585738 38218 586860 38454
rect -2936 38134 586860 38218
rect -2936 37898 -1814 38134
rect -1578 37898 986 38134
rect 1222 37898 36986 38134
rect 37222 37898 72986 38134
rect 73222 37898 108986 38134
rect 109222 37898 144986 38134
rect 145222 37898 180986 38134
rect 181222 37898 216986 38134
rect 217222 37898 252986 38134
rect 253222 37898 288986 38134
rect 289222 37898 324986 38134
rect 325222 37898 360986 38134
rect 361222 37898 396986 38134
rect 397222 37898 432986 38134
rect 433222 37898 468986 38134
rect 469222 37898 504986 38134
rect 505222 37898 540986 38134
rect 541222 37898 576986 38134
rect 577222 37898 585502 38134
rect 585738 37898 586860 38134
rect -2936 37876 586860 37898
rect -1996 37874 -1396 37876
rect 804 37874 1404 37876
rect 36804 37874 37404 37876
rect 72804 37874 73404 37876
rect 108804 37874 109404 37876
rect 144804 37874 145404 37876
rect 180804 37874 181404 37876
rect 216804 37874 217404 37876
rect 252804 37874 253404 37876
rect 288804 37874 289404 37876
rect 324804 37874 325404 37876
rect 360804 37874 361404 37876
rect 396804 37874 397404 37876
rect 432804 37874 433404 37876
rect 468804 37874 469404 37876
rect 504804 37874 505404 37876
rect 540804 37874 541404 37876
rect 576804 37874 577404 37876
rect 585320 37874 585920 37876
rect -8576 31276 -7976 31278
rect 29604 31276 30204 31278
rect 65604 31276 66204 31278
rect 101604 31276 102204 31278
rect 137604 31276 138204 31278
rect 173604 31276 174204 31278
rect 209604 31276 210204 31278
rect 245604 31276 246204 31278
rect 281604 31276 282204 31278
rect 317604 31276 318204 31278
rect 353604 31276 354204 31278
rect 389604 31276 390204 31278
rect 425604 31276 426204 31278
rect 461604 31276 462204 31278
rect 497604 31276 498204 31278
rect 533604 31276 534204 31278
rect 569604 31276 570204 31278
rect 591900 31276 592500 31278
rect -8576 31254 592500 31276
rect -8576 31018 -8394 31254
rect -8158 31018 29786 31254
rect 30022 31018 65786 31254
rect 66022 31018 101786 31254
rect 102022 31018 137786 31254
rect 138022 31018 173786 31254
rect 174022 31018 209786 31254
rect 210022 31018 245786 31254
rect 246022 31018 281786 31254
rect 282022 31018 317786 31254
rect 318022 31018 353786 31254
rect 354022 31018 389786 31254
rect 390022 31018 425786 31254
rect 426022 31018 461786 31254
rect 462022 31018 497786 31254
rect 498022 31018 533786 31254
rect 534022 31018 569786 31254
rect 570022 31018 592082 31254
rect 592318 31018 592500 31254
rect -8576 30934 592500 31018
rect -8576 30698 -8394 30934
rect -8158 30698 29786 30934
rect 30022 30698 65786 30934
rect 66022 30698 101786 30934
rect 102022 30698 137786 30934
rect 138022 30698 173786 30934
rect 174022 30698 209786 30934
rect 210022 30698 245786 30934
rect 246022 30698 281786 30934
rect 282022 30698 317786 30934
rect 318022 30698 353786 30934
rect 354022 30698 389786 30934
rect 390022 30698 425786 30934
rect 426022 30698 461786 30934
rect 462022 30698 497786 30934
rect 498022 30698 533786 30934
rect 534022 30698 569786 30934
rect 570022 30698 592082 30934
rect 592318 30698 592500 30934
rect -8576 30676 592500 30698
rect -8576 30674 -7976 30676
rect 29604 30674 30204 30676
rect 65604 30674 66204 30676
rect 101604 30674 102204 30676
rect 137604 30674 138204 30676
rect 173604 30674 174204 30676
rect 209604 30674 210204 30676
rect 245604 30674 246204 30676
rect 281604 30674 282204 30676
rect 317604 30674 318204 30676
rect 353604 30674 354204 30676
rect 389604 30674 390204 30676
rect 425604 30674 426204 30676
rect 461604 30674 462204 30676
rect 497604 30674 498204 30676
rect 533604 30674 534204 30676
rect 569604 30674 570204 30676
rect 591900 30674 592500 30676
rect -6696 27676 -6096 27678
rect 26004 27676 26604 27678
rect 62004 27676 62604 27678
rect 98004 27676 98604 27678
rect 134004 27676 134604 27678
rect 170004 27676 170604 27678
rect 206004 27676 206604 27678
rect 242004 27676 242604 27678
rect 278004 27676 278604 27678
rect 314004 27676 314604 27678
rect 350004 27676 350604 27678
rect 386004 27676 386604 27678
rect 422004 27676 422604 27678
rect 458004 27676 458604 27678
rect 494004 27676 494604 27678
rect 530004 27676 530604 27678
rect 566004 27676 566604 27678
rect 590020 27676 590620 27678
rect -6696 27654 590620 27676
rect -6696 27418 -6514 27654
rect -6278 27418 26186 27654
rect 26422 27418 62186 27654
rect 62422 27418 98186 27654
rect 98422 27418 134186 27654
rect 134422 27418 170186 27654
rect 170422 27418 206186 27654
rect 206422 27418 242186 27654
rect 242422 27418 278186 27654
rect 278422 27418 314186 27654
rect 314422 27418 350186 27654
rect 350422 27418 386186 27654
rect 386422 27418 422186 27654
rect 422422 27418 458186 27654
rect 458422 27418 494186 27654
rect 494422 27418 530186 27654
rect 530422 27418 566186 27654
rect 566422 27418 590202 27654
rect 590438 27418 590620 27654
rect -6696 27334 590620 27418
rect -6696 27098 -6514 27334
rect -6278 27098 26186 27334
rect 26422 27098 62186 27334
rect 62422 27098 98186 27334
rect 98422 27098 134186 27334
rect 134422 27098 170186 27334
rect 170422 27098 206186 27334
rect 206422 27098 242186 27334
rect 242422 27098 278186 27334
rect 278422 27098 314186 27334
rect 314422 27098 350186 27334
rect 350422 27098 386186 27334
rect 386422 27098 422186 27334
rect 422422 27098 458186 27334
rect 458422 27098 494186 27334
rect 494422 27098 530186 27334
rect 530422 27098 566186 27334
rect 566422 27098 590202 27334
rect 590438 27098 590620 27334
rect -6696 27076 590620 27098
rect -6696 27074 -6096 27076
rect 26004 27074 26604 27076
rect 62004 27074 62604 27076
rect 98004 27074 98604 27076
rect 134004 27074 134604 27076
rect 170004 27074 170604 27076
rect 206004 27074 206604 27076
rect 242004 27074 242604 27076
rect 278004 27074 278604 27076
rect 314004 27074 314604 27076
rect 350004 27074 350604 27076
rect 386004 27074 386604 27076
rect 422004 27074 422604 27076
rect 458004 27074 458604 27076
rect 494004 27074 494604 27076
rect 530004 27074 530604 27076
rect 566004 27074 566604 27076
rect 590020 27074 590620 27076
rect -4816 24076 -4216 24078
rect 22404 24076 23004 24078
rect 58404 24076 59004 24078
rect 94404 24076 95004 24078
rect 130404 24076 131004 24078
rect 166404 24076 167004 24078
rect 202404 24076 203004 24078
rect 238404 24076 239004 24078
rect 274404 24076 275004 24078
rect 310404 24076 311004 24078
rect 346404 24076 347004 24078
rect 382404 24076 383004 24078
rect 418404 24076 419004 24078
rect 454404 24076 455004 24078
rect 490404 24076 491004 24078
rect 526404 24076 527004 24078
rect 562404 24076 563004 24078
rect 588140 24076 588740 24078
rect -4816 24054 588740 24076
rect -4816 23818 -4634 24054
rect -4398 23818 22586 24054
rect 22822 23818 58586 24054
rect 58822 23818 94586 24054
rect 94822 23818 130586 24054
rect 130822 23818 166586 24054
rect 166822 23818 202586 24054
rect 202822 23818 238586 24054
rect 238822 23818 274586 24054
rect 274822 23818 310586 24054
rect 310822 23818 346586 24054
rect 346822 23818 382586 24054
rect 382822 23818 418586 24054
rect 418822 23818 454586 24054
rect 454822 23818 490586 24054
rect 490822 23818 526586 24054
rect 526822 23818 562586 24054
rect 562822 23818 588322 24054
rect 588558 23818 588740 24054
rect -4816 23734 588740 23818
rect -4816 23498 -4634 23734
rect -4398 23498 22586 23734
rect 22822 23498 58586 23734
rect 58822 23498 94586 23734
rect 94822 23498 130586 23734
rect 130822 23498 166586 23734
rect 166822 23498 202586 23734
rect 202822 23498 238586 23734
rect 238822 23498 274586 23734
rect 274822 23498 310586 23734
rect 310822 23498 346586 23734
rect 346822 23498 382586 23734
rect 382822 23498 418586 23734
rect 418822 23498 454586 23734
rect 454822 23498 490586 23734
rect 490822 23498 526586 23734
rect 526822 23498 562586 23734
rect 562822 23498 588322 23734
rect 588558 23498 588740 23734
rect -4816 23476 588740 23498
rect -4816 23474 -4216 23476
rect 22404 23474 23004 23476
rect 58404 23474 59004 23476
rect 94404 23474 95004 23476
rect 130404 23474 131004 23476
rect 166404 23474 167004 23476
rect 202404 23474 203004 23476
rect 238404 23474 239004 23476
rect 274404 23474 275004 23476
rect 310404 23474 311004 23476
rect 346404 23474 347004 23476
rect 382404 23474 383004 23476
rect 418404 23474 419004 23476
rect 454404 23474 455004 23476
rect 490404 23474 491004 23476
rect 526404 23474 527004 23476
rect 562404 23474 563004 23476
rect 588140 23474 588740 23476
rect -2936 20476 -2336 20478
rect 18804 20476 19404 20478
rect 54804 20476 55404 20478
rect 90804 20476 91404 20478
rect 126804 20476 127404 20478
rect 162804 20476 163404 20478
rect 198804 20476 199404 20478
rect 234804 20476 235404 20478
rect 270804 20476 271404 20478
rect 306804 20476 307404 20478
rect 342804 20476 343404 20478
rect 378804 20476 379404 20478
rect 414804 20476 415404 20478
rect 450804 20476 451404 20478
rect 486804 20476 487404 20478
rect 522804 20476 523404 20478
rect 558804 20476 559404 20478
rect 586260 20476 586860 20478
rect -2936 20454 586860 20476
rect -2936 20218 -2754 20454
rect -2518 20218 18986 20454
rect 19222 20218 54986 20454
rect 55222 20218 90986 20454
rect 91222 20218 126986 20454
rect 127222 20218 162986 20454
rect 163222 20218 198986 20454
rect 199222 20218 234986 20454
rect 235222 20218 270986 20454
rect 271222 20218 306986 20454
rect 307222 20218 342986 20454
rect 343222 20218 378986 20454
rect 379222 20218 414986 20454
rect 415222 20218 450986 20454
rect 451222 20218 486986 20454
rect 487222 20218 522986 20454
rect 523222 20218 558986 20454
rect 559222 20218 586442 20454
rect 586678 20218 586860 20454
rect -2936 20134 586860 20218
rect -2936 19898 -2754 20134
rect -2518 19898 18986 20134
rect 19222 19898 54986 20134
rect 55222 19898 90986 20134
rect 91222 19898 126986 20134
rect 127222 19898 162986 20134
rect 163222 19898 198986 20134
rect 199222 19898 234986 20134
rect 235222 19898 270986 20134
rect 271222 19898 306986 20134
rect 307222 19898 342986 20134
rect 343222 19898 378986 20134
rect 379222 19898 414986 20134
rect 415222 19898 450986 20134
rect 451222 19898 486986 20134
rect 487222 19898 522986 20134
rect 523222 19898 558986 20134
rect 559222 19898 586442 20134
rect 586678 19898 586860 20134
rect -2936 19876 586860 19898
rect -2936 19874 -2336 19876
rect 18804 19874 19404 19876
rect 54804 19874 55404 19876
rect 90804 19874 91404 19876
rect 126804 19874 127404 19876
rect 162804 19874 163404 19876
rect 198804 19874 199404 19876
rect 234804 19874 235404 19876
rect 270804 19874 271404 19876
rect 306804 19874 307404 19876
rect 342804 19874 343404 19876
rect 378804 19874 379404 19876
rect 414804 19874 415404 19876
rect 450804 19874 451404 19876
rect 486804 19874 487404 19876
rect 522804 19874 523404 19876
rect 558804 19874 559404 19876
rect 586260 19874 586860 19876
rect -7636 13276 -7036 13278
rect 11604 13276 12204 13278
rect 47604 13276 48204 13278
rect 83604 13276 84204 13278
rect 119604 13276 120204 13278
rect 155604 13276 156204 13278
rect 191604 13276 192204 13278
rect 227604 13276 228204 13278
rect 263604 13276 264204 13278
rect 299604 13276 300204 13278
rect 335604 13276 336204 13278
rect 371604 13276 372204 13278
rect 407604 13276 408204 13278
rect 443604 13276 444204 13278
rect 479604 13276 480204 13278
rect 515604 13276 516204 13278
rect 551604 13276 552204 13278
rect 590960 13276 591560 13278
rect -8576 13254 592500 13276
rect -8576 13018 -7454 13254
rect -7218 13018 11786 13254
rect 12022 13018 47786 13254
rect 48022 13018 83786 13254
rect 84022 13018 119786 13254
rect 120022 13018 155786 13254
rect 156022 13018 191786 13254
rect 192022 13018 227786 13254
rect 228022 13018 263786 13254
rect 264022 13018 299786 13254
rect 300022 13018 335786 13254
rect 336022 13018 371786 13254
rect 372022 13018 407786 13254
rect 408022 13018 443786 13254
rect 444022 13018 479786 13254
rect 480022 13018 515786 13254
rect 516022 13018 551786 13254
rect 552022 13018 591142 13254
rect 591378 13018 592500 13254
rect -8576 12934 592500 13018
rect -8576 12698 -7454 12934
rect -7218 12698 11786 12934
rect 12022 12698 47786 12934
rect 48022 12698 83786 12934
rect 84022 12698 119786 12934
rect 120022 12698 155786 12934
rect 156022 12698 191786 12934
rect 192022 12698 227786 12934
rect 228022 12698 263786 12934
rect 264022 12698 299786 12934
rect 300022 12698 335786 12934
rect 336022 12698 371786 12934
rect 372022 12698 407786 12934
rect 408022 12698 443786 12934
rect 444022 12698 479786 12934
rect 480022 12698 515786 12934
rect 516022 12698 551786 12934
rect 552022 12698 591142 12934
rect 591378 12698 592500 12934
rect -8576 12676 592500 12698
rect -7636 12674 -7036 12676
rect 11604 12674 12204 12676
rect 47604 12674 48204 12676
rect 83604 12674 84204 12676
rect 119604 12674 120204 12676
rect 155604 12674 156204 12676
rect 191604 12674 192204 12676
rect 227604 12674 228204 12676
rect 263604 12674 264204 12676
rect 299604 12674 300204 12676
rect 335604 12674 336204 12676
rect 371604 12674 372204 12676
rect 407604 12674 408204 12676
rect 443604 12674 444204 12676
rect 479604 12674 480204 12676
rect 515604 12674 516204 12676
rect 551604 12674 552204 12676
rect 590960 12674 591560 12676
rect -5756 9676 -5156 9678
rect 8004 9676 8604 9678
rect 44004 9676 44604 9678
rect 80004 9676 80604 9678
rect 116004 9676 116604 9678
rect 152004 9676 152604 9678
rect 188004 9676 188604 9678
rect 224004 9676 224604 9678
rect 260004 9676 260604 9678
rect 296004 9676 296604 9678
rect 332004 9676 332604 9678
rect 368004 9676 368604 9678
rect 404004 9676 404604 9678
rect 440004 9676 440604 9678
rect 476004 9676 476604 9678
rect 512004 9676 512604 9678
rect 548004 9676 548604 9678
rect 589080 9676 589680 9678
rect -6696 9654 590620 9676
rect -6696 9418 -5574 9654
rect -5338 9418 8186 9654
rect 8422 9418 44186 9654
rect 44422 9418 80186 9654
rect 80422 9418 116186 9654
rect 116422 9418 152186 9654
rect 152422 9418 188186 9654
rect 188422 9418 224186 9654
rect 224422 9418 260186 9654
rect 260422 9418 296186 9654
rect 296422 9418 332186 9654
rect 332422 9418 368186 9654
rect 368422 9418 404186 9654
rect 404422 9418 440186 9654
rect 440422 9418 476186 9654
rect 476422 9418 512186 9654
rect 512422 9418 548186 9654
rect 548422 9418 589262 9654
rect 589498 9418 590620 9654
rect -6696 9334 590620 9418
rect -6696 9098 -5574 9334
rect -5338 9098 8186 9334
rect 8422 9098 44186 9334
rect 44422 9098 80186 9334
rect 80422 9098 116186 9334
rect 116422 9098 152186 9334
rect 152422 9098 188186 9334
rect 188422 9098 224186 9334
rect 224422 9098 260186 9334
rect 260422 9098 296186 9334
rect 296422 9098 332186 9334
rect 332422 9098 368186 9334
rect 368422 9098 404186 9334
rect 404422 9098 440186 9334
rect 440422 9098 476186 9334
rect 476422 9098 512186 9334
rect 512422 9098 548186 9334
rect 548422 9098 589262 9334
rect 589498 9098 590620 9334
rect -6696 9076 590620 9098
rect -5756 9074 -5156 9076
rect 8004 9074 8604 9076
rect 44004 9074 44604 9076
rect 80004 9074 80604 9076
rect 116004 9074 116604 9076
rect 152004 9074 152604 9076
rect 188004 9074 188604 9076
rect 224004 9074 224604 9076
rect 260004 9074 260604 9076
rect 296004 9074 296604 9076
rect 332004 9074 332604 9076
rect 368004 9074 368604 9076
rect 404004 9074 404604 9076
rect 440004 9074 440604 9076
rect 476004 9074 476604 9076
rect 512004 9074 512604 9076
rect 548004 9074 548604 9076
rect 589080 9074 589680 9076
rect -3876 6076 -3276 6078
rect 4404 6076 5004 6078
rect 40404 6076 41004 6078
rect 76404 6076 77004 6078
rect 112404 6076 113004 6078
rect 148404 6076 149004 6078
rect 184404 6076 185004 6078
rect 220404 6076 221004 6078
rect 256404 6076 257004 6078
rect 292404 6076 293004 6078
rect 328404 6076 329004 6078
rect 364404 6076 365004 6078
rect 400404 6076 401004 6078
rect 436404 6076 437004 6078
rect 472404 6076 473004 6078
rect 508404 6076 509004 6078
rect 544404 6076 545004 6078
rect 580404 6076 581004 6078
rect 587200 6076 587800 6078
rect -4816 6054 588740 6076
rect -4816 5818 -3694 6054
rect -3458 5818 4586 6054
rect 4822 5818 40586 6054
rect 40822 5818 76586 6054
rect 76822 5818 112586 6054
rect 112822 5818 148586 6054
rect 148822 5818 184586 6054
rect 184822 5818 220586 6054
rect 220822 5818 256586 6054
rect 256822 5818 292586 6054
rect 292822 5818 328586 6054
rect 328822 5818 364586 6054
rect 364822 5818 400586 6054
rect 400822 5818 436586 6054
rect 436822 5818 472586 6054
rect 472822 5818 508586 6054
rect 508822 5818 544586 6054
rect 544822 5818 580586 6054
rect 580822 5818 587382 6054
rect 587618 5818 588740 6054
rect -4816 5734 588740 5818
rect -4816 5498 -3694 5734
rect -3458 5498 4586 5734
rect 4822 5498 40586 5734
rect 40822 5498 76586 5734
rect 76822 5498 112586 5734
rect 112822 5498 148586 5734
rect 148822 5498 184586 5734
rect 184822 5498 220586 5734
rect 220822 5498 256586 5734
rect 256822 5498 292586 5734
rect 292822 5498 328586 5734
rect 328822 5498 364586 5734
rect 364822 5498 400586 5734
rect 400822 5498 436586 5734
rect 436822 5498 472586 5734
rect 472822 5498 508586 5734
rect 508822 5498 544586 5734
rect 544822 5498 580586 5734
rect 580822 5498 587382 5734
rect 587618 5498 588740 5734
rect -4816 5476 588740 5498
rect -3876 5474 -3276 5476
rect 4404 5474 5004 5476
rect 40404 5474 41004 5476
rect 76404 5474 77004 5476
rect 112404 5474 113004 5476
rect 148404 5474 149004 5476
rect 184404 5474 185004 5476
rect 220404 5474 221004 5476
rect 256404 5474 257004 5476
rect 292404 5474 293004 5476
rect 328404 5474 329004 5476
rect 364404 5474 365004 5476
rect 400404 5474 401004 5476
rect 436404 5474 437004 5476
rect 472404 5474 473004 5476
rect 508404 5474 509004 5476
rect 544404 5474 545004 5476
rect 580404 5474 581004 5476
rect 587200 5474 587800 5476
rect -1996 2476 -1396 2478
rect 804 2476 1404 2478
rect 36804 2476 37404 2478
rect 72804 2476 73404 2478
rect 108804 2476 109404 2478
rect 144804 2476 145404 2478
rect 180804 2476 181404 2478
rect 216804 2476 217404 2478
rect 252804 2476 253404 2478
rect 288804 2476 289404 2478
rect 324804 2476 325404 2478
rect 360804 2476 361404 2478
rect 396804 2476 397404 2478
rect 432804 2476 433404 2478
rect 468804 2476 469404 2478
rect 504804 2476 505404 2478
rect 540804 2476 541404 2478
rect 576804 2476 577404 2478
rect 585320 2476 585920 2478
rect -2936 2454 586860 2476
rect -2936 2218 -1814 2454
rect -1578 2218 986 2454
rect 1222 2218 36986 2454
rect 37222 2218 72986 2454
rect 73222 2218 108986 2454
rect 109222 2218 144986 2454
rect 145222 2218 180986 2454
rect 181222 2218 216986 2454
rect 217222 2218 252986 2454
rect 253222 2218 288986 2454
rect 289222 2218 324986 2454
rect 325222 2218 360986 2454
rect 361222 2218 396986 2454
rect 397222 2218 432986 2454
rect 433222 2218 468986 2454
rect 469222 2218 504986 2454
rect 505222 2218 540986 2454
rect 541222 2218 576986 2454
rect 577222 2218 585502 2454
rect 585738 2218 586860 2454
rect -2936 2134 586860 2218
rect -2936 1898 -1814 2134
rect -1578 1898 986 2134
rect 1222 1898 36986 2134
rect 37222 1898 72986 2134
rect 73222 1898 108986 2134
rect 109222 1898 144986 2134
rect 145222 1898 180986 2134
rect 181222 1898 216986 2134
rect 217222 1898 252986 2134
rect 253222 1898 288986 2134
rect 289222 1898 324986 2134
rect 325222 1898 360986 2134
rect 361222 1898 396986 2134
rect 397222 1898 432986 2134
rect 433222 1898 468986 2134
rect 469222 1898 504986 2134
rect 505222 1898 540986 2134
rect 541222 1898 576986 2134
rect 577222 1898 585502 2134
rect 585738 1898 586860 2134
rect -2936 1876 586860 1898
rect -1996 1874 -1396 1876
rect 804 1874 1404 1876
rect 36804 1874 37404 1876
rect 72804 1874 73404 1876
rect 108804 1874 109404 1876
rect 144804 1874 145404 1876
rect 180804 1874 181404 1876
rect 216804 1874 217404 1876
rect 252804 1874 253404 1876
rect 288804 1874 289404 1876
rect 324804 1874 325404 1876
rect 360804 1874 361404 1876
rect 396804 1874 397404 1876
rect 432804 1874 433404 1876
rect 468804 1874 469404 1876
rect 504804 1874 505404 1876
rect 540804 1874 541404 1876
rect 576804 1874 577404 1876
rect 585320 1874 585920 1876
rect -1996 -324 -1396 -322
rect 804 -324 1404 -322
rect 36804 -324 37404 -322
rect 72804 -324 73404 -322
rect 108804 -324 109404 -322
rect 144804 -324 145404 -322
rect 180804 -324 181404 -322
rect 216804 -324 217404 -322
rect 252804 -324 253404 -322
rect 288804 -324 289404 -322
rect 324804 -324 325404 -322
rect 360804 -324 361404 -322
rect 396804 -324 397404 -322
rect 432804 -324 433404 -322
rect 468804 -324 469404 -322
rect 504804 -324 505404 -322
rect 540804 -324 541404 -322
rect 576804 -324 577404 -322
rect 585320 -324 585920 -322
rect -1996 -346 585920 -324
rect -1996 -582 -1814 -346
rect -1578 -582 986 -346
rect 1222 -582 36986 -346
rect 37222 -582 72986 -346
rect 73222 -582 108986 -346
rect 109222 -582 144986 -346
rect 145222 -582 180986 -346
rect 181222 -582 216986 -346
rect 217222 -582 252986 -346
rect 253222 -582 288986 -346
rect 289222 -582 324986 -346
rect 325222 -582 360986 -346
rect 361222 -582 396986 -346
rect 397222 -582 432986 -346
rect 433222 -582 468986 -346
rect 469222 -582 504986 -346
rect 505222 -582 540986 -346
rect 541222 -582 576986 -346
rect 577222 -582 585502 -346
rect 585738 -582 585920 -346
rect -1996 -666 585920 -582
rect -1996 -902 -1814 -666
rect -1578 -902 986 -666
rect 1222 -902 36986 -666
rect 37222 -902 72986 -666
rect 73222 -902 108986 -666
rect 109222 -902 144986 -666
rect 145222 -902 180986 -666
rect 181222 -902 216986 -666
rect 217222 -902 252986 -666
rect 253222 -902 288986 -666
rect 289222 -902 324986 -666
rect 325222 -902 360986 -666
rect 361222 -902 396986 -666
rect 397222 -902 432986 -666
rect 433222 -902 468986 -666
rect 469222 -902 504986 -666
rect 505222 -902 540986 -666
rect 541222 -902 576986 -666
rect 577222 -902 585502 -666
rect 585738 -902 585920 -666
rect -1996 -924 585920 -902
rect -1996 -926 -1396 -924
rect 804 -926 1404 -924
rect 36804 -926 37404 -924
rect 72804 -926 73404 -924
rect 108804 -926 109404 -924
rect 144804 -926 145404 -924
rect 180804 -926 181404 -924
rect 216804 -926 217404 -924
rect 252804 -926 253404 -924
rect 288804 -926 289404 -924
rect 324804 -926 325404 -924
rect 360804 -926 361404 -924
rect 396804 -926 397404 -924
rect 432804 -926 433404 -924
rect 468804 -926 469404 -924
rect 504804 -926 505404 -924
rect 540804 -926 541404 -924
rect 576804 -926 577404 -924
rect 585320 -926 585920 -924
rect -2936 -1264 -2336 -1262
rect 18804 -1264 19404 -1262
rect 54804 -1264 55404 -1262
rect 90804 -1264 91404 -1262
rect 126804 -1264 127404 -1262
rect 162804 -1264 163404 -1262
rect 198804 -1264 199404 -1262
rect 234804 -1264 235404 -1262
rect 270804 -1264 271404 -1262
rect 306804 -1264 307404 -1262
rect 342804 -1264 343404 -1262
rect 378804 -1264 379404 -1262
rect 414804 -1264 415404 -1262
rect 450804 -1264 451404 -1262
rect 486804 -1264 487404 -1262
rect 522804 -1264 523404 -1262
rect 558804 -1264 559404 -1262
rect 586260 -1264 586860 -1262
rect -2936 -1286 586860 -1264
rect -2936 -1522 -2754 -1286
rect -2518 -1522 18986 -1286
rect 19222 -1522 54986 -1286
rect 55222 -1522 90986 -1286
rect 91222 -1522 126986 -1286
rect 127222 -1522 162986 -1286
rect 163222 -1522 198986 -1286
rect 199222 -1522 234986 -1286
rect 235222 -1522 270986 -1286
rect 271222 -1522 306986 -1286
rect 307222 -1522 342986 -1286
rect 343222 -1522 378986 -1286
rect 379222 -1522 414986 -1286
rect 415222 -1522 450986 -1286
rect 451222 -1522 486986 -1286
rect 487222 -1522 522986 -1286
rect 523222 -1522 558986 -1286
rect 559222 -1522 586442 -1286
rect 586678 -1522 586860 -1286
rect -2936 -1606 586860 -1522
rect -2936 -1842 -2754 -1606
rect -2518 -1842 18986 -1606
rect 19222 -1842 54986 -1606
rect 55222 -1842 90986 -1606
rect 91222 -1842 126986 -1606
rect 127222 -1842 162986 -1606
rect 163222 -1842 198986 -1606
rect 199222 -1842 234986 -1606
rect 235222 -1842 270986 -1606
rect 271222 -1842 306986 -1606
rect 307222 -1842 342986 -1606
rect 343222 -1842 378986 -1606
rect 379222 -1842 414986 -1606
rect 415222 -1842 450986 -1606
rect 451222 -1842 486986 -1606
rect 487222 -1842 522986 -1606
rect 523222 -1842 558986 -1606
rect 559222 -1842 586442 -1606
rect 586678 -1842 586860 -1606
rect -2936 -1864 586860 -1842
rect -2936 -1866 -2336 -1864
rect 18804 -1866 19404 -1864
rect 54804 -1866 55404 -1864
rect 90804 -1866 91404 -1864
rect 126804 -1866 127404 -1864
rect 162804 -1866 163404 -1864
rect 198804 -1866 199404 -1864
rect 234804 -1866 235404 -1864
rect 270804 -1866 271404 -1864
rect 306804 -1866 307404 -1864
rect 342804 -1866 343404 -1864
rect 378804 -1866 379404 -1864
rect 414804 -1866 415404 -1864
rect 450804 -1866 451404 -1864
rect 486804 -1866 487404 -1864
rect 522804 -1866 523404 -1864
rect 558804 -1866 559404 -1864
rect 586260 -1866 586860 -1864
rect -3876 -2204 -3276 -2202
rect 4404 -2204 5004 -2202
rect 40404 -2204 41004 -2202
rect 76404 -2204 77004 -2202
rect 112404 -2204 113004 -2202
rect 148404 -2204 149004 -2202
rect 184404 -2204 185004 -2202
rect 220404 -2204 221004 -2202
rect 256404 -2204 257004 -2202
rect 292404 -2204 293004 -2202
rect 328404 -2204 329004 -2202
rect 364404 -2204 365004 -2202
rect 400404 -2204 401004 -2202
rect 436404 -2204 437004 -2202
rect 472404 -2204 473004 -2202
rect 508404 -2204 509004 -2202
rect 544404 -2204 545004 -2202
rect 580404 -2204 581004 -2202
rect 587200 -2204 587800 -2202
rect -3876 -2226 587800 -2204
rect -3876 -2462 -3694 -2226
rect -3458 -2462 4586 -2226
rect 4822 -2462 40586 -2226
rect 40822 -2462 76586 -2226
rect 76822 -2462 112586 -2226
rect 112822 -2462 148586 -2226
rect 148822 -2462 184586 -2226
rect 184822 -2462 220586 -2226
rect 220822 -2462 256586 -2226
rect 256822 -2462 292586 -2226
rect 292822 -2462 328586 -2226
rect 328822 -2462 364586 -2226
rect 364822 -2462 400586 -2226
rect 400822 -2462 436586 -2226
rect 436822 -2462 472586 -2226
rect 472822 -2462 508586 -2226
rect 508822 -2462 544586 -2226
rect 544822 -2462 580586 -2226
rect 580822 -2462 587382 -2226
rect 587618 -2462 587800 -2226
rect -3876 -2546 587800 -2462
rect -3876 -2782 -3694 -2546
rect -3458 -2782 4586 -2546
rect 4822 -2782 40586 -2546
rect 40822 -2782 76586 -2546
rect 76822 -2782 112586 -2546
rect 112822 -2782 148586 -2546
rect 148822 -2782 184586 -2546
rect 184822 -2782 220586 -2546
rect 220822 -2782 256586 -2546
rect 256822 -2782 292586 -2546
rect 292822 -2782 328586 -2546
rect 328822 -2782 364586 -2546
rect 364822 -2782 400586 -2546
rect 400822 -2782 436586 -2546
rect 436822 -2782 472586 -2546
rect 472822 -2782 508586 -2546
rect 508822 -2782 544586 -2546
rect 544822 -2782 580586 -2546
rect 580822 -2782 587382 -2546
rect 587618 -2782 587800 -2546
rect -3876 -2804 587800 -2782
rect -3876 -2806 -3276 -2804
rect 4404 -2806 5004 -2804
rect 40404 -2806 41004 -2804
rect 76404 -2806 77004 -2804
rect 112404 -2806 113004 -2804
rect 148404 -2806 149004 -2804
rect 184404 -2806 185004 -2804
rect 220404 -2806 221004 -2804
rect 256404 -2806 257004 -2804
rect 292404 -2806 293004 -2804
rect 328404 -2806 329004 -2804
rect 364404 -2806 365004 -2804
rect 400404 -2806 401004 -2804
rect 436404 -2806 437004 -2804
rect 472404 -2806 473004 -2804
rect 508404 -2806 509004 -2804
rect 544404 -2806 545004 -2804
rect 580404 -2806 581004 -2804
rect 587200 -2806 587800 -2804
rect -4816 -3144 -4216 -3142
rect 22404 -3144 23004 -3142
rect 58404 -3144 59004 -3142
rect 94404 -3144 95004 -3142
rect 130404 -3144 131004 -3142
rect 166404 -3144 167004 -3142
rect 202404 -3144 203004 -3142
rect 238404 -3144 239004 -3142
rect 274404 -3144 275004 -3142
rect 310404 -3144 311004 -3142
rect 346404 -3144 347004 -3142
rect 382404 -3144 383004 -3142
rect 418404 -3144 419004 -3142
rect 454404 -3144 455004 -3142
rect 490404 -3144 491004 -3142
rect 526404 -3144 527004 -3142
rect 562404 -3144 563004 -3142
rect 588140 -3144 588740 -3142
rect -4816 -3166 588740 -3144
rect -4816 -3402 -4634 -3166
rect -4398 -3402 22586 -3166
rect 22822 -3402 58586 -3166
rect 58822 -3402 94586 -3166
rect 94822 -3402 130586 -3166
rect 130822 -3402 166586 -3166
rect 166822 -3402 202586 -3166
rect 202822 -3402 238586 -3166
rect 238822 -3402 274586 -3166
rect 274822 -3402 310586 -3166
rect 310822 -3402 346586 -3166
rect 346822 -3402 382586 -3166
rect 382822 -3402 418586 -3166
rect 418822 -3402 454586 -3166
rect 454822 -3402 490586 -3166
rect 490822 -3402 526586 -3166
rect 526822 -3402 562586 -3166
rect 562822 -3402 588322 -3166
rect 588558 -3402 588740 -3166
rect -4816 -3486 588740 -3402
rect -4816 -3722 -4634 -3486
rect -4398 -3722 22586 -3486
rect 22822 -3722 58586 -3486
rect 58822 -3722 94586 -3486
rect 94822 -3722 130586 -3486
rect 130822 -3722 166586 -3486
rect 166822 -3722 202586 -3486
rect 202822 -3722 238586 -3486
rect 238822 -3722 274586 -3486
rect 274822 -3722 310586 -3486
rect 310822 -3722 346586 -3486
rect 346822 -3722 382586 -3486
rect 382822 -3722 418586 -3486
rect 418822 -3722 454586 -3486
rect 454822 -3722 490586 -3486
rect 490822 -3722 526586 -3486
rect 526822 -3722 562586 -3486
rect 562822 -3722 588322 -3486
rect 588558 -3722 588740 -3486
rect -4816 -3744 588740 -3722
rect -4816 -3746 -4216 -3744
rect 22404 -3746 23004 -3744
rect 58404 -3746 59004 -3744
rect 94404 -3746 95004 -3744
rect 130404 -3746 131004 -3744
rect 166404 -3746 167004 -3744
rect 202404 -3746 203004 -3744
rect 238404 -3746 239004 -3744
rect 274404 -3746 275004 -3744
rect 310404 -3746 311004 -3744
rect 346404 -3746 347004 -3744
rect 382404 -3746 383004 -3744
rect 418404 -3746 419004 -3744
rect 454404 -3746 455004 -3744
rect 490404 -3746 491004 -3744
rect 526404 -3746 527004 -3744
rect 562404 -3746 563004 -3744
rect 588140 -3746 588740 -3744
rect -5756 -4084 -5156 -4082
rect 8004 -4084 8604 -4082
rect 44004 -4084 44604 -4082
rect 80004 -4084 80604 -4082
rect 116004 -4084 116604 -4082
rect 152004 -4084 152604 -4082
rect 188004 -4084 188604 -4082
rect 224004 -4084 224604 -4082
rect 260004 -4084 260604 -4082
rect 296004 -4084 296604 -4082
rect 332004 -4084 332604 -4082
rect 368004 -4084 368604 -4082
rect 404004 -4084 404604 -4082
rect 440004 -4084 440604 -4082
rect 476004 -4084 476604 -4082
rect 512004 -4084 512604 -4082
rect 548004 -4084 548604 -4082
rect 589080 -4084 589680 -4082
rect -5756 -4106 589680 -4084
rect -5756 -4342 -5574 -4106
rect -5338 -4342 8186 -4106
rect 8422 -4342 44186 -4106
rect 44422 -4342 80186 -4106
rect 80422 -4342 116186 -4106
rect 116422 -4342 152186 -4106
rect 152422 -4342 188186 -4106
rect 188422 -4342 224186 -4106
rect 224422 -4342 260186 -4106
rect 260422 -4342 296186 -4106
rect 296422 -4342 332186 -4106
rect 332422 -4342 368186 -4106
rect 368422 -4342 404186 -4106
rect 404422 -4342 440186 -4106
rect 440422 -4342 476186 -4106
rect 476422 -4342 512186 -4106
rect 512422 -4342 548186 -4106
rect 548422 -4342 589262 -4106
rect 589498 -4342 589680 -4106
rect -5756 -4426 589680 -4342
rect -5756 -4662 -5574 -4426
rect -5338 -4662 8186 -4426
rect 8422 -4662 44186 -4426
rect 44422 -4662 80186 -4426
rect 80422 -4662 116186 -4426
rect 116422 -4662 152186 -4426
rect 152422 -4662 188186 -4426
rect 188422 -4662 224186 -4426
rect 224422 -4662 260186 -4426
rect 260422 -4662 296186 -4426
rect 296422 -4662 332186 -4426
rect 332422 -4662 368186 -4426
rect 368422 -4662 404186 -4426
rect 404422 -4662 440186 -4426
rect 440422 -4662 476186 -4426
rect 476422 -4662 512186 -4426
rect 512422 -4662 548186 -4426
rect 548422 -4662 589262 -4426
rect 589498 -4662 589680 -4426
rect -5756 -4684 589680 -4662
rect -5756 -4686 -5156 -4684
rect 8004 -4686 8604 -4684
rect 44004 -4686 44604 -4684
rect 80004 -4686 80604 -4684
rect 116004 -4686 116604 -4684
rect 152004 -4686 152604 -4684
rect 188004 -4686 188604 -4684
rect 224004 -4686 224604 -4684
rect 260004 -4686 260604 -4684
rect 296004 -4686 296604 -4684
rect 332004 -4686 332604 -4684
rect 368004 -4686 368604 -4684
rect 404004 -4686 404604 -4684
rect 440004 -4686 440604 -4684
rect 476004 -4686 476604 -4684
rect 512004 -4686 512604 -4684
rect 548004 -4686 548604 -4684
rect 589080 -4686 589680 -4684
rect -6696 -5024 -6096 -5022
rect 26004 -5024 26604 -5022
rect 62004 -5024 62604 -5022
rect 98004 -5024 98604 -5022
rect 134004 -5024 134604 -5022
rect 170004 -5024 170604 -5022
rect 206004 -5024 206604 -5022
rect 242004 -5024 242604 -5022
rect 278004 -5024 278604 -5022
rect 314004 -5024 314604 -5022
rect 350004 -5024 350604 -5022
rect 386004 -5024 386604 -5022
rect 422004 -5024 422604 -5022
rect 458004 -5024 458604 -5022
rect 494004 -5024 494604 -5022
rect 530004 -5024 530604 -5022
rect 566004 -5024 566604 -5022
rect 590020 -5024 590620 -5022
rect -6696 -5046 590620 -5024
rect -6696 -5282 -6514 -5046
rect -6278 -5282 26186 -5046
rect 26422 -5282 62186 -5046
rect 62422 -5282 98186 -5046
rect 98422 -5282 134186 -5046
rect 134422 -5282 170186 -5046
rect 170422 -5282 206186 -5046
rect 206422 -5282 242186 -5046
rect 242422 -5282 278186 -5046
rect 278422 -5282 314186 -5046
rect 314422 -5282 350186 -5046
rect 350422 -5282 386186 -5046
rect 386422 -5282 422186 -5046
rect 422422 -5282 458186 -5046
rect 458422 -5282 494186 -5046
rect 494422 -5282 530186 -5046
rect 530422 -5282 566186 -5046
rect 566422 -5282 590202 -5046
rect 590438 -5282 590620 -5046
rect -6696 -5366 590620 -5282
rect -6696 -5602 -6514 -5366
rect -6278 -5602 26186 -5366
rect 26422 -5602 62186 -5366
rect 62422 -5602 98186 -5366
rect 98422 -5602 134186 -5366
rect 134422 -5602 170186 -5366
rect 170422 -5602 206186 -5366
rect 206422 -5602 242186 -5366
rect 242422 -5602 278186 -5366
rect 278422 -5602 314186 -5366
rect 314422 -5602 350186 -5366
rect 350422 -5602 386186 -5366
rect 386422 -5602 422186 -5366
rect 422422 -5602 458186 -5366
rect 458422 -5602 494186 -5366
rect 494422 -5602 530186 -5366
rect 530422 -5602 566186 -5366
rect 566422 -5602 590202 -5366
rect 590438 -5602 590620 -5366
rect -6696 -5624 590620 -5602
rect -6696 -5626 -6096 -5624
rect 26004 -5626 26604 -5624
rect 62004 -5626 62604 -5624
rect 98004 -5626 98604 -5624
rect 134004 -5626 134604 -5624
rect 170004 -5626 170604 -5624
rect 206004 -5626 206604 -5624
rect 242004 -5626 242604 -5624
rect 278004 -5626 278604 -5624
rect 314004 -5626 314604 -5624
rect 350004 -5626 350604 -5624
rect 386004 -5626 386604 -5624
rect 422004 -5626 422604 -5624
rect 458004 -5626 458604 -5624
rect 494004 -5626 494604 -5624
rect 530004 -5626 530604 -5624
rect 566004 -5626 566604 -5624
rect 590020 -5626 590620 -5624
rect -7636 -5964 -7036 -5962
rect 11604 -5964 12204 -5962
rect 47604 -5964 48204 -5962
rect 83604 -5964 84204 -5962
rect 119604 -5964 120204 -5962
rect 155604 -5964 156204 -5962
rect 191604 -5964 192204 -5962
rect 227604 -5964 228204 -5962
rect 263604 -5964 264204 -5962
rect 299604 -5964 300204 -5962
rect 335604 -5964 336204 -5962
rect 371604 -5964 372204 -5962
rect 407604 -5964 408204 -5962
rect 443604 -5964 444204 -5962
rect 479604 -5964 480204 -5962
rect 515604 -5964 516204 -5962
rect 551604 -5964 552204 -5962
rect 590960 -5964 591560 -5962
rect -7636 -5986 591560 -5964
rect -7636 -6222 -7454 -5986
rect -7218 -6222 11786 -5986
rect 12022 -6222 47786 -5986
rect 48022 -6222 83786 -5986
rect 84022 -6222 119786 -5986
rect 120022 -6222 155786 -5986
rect 156022 -6222 191786 -5986
rect 192022 -6222 227786 -5986
rect 228022 -6222 263786 -5986
rect 264022 -6222 299786 -5986
rect 300022 -6222 335786 -5986
rect 336022 -6222 371786 -5986
rect 372022 -6222 407786 -5986
rect 408022 -6222 443786 -5986
rect 444022 -6222 479786 -5986
rect 480022 -6222 515786 -5986
rect 516022 -6222 551786 -5986
rect 552022 -6222 591142 -5986
rect 591378 -6222 591560 -5986
rect -7636 -6306 591560 -6222
rect -7636 -6542 -7454 -6306
rect -7218 -6542 11786 -6306
rect 12022 -6542 47786 -6306
rect 48022 -6542 83786 -6306
rect 84022 -6542 119786 -6306
rect 120022 -6542 155786 -6306
rect 156022 -6542 191786 -6306
rect 192022 -6542 227786 -6306
rect 228022 -6542 263786 -6306
rect 264022 -6542 299786 -6306
rect 300022 -6542 335786 -6306
rect 336022 -6542 371786 -6306
rect 372022 -6542 407786 -6306
rect 408022 -6542 443786 -6306
rect 444022 -6542 479786 -6306
rect 480022 -6542 515786 -6306
rect 516022 -6542 551786 -6306
rect 552022 -6542 591142 -6306
rect 591378 -6542 591560 -6306
rect -7636 -6564 591560 -6542
rect -7636 -6566 -7036 -6564
rect 11604 -6566 12204 -6564
rect 47604 -6566 48204 -6564
rect 83604 -6566 84204 -6564
rect 119604 -6566 120204 -6564
rect 155604 -6566 156204 -6564
rect 191604 -6566 192204 -6564
rect 227604 -6566 228204 -6564
rect 263604 -6566 264204 -6564
rect 299604 -6566 300204 -6564
rect 335604 -6566 336204 -6564
rect 371604 -6566 372204 -6564
rect 407604 -6566 408204 -6564
rect 443604 -6566 444204 -6564
rect 479604 -6566 480204 -6564
rect 515604 -6566 516204 -6564
rect 551604 -6566 552204 -6564
rect 590960 -6566 591560 -6564
rect -8576 -6904 -7976 -6902
rect 29604 -6904 30204 -6902
rect 65604 -6904 66204 -6902
rect 101604 -6904 102204 -6902
rect 137604 -6904 138204 -6902
rect 173604 -6904 174204 -6902
rect 209604 -6904 210204 -6902
rect 245604 -6904 246204 -6902
rect 281604 -6904 282204 -6902
rect 317604 -6904 318204 -6902
rect 353604 -6904 354204 -6902
rect 389604 -6904 390204 -6902
rect 425604 -6904 426204 -6902
rect 461604 -6904 462204 -6902
rect 497604 -6904 498204 -6902
rect 533604 -6904 534204 -6902
rect 569604 -6904 570204 -6902
rect 591900 -6904 592500 -6902
rect -8576 -6926 592500 -6904
rect -8576 -7162 -8394 -6926
rect -8158 -7162 29786 -6926
rect 30022 -7162 65786 -6926
rect 66022 -7162 101786 -6926
rect 102022 -7162 137786 -6926
rect 138022 -7162 173786 -6926
rect 174022 -7162 209786 -6926
rect 210022 -7162 245786 -6926
rect 246022 -7162 281786 -6926
rect 282022 -7162 317786 -6926
rect 318022 -7162 353786 -6926
rect 354022 -7162 389786 -6926
rect 390022 -7162 425786 -6926
rect 426022 -7162 461786 -6926
rect 462022 -7162 497786 -6926
rect 498022 -7162 533786 -6926
rect 534022 -7162 569786 -6926
rect 570022 -7162 592082 -6926
rect 592318 -7162 592500 -6926
rect -8576 -7246 592500 -7162
rect -8576 -7482 -8394 -7246
rect -8158 -7482 29786 -7246
rect 30022 -7482 65786 -7246
rect 66022 -7482 101786 -7246
rect 102022 -7482 137786 -7246
rect 138022 -7482 173786 -7246
rect 174022 -7482 209786 -7246
rect 210022 -7482 245786 -7246
rect 246022 -7482 281786 -7246
rect 282022 -7482 317786 -7246
rect 318022 -7482 353786 -7246
rect 354022 -7482 389786 -7246
rect 390022 -7482 425786 -7246
rect 426022 -7482 461786 -7246
rect 462022 -7482 497786 -7246
rect 498022 -7482 533786 -7246
rect 534022 -7482 569786 -7246
rect 570022 -7482 592082 -7246
rect 592318 -7482 592500 -7246
rect -8576 -7504 592500 -7482
rect -8576 -7506 -7976 -7504
rect 29604 -7506 30204 -7504
rect 65604 -7506 66204 -7504
rect 101604 -7506 102204 -7504
rect 137604 -7506 138204 -7504
rect 173604 -7506 174204 -7504
rect 209604 -7506 210204 -7504
rect 245604 -7506 246204 -7504
rect 281604 -7506 282204 -7504
rect 317604 -7506 318204 -7504
rect 353604 -7506 354204 -7504
rect 389604 -7506 390204 -7504
rect 425604 -7506 426204 -7504
rect 461604 -7506 462204 -7504
rect 497604 -7506 498204 -7504
rect 533604 -7506 534204 -7504
rect 569604 -7506 570204 -7504
rect 591900 -7506 592500 -7504
use MM2hdmi  proj_7
timestamp 1608040051
transform 1 0 200000 0 1 520000
box 0 0 20000 40000
use challenge  proj_6
timestamp 1608040051
transform 1 0 480000 0 1 520000
box 0 0 31344 34764
use watch_hhmm  proj_5
timestamp 1608040051
transform 1 0 360000 0 1 360000
box 0 0 31275 33419
use asic_freq  proj_4
timestamp 1608040051
transform 1 0 300000 0 1 500000
box 0 0 77867 80011
use spinet5  proj_3
timestamp 1608040051
transform 1 0 200000 0 1 340000
box 0 0 66678 68822
use vga_clock  proj_2
timestamp 1608040051
transform 1 0 460000 0 1 340000
box 0 0 45405 47549
use ws2812  proj_1
timestamp 1608040051
transform 1 0 72000 0 1 340000
box 0 0 54206 56350
use seven_segment_seconds  proj_0
timestamp 1608040051
transform 1 0 86000 0 1 520000
box 0 0 29760 31904
use multi_project_harness  mprj
timestamp 1608040051
transform 1 0 134000 0 1 120000
box 0 0 300000 80000
<< labels >>
rlabel metal3 s 583520 5796 584960 6036 6 analog_io[0]
port 0 nsew default bidirectional
rlabel metal3 s 583520 474996 584960 475236 6 analog_io[10]
port 1 nsew default bidirectional
rlabel metal3 s 583520 521916 584960 522156 6 analog_io[11]
port 2 nsew default bidirectional
rlabel metal3 s 583520 568836 584960 569076 6 analog_io[12]
port 3 nsew default bidirectional
rlabel metal3 s 583520 615756 584960 615996 6 analog_io[13]
port 4 nsew default bidirectional
rlabel metal3 s 583520 662676 584960 662916 6 analog_io[14]
port 5 nsew default bidirectional
rlabel metal2 s 575818 703520 575930 704960 6 analog_io[15]
port 6 nsew default bidirectional
rlabel metal2 s 510958 703520 511070 704960 6 analog_io[16]
port 7 nsew default bidirectional
rlabel metal2 s 446098 703520 446210 704960 6 analog_io[17]
port 8 nsew default bidirectional
rlabel metal2 s 381146 703520 381258 704960 6 analog_io[18]
port 9 nsew default bidirectional
rlabel metal2 s 316286 703520 316398 704960 6 analog_io[19]
port 10 nsew default bidirectional
rlabel metal3 s 583520 52716 584960 52956 6 analog_io[1]
port 11 nsew default bidirectional
rlabel metal2 s 251426 703520 251538 704960 6 analog_io[20]
port 12 nsew default bidirectional
rlabel metal2 s 186474 703520 186586 704960 6 analog_io[21]
port 13 nsew default bidirectional
rlabel metal2 s 121614 703520 121726 704960 6 analog_io[22]
port 14 nsew default bidirectional
rlabel metal2 s 56754 703520 56866 704960 6 analog_io[23]
port 15 nsew default bidirectional
rlabel metal3 s -960 696540 480 696780 4 analog_io[24]
port 16 nsew default bidirectional
rlabel metal3 s -960 639012 480 639252 4 analog_io[25]
port 17 nsew default bidirectional
rlabel metal3 s -960 581620 480 581860 4 analog_io[26]
port 18 nsew default bidirectional
rlabel metal3 s -960 524092 480 524332 4 analog_io[27]
port 19 nsew default bidirectional
rlabel metal3 s -960 466700 480 466940 4 analog_io[28]
port 20 nsew default bidirectional
rlabel metal3 s -960 409172 480 409412 4 analog_io[29]
port 21 nsew default bidirectional
rlabel metal3 s 583520 99636 584960 99876 6 analog_io[2]
port 22 nsew default bidirectional
rlabel metal3 s -960 351780 480 352020 4 analog_io[30]
port 23 nsew default bidirectional
rlabel metal3 s 583520 146556 584960 146796 6 analog_io[3]
port 24 nsew default bidirectional
rlabel metal3 s 583520 193476 584960 193716 6 analog_io[4]
port 25 nsew default bidirectional
rlabel metal3 s 583520 240396 584960 240636 6 analog_io[5]
port 26 nsew default bidirectional
rlabel metal3 s 583520 287316 584960 287556 6 analog_io[6]
port 27 nsew default bidirectional
rlabel metal3 s 583520 334236 584960 334476 6 analog_io[7]
port 28 nsew default bidirectional
rlabel metal3 s 583520 381156 584960 381396 6 analog_io[8]
port 29 nsew default bidirectional
rlabel metal3 s 583520 428076 584960 428316 6 analog_io[9]
port 30 nsew default bidirectional
rlabel metal3 s 583520 17492 584960 17732 6 io_in[0]
port 31 nsew default input
rlabel metal3 s 583520 486692 584960 486932 6 io_in[10]
port 32 nsew default input
rlabel metal3 s 583520 533748 584960 533988 6 io_in[11]
port 33 nsew default input
rlabel metal3 s 583520 580668 584960 580908 6 io_in[12]
port 34 nsew default input
rlabel metal3 s 583520 627588 584960 627828 6 io_in[13]
port 35 nsew default input
rlabel metal3 s 583520 674508 584960 674748 6 io_in[14]
port 36 nsew default input
rlabel metal2 s 559626 703520 559738 704960 6 io_in[15]
port 37 nsew default input
rlabel metal2 s 494766 703520 494878 704960 6 io_in[16]
port 38 nsew default input
rlabel metal2 s 429814 703520 429926 704960 6 io_in[17]
port 39 nsew default input
rlabel metal2 s 364954 703520 365066 704960 6 io_in[18]
port 40 nsew default input
rlabel metal2 s 300094 703520 300206 704960 6 io_in[19]
port 41 nsew default input
rlabel metal3 s 583520 64412 584960 64652 6 io_in[1]
port 42 nsew default input
rlabel metal2 s 235142 703520 235254 704960 6 io_in[20]
port 43 nsew default input
rlabel metal2 s 170282 703520 170394 704960 6 io_in[21]
port 44 nsew default input
rlabel metal2 s 105422 703520 105534 704960 6 io_in[22]
port 45 nsew default input
rlabel metal2 s 40470 703520 40582 704960 6 io_in[23]
port 46 nsew default input
rlabel metal3 s -960 682124 480 682364 4 io_in[24]
port 47 nsew default input
rlabel metal3 s -960 624732 480 624972 4 io_in[25]
port 48 nsew default input
rlabel metal3 s -960 567204 480 567444 4 io_in[26]
port 49 nsew default input
rlabel metal3 s -960 509812 480 510052 4 io_in[27]
port 50 nsew default input
rlabel metal3 s -960 452284 480 452524 4 io_in[28]
port 51 nsew default input
rlabel metal3 s -960 394892 480 395132 4 io_in[29]
port 52 nsew default input
rlabel metal3 s 583520 111332 584960 111572 6 io_in[2]
port 53 nsew default input
rlabel metal3 s -960 337364 480 337604 4 io_in[30]
port 54 nsew default input
rlabel metal3 s -960 294252 480 294492 4 io_in[31]
port 55 nsew default input
rlabel metal3 s -960 251140 480 251380 4 io_in[32]
port 56 nsew default input
rlabel metal3 s -960 208028 480 208268 4 io_in[33]
port 57 nsew default input
rlabel metal3 s -960 164916 480 165156 4 io_in[34]
port 58 nsew default input
rlabel metal3 s -960 121940 480 122180 4 io_in[35]
port 59 nsew default input
rlabel metal3 s -960 78828 480 79068 4 io_in[36]
port 60 nsew default input
rlabel metal3 s -960 35716 480 35956 4 io_in[37]
port 61 nsew default input
rlabel metal3 s 583520 158252 584960 158492 6 io_in[3]
port 62 nsew default input
rlabel metal3 s 583520 205172 584960 205412 6 io_in[4]
port 63 nsew default input
rlabel metal3 s 583520 252092 584960 252332 6 io_in[5]
port 64 nsew default input
rlabel metal3 s 583520 299012 584960 299252 6 io_in[6]
port 65 nsew default input
rlabel metal3 s 583520 345932 584960 346172 6 io_in[7]
port 66 nsew default input
rlabel metal3 s 583520 392852 584960 393092 6 io_in[8]
port 67 nsew default input
rlabel metal3 s 583520 439772 584960 440012 6 io_in[9]
port 68 nsew default input
rlabel metal3 s 583520 40884 584960 41124 6 io_oeb[0]
port 69 nsew default tristate
rlabel metal3 s 583520 510220 584960 510460 6 io_oeb[10]
port 70 nsew default tristate
rlabel metal3 s 583520 557140 584960 557380 6 io_oeb[11]
port 71 nsew default tristate
rlabel metal3 s 583520 604060 584960 604300 6 io_oeb[12]
port 72 nsew default tristate
rlabel metal3 s 583520 650980 584960 651220 6 io_oeb[13]
port 73 nsew default tristate
rlabel metal3 s 583520 697900 584960 698140 6 io_oeb[14]
port 74 nsew default tristate
rlabel metal2 s 527150 703520 527262 704960 6 io_oeb[15]
port 75 nsew default tristate
rlabel metal2 s 462290 703520 462402 704960 6 io_oeb[16]
port 76 nsew default tristate
rlabel metal2 s 397430 703520 397542 704960 6 io_oeb[17]
port 77 nsew default tristate
rlabel metal2 s 332478 703520 332590 704960 6 io_oeb[18]
port 78 nsew default tristate
rlabel metal2 s 267618 703520 267730 704960 6 io_oeb[19]
port 79 nsew default tristate
rlabel metal3 s 583520 87804 584960 88044 6 io_oeb[1]
port 80 nsew default tristate
rlabel metal2 s 202758 703520 202870 704960 6 io_oeb[20]
port 81 nsew default tristate
rlabel metal2 s 137806 703520 137918 704960 6 io_oeb[21]
port 82 nsew default tristate
rlabel metal2 s 72946 703520 73058 704960 6 io_oeb[22]
port 83 nsew default tristate
rlabel metal2 s 8086 703520 8198 704960 6 io_oeb[23]
port 84 nsew default tristate
rlabel metal3 s -960 653428 480 653668 4 io_oeb[24]
port 85 nsew default tristate
rlabel metal3 s -960 595900 480 596140 4 io_oeb[25]
port 86 nsew default tristate
rlabel metal3 s -960 538508 480 538748 4 io_oeb[26]
port 87 nsew default tristate
rlabel metal3 s -960 480980 480 481220 4 io_oeb[27]
port 88 nsew default tristate
rlabel metal3 s -960 423588 480 423828 4 io_oeb[28]
port 89 nsew default tristate
rlabel metal3 s -960 366060 480 366300 4 io_oeb[29]
port 90 nsew default tristate
rlabel metal3 s 583520 134724 584960 134964 6 io_oeb[2]
port 91 nsew default tristate
rlabel metal3 s -960 308668 480 308908 4 io_oeb[30]
port 92 nsew default tristate
rlabel metal3 s -960 265556 480 265796 4 io_oeb[31]
port 93 nsew default tristate
rlabel metal3 s -960 222444 480 222684 4 io_oeb[32]
port 94 nsew default tristate
rlabel metal3 s -960 179332 480 179572 4 io_oeb[33]
port 95 nsew default tristate
rlabel metal3 s -960 136220 480 136460 4 io_oeb[34]
port 96 nsew default tristate
rlabel metal3 s -960 93108 480 93348 4 io_oeb[35]
port 97 nsew default tristate
rlabel metal3 s -960 49996 480 50236 4 io_oeb[36]
port 98 nsew default tristate
rlabel metal3 s -960 7020 480 7260 4 io_oeb[37]
port 99 nsew default tristate
rlabel metal3 s 583520 181780 584960 182020 6 io_oeb[3]
port 100 nsew default tristate
rlabel metal3 s 583520 228700 584960 228940 6 io_oeb[4]
port 101 nsew default tristate
rlabel metal3 s 583520 275620 584960 275860 6 io_oeb[5]
port 102 nsew default tristate
rlabel metal3 s 583520 322540 584960 322780 6 io_oeb[6]
port 103 nsew default tristate
rlabel metal3 s 583520 369460 584960 369700 6 io_oeb[7]
port 104 nsew default tristate
rlabel metal3 s 583520 416380 584960 416620 6 io_oeb[8]
port 105 nsew default tristate
rlabel metal3 s 583520 463300 584960 463540 6 io_oeb[9]
port 106 nsew default tristate
rlabel metal3 s 583520 29188 584960 29428 6 io_out[0]
port 107 nsew default tristate
rlabel metal3 s 583520 498524 584960 498764 6 io_out[10]
port 108 nsew default tristate
rlabel metal3 s 583520 545444 584960 545684 6 io_out[11]
port 109 nsew default tristate
rlabel metal3 s 583520 592364 584960 592604 6 io_out[12]
port 110 nsew default tristate
rlabel metal3 s 583520 639284 584960 639524 6 io_out[13]
port 111 nsew default tristate
rlabel metal3 s 583520 686204 584960 686444 6 io_out[14]
port 112 nsew default tristate
rlabel metal2 s 543434 703520 543546 704960 6 io_out[15]
port 113 nsew default tristate
rlabel metal2 s 478482 703520 478594 704960 6 io_out[16]
port 114 nsew default tristate
rlabel metal2 s 413622 703520 413734 704960 6 io_out[17]
port 115 nsew default tristate
rlabel metal2 s 348762 703520 348874 704960 6 io_out[18]
port 116 nsew default tristate
rlabel metal2 s 283810 703520 283922 704960 6 io_out[19]
port 117 nsew default tristate
rlabel metal3 s 583520 76108 584960 76348 6 io_out[1]
port 118 nsew default tristate
rlabel metal2 s 218950 703520 219062 704960 6 io_out[20]
port 119 nsew default tristate
rlabel metal2 s 154090 703520 154202 704960 6 io_out[21]
port 120 nsew default tristate
rlabel metal2 s 89138 703520 89250 704960 6 io_out[22]
port 121 nsew default tristate
rlabel metal2 s 24278 703520 24390 704960 6 io_out[23]
port 122 nsew default tristate
rlabel metal3 s -960 667844 480 668084 4 io_out[24]
port 123 nsew default tristate
rlabel metal3 s -960 610316 480 610556 4 io_out[25]
port 124 nsew default tristate
rlabel metal3 s -960 552924 480 553164 4 io_out[26]
port 125 nsew default tristate
rlabel metal3 s -960 495396 480 495636 4 io_out[27]
port 126 nsew default tristate
rlabel metal3 s -960 437868 480 438108 4 io_out[28]
port 127 nsew default tristate
rlabel metal3 s -960 380476 480 380716 4 io_out[29]
port 128 nsew default tristate
rlabel metal3 s 583520 123028 584960 123268 6 io_out[2]
port 129 nsew default tristate
rlabel metal3 s -960 322948 480 323188 4 io_out[30]
port 130 nsew default tristate
rlabel metal3 s -960 279972 480 280212 4 io_out[31]
port 131 nsew default tristate
rlabel metal3 s -960 236860 480 237100 4 io_out[32]
port 132 nsew default tristate
rlabel metal3 s -960 193748 480 193988 4 io_out[33]
port 133 nsew default tristate
rlabel metal3 s -960 150636 480 150876 4 io_out[34]
port 134 nsew default tristate
rlabel metal3 s -960 107524 480 107764 4 io_out[35]
port 135 nsew default tristate
rlabel metal3 s -960 64412 480 64652 4 io_out[36]
port 136 nsew default tristate
rlabel metal3 s -960 21300 480 21540 4 io_out[37]
port 137 nsew default tristate
rlabel metal3 s 583520 169948 584960 170188 6 io_out[3]
port 138 nsew default tristate
rlabel metal3 s 583520 216868 584960 217108 6 io_out[4]
port 139 nsew default tristate
rlabel metal3 s 583520 263788 584960 264028 6 io_out[5]
port 140 nsew default tristate
rlabel metal3 s 583520 310708 584960 310948 6 io_out[6]
port 141 nsew default tristate
rlabel metal3 s 583520 357764 584960 358004 6 io_out[7]
port 142 nsew default tristate
rlabel metal3 s 583520 404684 584960 404924 6 io_out[8]
port 143 nsew default tristate
rlabel metal3 s 583520 451604 584960 451844 6 io_out[9]
port 144 nsew default tristate
rlabel metal2 s 126582 -960 126694 480 8 la_data_in[0]
port 145 nsew default input
rlabel metal2 s 483450 -960 483562 480 8 la_data_in[100]
port 146 nsew default input
rlabel metal2 s 486946 -960 487058 480 8 la_data_in[101]
port 147 nsew default input
rlabel metal2 s 490534 -960 490646 480 8 la_data_in[102]
port 148 nsew default input
rlabel metal2 s 494122 -960 494234 480 8 la_data_in[103]
port 149 nsew default input
rlabel metal2 s 497710 -960 497822 480 8 la_data_in[104]
port 150 nsew default input
rlabel metal2 s 501206 -960 501318 480 8 la_data_in[105]
port 151 nsew default input
rlabel metal2 s 504794 -960 504906 480 8 la_data_in[106]
port 152 nsew default input
rlabel metal2 s 508382 -960 508494 480 8 la_data_in[107]
port 153 nsew default input
rlabel metal2 s 511970 -960 512082 480 8 la_data_in[108]
port 154 nsew default input
rlabel metal2 s 515558 -960 515670 480 8 la_data_in[109]
port 155 nsew default input
rlabel metal2 s 162278 -960 162390 480 8 la_data_in[10]
port 156 nsew default input
rlabel metal2 s 519054 -960 519166 480 8 la_data_in[110]
port 157 nsew default input
rlabel metal2 s 522642 -960 522754 480 8 la_data_in[111]
port 158 nsew default input
rlabel metal2 s 526230 -960 526342 480 8 la_data_in[112]
port 159 nsew default input
rlabel metal2 s 529818 -960 529930 480 8 la_data_in[113]
port 160 nsew default input
rlabel metal2 s 533406 -960 533518 480 8 la_data_in[114]
port 161 nsew default input
rlabel metal2 s 536902 -960 537014 480 8 la_data_in[115]
port 162 nsew default input
rlabel metal2 s 540490 -960 540602 480 8 la_data_in[116]
port 163 nsew default input
rlabel metal2 s 544078 -960 544190 480 8 la_data_in[117]
port 164 nsew default input
rlabel metal2 s 547666 -960 547778 480 8 la_data_in[118]
port 165 nsew default input
rlabel metal2 s 551162 -960 551274 480 8 la_data_in[119]
port 166 nsew default input
rlabel metal2 s 165866 -960 165978 480 8 la_data_in[11]
port 167 nsew default input
rlabel metal2 s 554750 -960 554862 480 8 la_data_in[120]
port 168 nsew default input
rlabel metal2 s 558338 -960 558450 480 8 la_data_in[121]
port 169 nsew default input
rlabel metal2 s 561926 -960 562038 480 8 la_data_in[122]
port 170 nsew default input
rlabel metal2 s 565514 -960 565626 480 8 la_data_in[123]
port 171 nsew default input
rlabel metal2 s 569010 -960 569122 480 8 la_data_in[124]
port 172 nsew default input
rlabel metal2 s 572598 -960 572710 480 8 la_data_in[125]
port 173 nsew default input
rlabel metal2 s 576186 -960 576298 480 8 la_data_in[126]
port 174 nsew default input
rlabel metal2 s 579774 -960 579886 480 8 la_data_in[127]
port 175 nsew default input
rlabel metal2 s 169362 -960 169474 480 8 la_data_in[12]
port 176 nsew default input
rlabel metal2 s 172950 -960 173062 480 8 la_data_in[13]
port 177 nsew default input
rlabel metal2 s 176538 -960 176650 480 8 la_data_in[14]
port 178 nsew default input
rlabel metal2 s 180126 -960 180238 480 8 la_data_in[15]
port 179 nsew default input
rlabel metal2 s 183714 -960 183826 480 8 la_data_in[16]
port 180 nsew default input
rlabel metal2 s 187210 -960 187322 480 8 la_data_in[17]
port 181 nsew default input
rlabel metal2 s 190798 -960 190910 480 8 la_data_in[18]
port 182 nsew default input
rlabel metal2 s 194386 -960 194498 480 8 la_data_in[19]
port 183 nsew default input
rlabel metal2 s 130170 -960 130282 480 8 la_data_in[1]
port 184 nsew default input
rlabel metal2 s 197974 -960 198086 480 8 la_data_in[20]
port 185 nsew default input
rlabel metal2 s 201470 -960 201582 480 8 la_data_in[21]
port 186 nsew default input
rlabel metal2 s 205058 -960 205170 480 8 la_data_in[22]
port 187 nsew default input
rlabel metal2 s 208646 -960 208758 480 8 la_data_in[23]
port 188 nsew default input
rlabel metal2 s 212234 -960 212346 480 8 la_data_in[24]
port 189 nsew default input
rlabel metal2 s 215822 -960 215934 480 8 la_data_in[25]
port 190 nsew default input
rlabel metal2 s 219318 -960 219430 480 8 la_data_in[26]
port 191 nsew default input
rlabel metal2 s 222906 -960 223018 480 8 la_data_in[27]
port 192 nsew default input
rlabel metal2 s 226494 -960 226606 480 8 la_data_in[28]
port 193 nsew default input
rlabel metal2 s 230082 -960 230194 480 8 la_data_in[29]
port 194 nsew default input
rlabel metal2 s 133758 -960 133870 480 8 la_data_in[2]
port 195 nsew default input
rlabel metal2 s 233670 -960 233782 480 8 la_data_in[30]
port 196 nsew default input
rlabel metal2 s 237166 -960 237278 480 8 la_data_in[31]
port 197 nsew default input
rlabel metal2 s 240754 -960 240866 480 8 la_data_in[32]
port 198 nsew default input
rlabel metal2 s 244342 -960 244454 480 8 la_data_in[33]
port 199 nsew default input
rlabel metal2 s 247930 -960 248042 480 8 la_data_in[34]
port 200 nsew default input
rlabel metal2 s 251426 -960 251538 480 8 la_data_in[35]
port 201 nsew default input
rlabel metal2 s 255014 -960 255126 480 8 la_data_in[36]
port 202 nsew default input
rlabel metal2 s 258602 -960 258714 480 8 la_data_in[37]
port 203 nsew default input
rlabel metal2 s 262190 -960 262302 480 8 la_data_in[38]
port 204 nsew default input
rlabel metal2 s 265778 -960 265890 480 8 la_data_in[39]
port 205 nsew default input
rlabel metal2 s 137254 -960 137366 480 8 la_data_in[3]
port 206 nsew default input
rlabel metal2 s 269274 -960 269386 480 8 la_data_in[40]
port 207 nsew default input
rlabel metal2 s 272862 -960 272974 480 8 la_data_in[41]
port 208 nsew default input
rlabel metal2 s 276450 -960 276562 480 8 la_data_in[42]
port 209 nsew default input
rlabel metal2 s 280038 -960 280150 480 8 la_data_in[43]
port 210 nsew default input
rlabel metal2 s 283626 -960 283738 480 8 la_data_in[44]
port 211 nsew default input
rlabel metal2 s 287122 -960 287234 480 8 la_data_in[45]
port 212 nsew default input
rlabel metal2 s 290710 -960 290822 480 8 la_data_in[46]
port 213 nsew default input
rlabel metal2 s 294298 -960 294410 480 8 la_data_in[47]
port 214 nsew default input
rlabel metal2 s 297886 -960 297998 480 8 la_data_in[48]
port 215 nsew default input
rlabel metal2 s 301382 -960 301494 480 8 la_data_in[49]
port 216 nsew default input
rlabel metal2 s 140842 -960 140954 480 8 la_data_in[4]
port 217 nsew default input
rlabel metal2 s 304970 -960 305082 480 8 la_data_in[50]
port 218 nsew default input
rlabel metal2 s 308558 -960 308670 480 8 la_data_in[51]
port 219 nsew default input
rlabel metal2 s 312146 -960 312258 480 8 la_data_in[52]
port 220 nsew default input
rlabel metal2 s 315734 -960 315846 480 8 la_data_in[53]
port 221 nsew default input
rlabel metal2 s 319230 -960 319342 480 8 la_data_in[54]
port 222 nsew default input
rlabel metal2 s 322818 -960 322930 480 8 la_data_in[55]
port 223 nsew default input
rlabel metal2 s 326406 -960 326518 480 8 la_data_in[56]
port 224 nsew default input
rlabel metal2 s 329994 -960 330106 480 8 la_data_in[57]
port 225 nsew default input
rlabel metal2 s 333582 -960 333694 480 8 la_data_in[58]
port 226 nsew default input
rlabel metal2 s 337078 -960 337190 480 8 la_data_in[59]
port 227 nsew default input
rlabel metal2 s 144430 -960 144542 480 8 la_data_in[5]
port 228 nsew default input
rlabel metal2 s 340666 -960 340778 480 8 la_data_in[60]
port 229 nsew default input
rlabel metal2 s 344254 -960 344366 480 8 la_data_in[61]
port 230 nsew default input
rlabel metal2 s 347842 -960 347954 480 8 la_data_in[62]
port 231 nsew default input
rlabel metal2 s 351338 -960 351450 480 8 la_data_in[63]
port 232 nsew default input
rlabel metal2 s 354926 -960 355038 480 8 la_data_in[64]
port 233 nsew default input
rlabel metal2 s 358514 -960 358626 480 8 la_data_in[65]
port 234 nsew default input
rlabel metal2 s 362102 -960 362214 480 8 la_data_in[66]
port 235 nsew default input
rlabel metal2 s 365690 -960 365802 480 8 la_data_in[67]
port 236 nsew default input
rlabel metal2 s 369186 -960 369298 480 8 la_data_in[68]
port 237 nsew default input
rlabel metal2 s 372774 -960 372886 480 8 la_data_in[69]
port 238 nsew default input
rlabel metal2 s 148018 -960 148130 480 8 la_data_in[6]
port 239 nsew default input
rlabel metal2 s 376362 -960 376474 480 8 la_data_in[70]
port 240 nsew default input
rlabel metal2 s 379950 -960 380062 480 8 la_data_in[71]
port 241 nsew default input
rlabel metal2 s 383538 -960 383650 480 8 la_data_in[72]
port 242 nsew default input
rlabel metal2 s 387034 -960 387146 480 8 la_data_in[73]
port 243 nsew default input
rlabel metal2 s 390622 -960 390734 480 8 la_data_in[74]
port 244 nsew default input
rlabel metal2 s 394210 -960 394322 480 8 la_data_in[75]
port 245 nsew default input
rlabel metal2 s 397798 -960 397910 480 8 la_data_in[76]
port 246 nsew default input
rlabel metal2 s 401294 -960 401406 480 8 la_data_in[77]
port 247 nsew default input
rlabel metal2 s 404882 -960 404994 480 8 la_data_in[78]
port 248 nsew default input
rlabel metal2 s 408470 -960 408582 480 8 la_data_in[79]
port 249 nsew default input
rlabel metal2 s 151514 -960 151626 480 8 la_data_in[7]
port 250 nsew default input
rlabel metal2 s 412058 -960 412170 480 8 la_data_in[80]
port 251 nsew default input
rlabel metal2 s 415646 -960 415758 480 8 la_data_in[81]
port 252 nsew default input
rlabel metal2 s 419142 -960 419254 480 8 la_data_in[82]
port 253 nsew default input
rlabel metal2 s 422730 -960 422842 480 8 la_data_in[83]
port 254 nsew default input
rlabel metal2 s 426318 -960 426430 480 8 la_data_in[84]
port 255 nsew default input
rlabel metal2 s 429906 -960 430018 480 8 la_data_in[85]
port 256 nsew default input
rlabel metal2 s 433494 -960 433606 480 8 la_data_in[86]
port 257 nsew default input
rlabel metal2 s 436990 -960 437102 480 8 la_data_in[87]
port 258 nsew default input
rlabel metal2 s 440578 -960 440690 480 8 la_data_in[88]
port 259 nsew default input
rlabel metal2 s 444166 -960 444278 480 8 la_data_in[89]
port 260 nsew default input
rlabel metal2 s 155102 -960 155214 480 8 la_data_in[8]
port 261 nsew default input
rlabel metal2 s 447754 -960 447866 480 8 la_data_in[90]
port 262 nsew default input
rlabel metal2 s 451250 -960 451362 480 8 la_data_in[91]
port 263 nsew default input
rlabel metal2 s 454838 -960 454950 480 8 la_data_in[92]
port 264 nsew default input
rlabel metal2 s 458426 -960 458538 480 8 la_data_in[93]
port 265 nsew default input
rlabel metal2 s 462014 -960 462126 480 8 la_data_in[94]
port 266 nsew default input
rlabel metal2 s 465602 -960 465714 480 8 la_data_in[95]
port 267 nsew default input
rlabel metal2 s 469098 -960 469210 480 8 la_data_in[96]
port 268 nsew default input
rlabel metal2 s 472686 -960 472798 480 8 la_data_in[97]
port 269 nsew default input
rlabel metal2 s 476274 -960 476386 480 8 la_data_in[98]
port 270 nsew default input
rlabel metal2 s 479862 -960 479974 480 8 la_data_in[99]
port 271 nsew default input
rlabel metal2 s 158690 -960 158802 480 8 la_data_in[9]
port 272 nsew default input
rlabel metal2 s 127778 -960 127890 480 8 la_data_out[0]
port 273 nsew default tristate
rlabel metal2 s 484554 -960 484666 480 8 la_data_out[100]
port 274 nsew default tristate
rlabel metal2 s 488142 -960 488254 480 8 la_data_out[101]
port 275 nsew default tristate
rlabel metal2 s 491730 -960 491842 480 8 la_data_out[102]
port 276 nsew default tristate
rlabel metal2 s 495318 -960 495430 480 8 la_data_out[103]
port 277 nsew default tristate
rlabel metal2 s 498906 -960 499018 480 8 la_data_out[104]
port 278 nsew default tristate
rlabel metal2 s 502402 -960 502514 480 8 la_data_out[105]
port 279 nsew default tristate
rlabel metal2 s 505990 -960 506102 480 8 la_data_out[106]
port 280 nsew default tristate
rlabel metal2 s 509578 -960 509690 480 8 la_data_out[107]
port 281 nsew default tristate
rlabel metal2 s 513166 -960 513278 480 8 la_data_out[108]
port 282 nsew default tristate
rlabel metal2 s 516754 -960 516866 480 8 la_data_out[109]
port 283 nsew default tristate
rlabel metal2 s 163474 -960 163586 480 8 la_data_out[10]
port 284 nsew default tristate
rlabel metal2 s 520250 -960 520362 480 8 la_data_out[110]
port 285 nsew default tristate
rlabel metal2 s 523838 -960 523950 480 8 la_data_out[111]
port 286 nsew default tristate
rlabel metal2 s 527426 -960 527538 480 8 la_data_out[112]
port 287 nsew default tristate
rlabel metal2 s 531014 -960 531126 480 8 la_data_out[113]
port 288 nsew default tristate
rlabel metal2 s 534510 -960 534622 480 8 la_data_out[114]
port 289 nsew default tristate
rlabel metal2 s 538098 -960 538210 480 8 la_data_out[115]
port 290 nsew default tristate
rlabel metal2 s 541686 -960 541798 480 8 la_data_out[116]
port 291 nsew default tristate
rlabel metal2 s 545274 -960 545386 480 8 la_data_out[117]
port 292 nsew default tristate
rlabel metal2 s 548862 -960 548974 480 8 la_data_out[118]
port 293 nsew default tristate
rlabel metal2 s 552358 -960 552470 480 8 la_data_out[119]
port 294 nsew default tristate
rlabel metal2 s 167062 -960 167174 480 8 la_data_out[11]
port 295 nsew default tristate
rlabel metal2 s 555946 -960 556058 480 8 la_data_out[120]
port 296 nsew default tristate
rlabel metal2 s 559534 -960 559646 480 8 la_data_out[121]
port 297 nsew default tristate
rlabel metal2 s 563122 -960 563234 480 8 la_data_out[122]
port 298 nsew default tristate
rlabel metal2 s 566710 -960 566822 480 8 la_data_out[123]
port 299 nsew default tristate
rlabel metal2 s 570206 -960 570318 480 8 la_data_out[124]
port 300 nsew default tristate
rlabel metal2 s 573794 -960 573906 480 8 la_data_out[125]
port 301 nsew default tristate
rlabel metal2 s 577382 -960 577494 480 8 la_data_out[126]
port 302 nsew default tristate
rlabel metal2 s 580970 -960 581082 480 8 la_data_out[127]
port 303 nsew default tristate
rlabel metal2 s 170558 -960 170670 480 8 la_data_out[12]
port 304 nsew default tristate
rlabel metal2 s 174146 -960 174258 480 8 la_data_out[13]
port 305 nsew default tristate
rlabel metal2 s 177734 -960 177846 480 8 la_data_out[14]
port 306 nsew default tristate
rlabel metal2 s 181322 -960 181434 480 8 la_data_out[15]
port 307 nsew default tristate
rlabel metal2 s 184818 -960 184930 480 8 la_data_out[16]
port 308 nsew default tristate
rlabel metal2 s 188406 -960 188518 480 8 la_data_out[17]
port 309 nsew default tristate
rlabel metal2 s 191994 -960 192106 480 8 la_data_out[18]
port 310 nsew default tristate
rlabel metal2 s 195582 -960 195694 480 8 la_data_out[19]
port 311 nsew default tristate
rlabel metal2 s 131366 -960 131478 480 8 la_data_out[1]
port 312 nsew default tristate
rlabel metal2 s 199170 -960 199282 480 8 la_data_out[20]
port 313 nsew default tristate
rlabel metal2 s 202666 -960 202778 480 8 la_data_out[21]
port 314 nsew default tristate
rlabel metal2 s 206254 -960 206366 480 8 la_data_out[22]
port 315 nsew default tristate
rlabel metal2 s 209842 -960 209954 480 8 la_data_out[23]
port 316 nsew default tristate
rlabel metal2 s 213430 -960 213542 480 8 la_data_out[24]
port 317 nsew default tristate
rlabel metal2 s 217018 -960 217130 480 8 la_data_out[25]
port 318 nsew default tristate
rlabel metal2 s 220514 -960 220626 480 8 la_data_out[26]
port 319 nsew default tristate
rlabel metal2 s 224102 -960 224214 480 8 la_data_out[27]
port 320 nsew default tristate
rlabel metal2 s 227690 -960 227802 480 8 la_data_out[28]
port 321 nsew default tristate
rlabel metal2 s 231278 -960 231390 480 8 la_data_out[29]
port 322 nsew default tristate
rlabel metal2 s 134862 -960 134974 480 8 la_data_out[2]
port 323 nsew default tristate
rlabel metal2 s 234774 -960 234886 480 8 la_data_out[30]
port 324 nsew default tristate
rlabel metal2 s 238362 -960 238474 480 8 la_data_out[31]
port 325 nsew default tristate
rlabel metal2 s 241950 -960 242062 480 8 la_data_out[32]
port 326 nsew default tristate
rlabel metal2 s 245538 -960 245650 480 8 la_data_out[33]
port 327 nsew default tristate
rlabel metal2 s 249126 -960 249238 480 8 la_data_out[34]
port 328 nsew default tristate
rlabel metal2 s 252622 -960 252734 480 8 la_data_out[35]
port 329 nsew default tristate
rlabel metal2 s 256210 -960 256322 480 8 la_data_out[36]
port 330 nsew default tristate
rlabel metal2 s 259798 -960 259910 480 8 la_data_out[37]
port 331 nsew default tristate
rlabel metal2 s 263386 -960 263498 480 8 la_data_out[38]
port 332 nsew default tristate
rlabel metal2 s 266974 -960 267086 480 8 la_data_out[39]
port 333 nsew default tristate
rlabel metal2 s 138450 -960 138562 480 8 la_data_out[3]
port 334 nsew default tristate
rlabel metal2 s 270470 -960 270582 480 8 la_data_out[40]
port 335 nsew default tristate
rlabel metal2 s 274058 -960 274170 480 8 la_data_out[41]
port 336 nsew default tristate
rlabel metal2 s 277646 -960 277758 480 8 la_data_out[42]
port 337 nsew default tristate
rlabel metal2 s 281234 -960 281346 480 8 la_data_out[43]
port 338 nsew default tristate
rlabel metal2 s 284730 -960 284842 480 8 la_data_out[44]
port 339 nsew default tristate
rlabel metal2 s 288318 -960 288430 480 8 la_data_out[45]
port 340 nsew default tristate
rlabel metal2 s 291906 -960 292018 480 8 la_data_out[46]
port 341 nsew default tristate
rlabel metal2 s 295494 -960 295606 480 8 la_data_out[47]
port 342 nsew default tristate
rlabel metal2 s 299082 -960 299194 480 8 la_data_out[48]
port 343 nsew default tristate
rlabel metal2 s 302578 -960 302690 480 8 la_data_out[49]
port 344 nsew default tristate
rlabel metal2 s 142038 -960 142150 480 8 la_data_out[4]
port 345 nsew default tristate
rlabel metal2 s 306166 -960 306278 480 8 la_data_out[50]
port 346 nsew default tristate
rlabel metal2 s 309754 -960 309866 480 8 la_data_out[51]
port 347 nsew default tristate
rlabel metal2 s 313342 -960 313454 480 8 la_data_out[52]
port 348 nsew default tristate
rlabel metal2 s 316930 -960 317042 480 8 la_data_out[53]
port 349 nsew default tristate
rlabel metal2 s 320426 -960 320538 480 8 la_data_out[54]
port 350 nsew default tristate
rlabel metal2 s 324014 -960 324126 480 8 la_data_out[55]
port 351 nsew default tristate
rlabel metal2 s 327602 -960 327714 480 8 la_data_out[56]
port 352 nsew default tristate
rlabel metal2 s 331190 -960 331302 480 8 la_data_out[57]
port 353 nsew default tristate
rlabel metal2 s 334686 -960 334798 480 8 la_data_out[58]
port 354 nsew default tristate
rlabel metal2 s 338274 -960 338386 480 8 la_data_out[59]
port 355 nsew default tristate
rlabel metal2 s 145626 -960 145738 480 8 la_data_out[5]
port 356 nsew default tristate
rlabel metal2 s 341862 -960 341974 480 8 la_data_out[60]
port 357 nsew default tristate
rlabel metal2 s 345450 -960 345562 480 8 la_data_out[61]
port 358 nsew default tristate
rlabel metal2 s 349038 -960 349150 480 8 la_data_out[62]
port 359 nsew default tristate
rlabel metal2 s 352534 -960 352646 480 8 la_data_out[63]
port 360 nsew default tristate
rlabel metal2 s 356122 -960 356234 480 8 la_data_out[64]
port 361 nsew default tristate
rlabel metal2 s 359710 -960 359822 480 8 la_data_out[65]
port 362 nsew default tristate
rlabel metal2 s 363298 -960 363410 480 8 la_data_out[66]
port 363 nsew default tristate
rlabel metal2 s 366886 -960 366998 480 8 la_data_out[67]
port 364 nsew default tristate
rlabel metal2 s 370382 -960 370494 480 8 la_data_out[68]
port 365 nsew default tristate
rlabel metal2 s 373970 -960 374082 480 8 la_data_out[69]
port 366 nsew default tristate
rlabel metal2 s 149214 -960 149326 480 8 la_data_out[6]
port 367 nsew default tristate
rlabel metal2 s 377558 -960 377670 480 8 la_data_out[70]
port 368 nsew default tristate
rlabel metal2 s 381146 -960 381258 480 8 la_data_out[71]
port 369 nsew default tristate
rlabel metal2 s 384642 -960 384754 480 8 la_data_out[72]
port 370 nsew default tristate
rlabel metal2 s 388230 -960 388342 480 8 la_data_out[73]
port 371 nsew default tristate
rlabel metal2 s 391818 -960 391930 480 8 la_data_out[74]
port 372 nsew default tristate
rlabel metal2 s 395406 -960 395518 480 8 la_data_out[75]
port 373 nsew default tristate
rlabel metal2 s 398994 -960 399106 480 8 la_data_out[76]
port 374 nsew default tristate
rlabel metal2 s 402490 -960 402602 480 8 la_data_out[77]
port 375 nsew default tristate
rlabel metal2 s 406078 -960 406190 480 8 la_data_out[78]
port 376 nsew default tristate
rlabel metal2 s 409666 -960 409778 480 8 la_data_out[79]
port 377 nsew default tristate
rlabel metal2 s 152710 -960 152822 480 8 la_data_out[7]
port 378 nsew default tristate
rlabel metal2 s 413254 -960 413366 480 8 la_data_out[80]
port 379 nsew default tristate
rlabel metal2 s 416842 -960 416954 480 8 la_data_out[81]
port 380 nsew default tristate
rlabel metal2 s 420338 -960 420450 480 8 la_data_out[82]
port 381 nsew default tristate
rlabel metal2 s 423926 -960 424038 480 8 la_data_out[83]
port 382 nsew default tristate
rlabel metal2 s 427514 -960 427626 480 8 la_data_out[84]
port 383 nsew default tristate
rlabel metal2 s 431102 -960 431214 480 8 la_data_out[85]
port 384 nsew default tristate
rlabel metal2 s 434598 -960 434710 480 8 la_data_out[86]
port 385 nsew default tristate
rlabel metal2 s 438186 -960 438298 480 8 la_data_out[87]
port 386 nsew default tristate
rlabel metal2 s 441774 -960 441886 480 8 la_data_out[88]
port 387 nsew default tristate
rlabel metal2 s 445362 -960 445474 480 8 la_data_out[89]
port 388 nsew default tristate
rlabel metal2 s 156298 -960 156410 480 8 la_data_out[8]
port 389 nsew default tristate
rlabel metal2 s 448950 -960 449062 480 8 la_data_out[90]
port 390 nsew default tristate
rlabel metal2 s 452446 -960 452558 480 8 la_data_out[91]
port 391 nsew default tristate
rlabel metal2 s 456034 -960 456146 480 8 la_data_out[92]
port 392 nsew default tristate
rlabel metal2 s 459622 -960 459734 480 8 la_data_out[93]
port 393 nsew default tristate
rlabel metal2 s 463210 -960 463322 480 8 la_data_out[94]
port 394 nsew default tristate
rlabel metal2 s 466798 -960 466910 480 8 la_data_out[95]
port 395 nsew default tristate
rlabel metal2 s 470294 -960 470406 480 8 la_data_out[96]
port 396 nsew default tristate
rlabel metal2 s 473882 -960 473994 480 8 la_data_out[97]
port 397 nsew default tristate
rlabel metal2 s 477470 -960 477582 480 8 la_data_out[98]
port 398 nsew default tristate
rlabel metal2 s 481058 -960 481170 480 8 la_data_out[99]
port 399 nsew default tristate
rlabel metal2 s 159886 -960 159998 480 8 la_data_out[9]
port 400 nsew default tristate
rlabel metal2 s 128974 -960 129086 480 8 la_oen[0]
port 401 nsew default input
rlabel metal2 s 485750 -960 485862 480 8 la_oen[100]
port 402 nsew default input
rlabel metal2 s 489338 -960 489450 480 8 la_oen[101]
port 403 nsew default input
rlabel metal2 s 492926 -960 493038 480 8 la_oen[102]
port 404 nsew default input
rlabel metal2 s 496514 -960 496626 480 8 la_oen[103]
port 405 nsew default input
rlabel metal2 s 500102 -960 500214 480 8 la_oen[104]
port 406 nsew default input
rlabel metal2 s 503598 -960 503710 480 8 la_oen[105]
port 407 nsew default input
rlabel metal2 s 507186 -960 507298 480 8 la_oen[106]
port 408 nsew default input
rlabel metal2 s 510774 -960 510886 480 8 la_oen[107]
port 409 nsew default input
rlabel metal2 s 514362 -960 514474 480 8 la_oen[108]
port 410 nsew default input
rlabel metal2 s 517858 -960 517970 480 8 la_oen[109]
port 411 nsew default input
rlabel metal2 s 164670 -960 164782 480 8 la_oen[10]
port 412 nsew default input
rlabel metal2 s 521446 -960 521558 480 8 la_oen[110]
port 413 nsew default input
rlabel metal2 s 525034 -960 525146 480 8 la_oen[111]
port 414 nsew default input
rlabel metal2 s 528622 -960 528734 480 8 la_oen[112]
port 415 nsew default input
rlabel metal2 s 532210 -960 532322 480 8 la_oen[113]
port 416 nsew default input
rlabel metal2 s 535706 -960 535818 480 8 la_oen[114]
port 417 nsew default input
rlabel metal2 s 539294 -960 539406 480 8 la_oen[115]
port 418 nsew default input
rlabel metal2 s 542882 -960 542994 480 8 la_oen[116]
port 419 nsew default input
rlabel metal2 s 546470 -960 546582 480 8 la_oen[117]
port 420 nsew default input
rlabel metal2 s 550058 -960 550170 480 8 la_oen[118]
port 421 nsew default input
rlabel metal2 s 553554 -960 553666 480 8 la_oen[119]
port 422 nsew default input
rlabel metal2 s 168166 -960 168278 480 8 la_oen[11]
port 423 nsew default input
rlabel metal2 s 557142 -960 557254 480 8 la_oen[120]
port 424 nsew default input
rlabel metal2 s 560730 -960 560842 480 8 la_oen[121]
port 425 nsew default input
rlabel metal2 s 564318 -960 564430 480 8 la_oen[122]
port 426 nsew default input
rlabel metal2 s 567814 -960 567926 480 8 la_oen[123]
port 427 nsew default input
rlabel metal2 s 571402 -960 571514 480 8 la_oen[124]
port 428 nsew default input
rlabel metal2 s 574990 -960 575102 480 8 la_oen[125]
port 429 nsew default input
rlabel metal2 s 578578 -960 578690 480 8 la_oen[126]
port 430 nsew default input
rlabel metal2 s 582166 -960 582278 480 8 la_oen[127]
port 431 nsew default input
rlabel metal2 s 171754 -960 171866 480 8 la_oen[12]
port 432 nsew default input
rlabel metal2 s 175342 -960 175454 480 8 la_oen[13]
port 433 nsew default input
rlabel metal2 s 178930 -960 179042 480 8 la_oen[14]
port 434 nsew default input
rlabel metal2 s 182518 -960 182630 480 8 la_oen[15]
port 435 nsew default input
rlabel metal2 s 186014 -960 186126 480 8 la_oen[16]
port 436 nsew default input
rlabel metal2 s 189602 -960 189714 480 8 la_oen[17]
port 437 nsew default input
rlabel metal2 s 193190 -960 193302 480 8 la_oen[18]
port 438 nsew default input
rlabel metal2 s 196778 -960 196890 480 8 la_oen[19]
port 439 nsew default input
rlabel metal2 s 132562 -960 132674 480 8 la_oen[1]
port 440 nsew default input
rlabel metal2 s 200366 -960 200478 480 8 la_oen[20]
port 441 nsew default input
rlabel metal2 s 203862 -960 203974 480 8 la_oen[21]
port 442 nsew default input
rlabel metal2 s 207450 -960 207562 480 8 la_oen[22]
port 443 nsew default input
rlabel metal2 s 211038 -960 211150 480 8 la_oen[23]
port 444 nsew default input
rlabel metal2 s 214626 -960 214738 480 8 la_oen[24]
port 445 nsew default input
rlabel metal2 s 218122 -960 218234 480 8 la_oen[25]
port 446 nsew default input
rlabel metal2 s 221710 -960 221822 480 8 la_oen[26]
port 447 nsew default input
rlabel metal2 s 225298 -960 225410 480 8 la_oen[27]
port 448 nsew default input
rlabel metal2 s 228886 -960 228998 480 8 la_oen[28]
port 449 nsew default input
rlabel metal2 s 232474 -960 232586 480 8 la_oen[29]
port 450 nsew default input
rlabel metal2 s 136058 -960 136170 480 8 la_oen[2]
port 451 nsew default input
rlabel metal2 s 235970 -960 236082 480 8 la_oen[30]
port 452 nsew default input
rlabel metal2 s 239558 -960 239670 480 8 la_oen[31]
port 453 nsew default input
rlabel metal2 s 243146 -960 243258 480 8 la_oen[32]
port 454 nsew default input
rlabel metal2 s 246734 -960 246846 480 8 la_oen[33]
port 455 nsew default input
rlabel metal2 s 250322 -960 250434 480 8 la_oen[34]
port 456 nsew default input
rlabel metal2 s 253818 -960 253930 480 8 la_oen[35]
port 457 nsew default input
rlabel metal2 s 257406 -960 257518 480 8 la_oen[36]
port 458 nsew default input
rlabel metal2 s 260994 -960 261106 480 8 la_oen[37]
port 459 nsew default input
rlabel metal2 s 264582 -960 264694 480 8 la_oen[38]
port 460 nsew default input
rlabel metal2 s 268078 -960 268190 480 8 la_oen[39]
port 461 nsew default input
rlabel metal2 s 139646 -960 139758 480 8 la_oen[3]
port 462 nsew default input
rlabel metal2 s 271666 -960 271778 480 8 la_oen[40]
port 463 nsew default input
rlabel metal2 s 275254 -960 275366 480 8 la_oen[41]
port 464 nsew default input
rlabel metal2 s 278842 -960 278954 480 8 la_oen[42]
port 465 nsew default input
rlabel metal2 s 282430 -960 282542 480 8 la_oen[43]
port 466 nsew default input
rlabel metal2 s 285926 -960 286038 480 8 la_oen[44]
port 467 nsew default input
rlabel metal2 s 289514 -960 289626 480 8 la_oen[45]
port 468 nsew default input
rlabel metal2 s 293102 -960 293214 480 8 la_oen[46]
port 469 nsew default input
rlabel metal2 s 296690 -960 296802 480 8 la_oen[47]
port 470 nsew default input
rlabel metal2 s 300278 -960 300390 480 8 la_oen[48]
port 471 nsew default input
rlabel metal2 s 303774 -960 303886 480 8 la_oen[49]
port 472 nsew default input
rlabel metal2 s 143234 -960 143346 480 8 la_oen[4]
port 473 nsew default input
rlabel metal2 s 307362 -960 307474 480 8 la_oen[50]
port 474 nsew default input
rlabel metal2 s 310950 -960 311062 480 8 la_oen[51]
port 475 nsew default input
rlabel metal2 s 314538 -960 314650 480 8 la_oen[52]
port 476 nsew default input
rlabel metal2 s 318034 -960 318146 480 8 la_oen[53]
port 477 nsew default input
rlabel metal2 s 321622 -960 321734 480 8 la_oen[54]
port 478 nsew default input
rlabel metal2 s 325210 -960 325322 480 8 la_oen[55]
port 479 nsew default input
rlabel metal2 s 328798 -960 328910 480 8 la_oen[56]
port 480 nsew default input
rlabel metal2 s 332386 -960 332498 480 8 la_oen[57]
port 481 nsew default input
rlabel metal2 s 335882 -960 335994 480 8 la_oen[58]
port 482 nsew default input
rlabel metal2 s 339470 -960 339582 480 8 la_oen[59]
port 483 nsew default input
rlabel metal2 s 146822 -960 146934 480 8 la_oen[5]
port 484 nsew default input
rlabel metal2 s 343058 -960 343170 480 8 la_oen[60]
port 485 nsew default input
rlabel metal2 s 346646 -960 346758 480 8 la_oen[61]
port 486 nsew default input
rlabel metal2 s 350234 -960 350346 480 8 la_oen[62]
port 487 nsew default input
rlabel metal2 s 353730 -960 353842 480 8 la_oen[63]
port 488 nsew default input
rlabel metal2 s 357318 -960 357430 480 8 la_oen[64]
port 489 nsew default input
rlabel metal2 s 360906 -960 361018 480 8 la_oen[65]
port 490 nsew default input
rlabel metal2 s 364494 -960 364606 480 8 la_oen[66]
port 491 nsew default input
rlabel metal2 s 367990 -960 368102 480 8 la_oen[67]
port 492 nsew default input
rlabel metal2 s 371578 -960 371690 480 8 la_oen[68]
port 493 nsew default input
rlabel metal2 s 375166 -960 375278 480 8 la_oen[69]
port 494 nsew default input
rlabel metal2 s 150410 -960 150522 480 8 la_oen[6]
port 495 nsew default input
rlabel metal2 s 378754 -960 378866 480 8 la_oen[70]
port 496 nsew default input
rlabel metal2 s 382342 -960 382454 480 8 la_oen[71]
port 497 nsew default input
rlabel metal2 s 385838 -960 385950 480 8 la_oen[72]
port 498 nsew default input
rlabel metal2 s 389426 -960 389538 480 8 la_oen[73]
port 499 nsew default input
rlabel metal2 s 393014 -960 393126 480 8 la_oen[74]
port 500 nsew default input
rlabel metal2 s 396602 -960 396714 480 8 la_oen[75]
port 501 nsew default input
rlabel metal2 s 400190 -960 400302 480 8 la_oen[76]
port 502 nsew default input
rlabel metal2 s 403686 -960 403798 480 8 la_oen[77]
port 503 nsew default input
rlabel metal2 s 407274 -960 407386 480 8 la_oen[78]
port 504 nsew default input
rlabel metal2 s 410862 -960 410974 480 8 la_oen[79]
port 505 nsew default input
rlabel metal2 s 153906 -960 154018 480 8 la_oen[7]
port 506 nsew default input
rlabel metal2 s 414450 -960 414562 480 8 la_oen[80]
port 507 nsew default input
rlabel metal2 s 417946 -960 418058 480 8 la_oen[81]
port 508 nsew default input
rlabel metal2 s 421534 -960 421646 480 8 la_oen[82]
port 509 nsew default input
rlabel metal2 s 425122 -960 425234 480 8 la_oen[83]
port 510 nsew default input
rlabel metal2 s 428710 -960 428822 480 8 la_oen[84]
port 511 nsew default input
rlabel metal2 s 432298 -960 432410 480 8 la_oen[85]
port 512 nsew default input
rlabel metal2 s 435794 -960 435906 480 8 la_oen[86]
port 513 nsew default input
rlabel metal2 s 439382 -960 439494 480 8 la_oen[87]
port 514 nsew default input
rlabel metal2 s 442970 -960 443082 480 8 la_oen[88]
port 515 nsew default input
rlabel metal2 s 446558 -960 446670 480 8 la_oen[89]
port 516 nsew default input
rlabel metal2 s 157494 -960 157606 480 8 la_oen[8]
port 517 nsew default input
rlabel metal2 s 450146 -960 450258 480 8 la_oen[90]
port 518 nsew default input
rlabel metal2 s 453642 -960 453754 480 8 la_oen[91]
port 519 nsew default input
rlabel metal2 s 457230 -960 457342 480 8 la_oen[92]
port 520 nsew default input
rlabel metal2 s 460818 -960 460930 480 8 la_oen[93]
port 521 nsew default input
rlabel metal2 s 464406 -960 464518 480 8 la_oen[94]
port 522 nsew default input
rlabel metal2 s 467902 -960 468014 480 8 la_oen[95]
port 523 nsew default input
rlabel metal2 s 471490 -960 471602 480 8 la_oen[96]
port 524 nsew default input
rlabel metal2 s 475078 -960 475190 480 8 la_oen[97]
port 525 nsew default input
rlabel metal2 s 478666 -960 478778 480 8 la_oen[98]
port 526 nsew default input
rlabel metal2 s 482254 -960 482366 480 8 la_oen[99]
port 527 nsew default input
rlabel metal2 s 161082 -960 161194 480 8 la_oen[9]
port 528 nsew default input
rlabel metal2 s 583362 -960 583474 480 8 user_clock2
port 529 nsew default input
rlabel metal2 s 542 -960 654 480 8 wb_clk_i
port 530 nsew default input
rlabel metal2 s 1646 -960 1758 480 8 wb_rst_i
port 531 nsew default input
rlabel metal2 s 2842 -960 2954 480 8 wbs_ack_o
port 532 nsew default tristate
rlabel metal2 s 7626 -960 7738 480 8 wbs_adr_i[0]
port 533 nsew default input
rlabel metal2 s 48106 -960 48218 480 8 wbs_adr_i[10]
port 534 nsew default input
rlabel metal2 s 51602 -960 51714 480 8 wbs_adr_i[11]
port 535 nsew default input
rlabel metal2 s 55190 -960 55302 480 8 wbs_adr_i[12]
port 536 nsew default input
rlabel metal2 s 58778 -960 58890 480 8 wbs_adr_i[13]
port 537 nsew default input
rlabel metal2 s 62366 -960 62478 480 8 wbs_adr_i[14]
port 538 nsew default input
rlabel metal2 s 65954 -960 66066 480 8 wbs_adr_i[15]
port 539 nsew default input
rlabel metal2 s 69450 -960 69562 480 8 wbs_adr_i[16]
port 540 nsew default input
rlabel metal2 s 73038 -960 73150 480 8 wbs_adr_i[17]
port 541 nsew default input
rlabel metal2 s 76626 -960 76738 480 8 wbs_adr_i[18]
port 542 nsew default input
rlabel metal2 s 80214 -960 80326 480 8 wbs_adr_i[19]
port 543 nsew default input
rlabel metal2 s 12410 -960 12522 480 8 wbs_adr_i[1]
port 544 nsew default input
rlabel metal2 s 83802 -960 83914 480 8 wbs_adr_i[20]
port 545 nsew default input
rlabel metal2 s 87298 -960 87410 480 8 wbs_adr_i[21]
port 546 nsew default input
rlabel metal2 s 90886 -960 90998 480 8 wbs_adr_i[22]
port 547 nsew default input
rlabel metal2 s 94474 -960 94586 480 8 wbs_adr_i[23]
port 548 nsew default input
rlabel metal2 s 98062 -960 98174 480 8 wbs_adr_i[24]
port 549 nsew default input
rlabel metal2 s 101558 -960 101670 480 8 wbs_adr_i[25]
port 550 nsew default input
rlabel metal2 s 105146 -960 105258 480 8 wbs_adr_i[26]
port 551 nsew default input
rlabel metal2 s 108734 -960 108846 480 8 wbs_adr_i[27]
port 552 nsew default input
rlabel metal2 s 112322 -960 112434 480 8 wbs_adr_i[28]
port 553 nsew default input
rlabel metal2 s 115910 -960 116022 480 8 wbs_adr_i[29]
port 554 nsew default input
rlabel metal2 s 17194 -960 17306 480 8 wbs_adr_i[2]
port 555 nsew default input
rlabel metal2 s 119406 -960 119518 480 8 wbs_adr_i[30]
port 556 nsew default input
rlabel metal2 s 122994 -960 123106 480 8 wbs_adr_i[31]
port 557 nsew default input
rlabel metal2 s 21886 -960 21998 480 8 wbs_adr_i[3]
port 558 nsew default input
rlabel metal2 s 26670 -960 26782 480 8 wbs_adr_i[4]
port 559 nsew default input
rlabel metal2 s 30258 -960 30370 480 8 wbs_adr_i[5]
port 560 nsew default input
rlabel metal2 s 33846 -960 33958 480 8 wbs_adr_i[6]
port 561 nsew default input
rlabel metal2 s 37342 -960 37454 480 8 wbs_adr_i[7]
port 562 nsew default input
rlabel metal2 s 40930 -960 41042 480 8 wbs_adr_i[8]
port 563 nsew default input
rlabel metal2 s 44518 -960 44630 480 8 wbs_adr_i[9]
port 564 nsew default input
rlabel metal2 s 4038 -960 4150 480 8 wbs_cyc_i
port 565 nsew default input
rlabel metal2 s 8822 -960 8934 480 8 wbs_dat_i[0]
port 566 nsew default input
rlabel metal2 s 49302 -960 49414 480 8 wbs_dat_i[10]
port 567 nsew default input
rlabel metal2 s 52798 -960 52910 480 8 wbs_dat_i[11]
port 568 nsew default input
rlabel metal2 s 56386 -960 56498 480 8 wbs_dat_i[12]
port 569 nsew default input
rlabel metal2 s 59974 -960 60086 480 8 wbs_dat_i[13]
port 570 nsew default input
rlabel metal2 s 63562 -960 63674 480 8 wbs_dat_i[14]
port 571 nsew default input
rlabel metal2 s 67150 -960 67262 480 8 wbs_dat_i[15]
port 572 nsew default input
rlabel metal2 s 70646 -960 70758 480 8 wbs_dat_i[16]
port 573 nsew default input
rlabel metal2 s 74234 -960 74346 480 8 wbs_dat_i[17]
port 574 nsew default input
rlabel metal2 s 77822 -960 77934 480 8 wbs_dat_i[18]
port 575 nsew default input
rlabel metal2 s 81410 -960 81522 480 8 wbs_dat_i[19]
port 576 nsew default input
rlabel metal2 s 13606 -960 13718 480 8 wbs_dat_i[1]
port 577 nsew default input
rlabel metal2 s 84906 -960 85018 480 8 wbs_dat_i[20]
port 578 nsew default input
rlabel metal2 s 88494 -960 88606 480 8 wbs_dat_i[21]
port 579 nsew default input
rlabel metal2 s 92082 -960 92194 480 8 wbs_dat_i[22]
port 580 nsew default input
rlabel metal2 s 95670 -960 95782 480 8 wbs_dat_i[23]
port 581 nsew default input
rlabel metal2 s 99258 -960 99370 480 8 wbs_dat_i[24]
port 582 nsew default input
rlabel metal2 s 102754 -960 102866 480 8 wbs_dat_i[25]
port 583 nsew default input
rlabel metal2 s 106342 -960 106454 480 8 wbs_dat_i[26]
port 584 nsew default input
rlabel metal2 s 109930 -960 110042 480 8 wbs_dat_i[27]
port 585 nsew default input
rlabel metal2 s 113518 -960 113630 480 8 wbs_dat_i[28]
port 586 nsew default input
rlabel metal2 s 117106 -960 117218 480 8 wbs_dat_i[29]
port 587 nsew default input
rlabel metal2 s 18298 -960 18410 480 8 wbs_dat_i[2]
port 588 nsew default input
rlabel metal2 s 120602 -960 120714 480 8 wbs_dat_i[30]
port 589 nsew default input
rlabel metal2 s 124190 -960 124302 480 8 wbs_dat_i[31]
port 590 nsew default input
rlabel metal2 s 23082 -960 23194 480 8 wbs_dat_i[3]
port 591 nsew default input
rlabel metal2 s 27866 -960 27978 480 8 wbs_dat_i[4]
port 592 nsew default input
rlabel metal2 s 31454 -960 31566 480 8 wbs_dat_i[5]
port 593 nsew default input
rlabel metal2 s 34950 -960 35062 480 8 wbs_dat_i[6]
port 594 nsew default input
rlabel metal2 s 38538 -960 38650 480 8 wbs_dat_i[7]
port 595 nsew default input
rlabel metal2 s 42126 -960 42238 480 8 wbs_dat_i[8]
port 596 nsew default input
rlabel metal2 s 45714 -960 45826 480 8 wbs_dat_i[9]
port 597 nsew default input
rlabel metal2 s 10018 -960 10130 480 8 wbs_dat_o[0]
port 598 nsew default tristate
rlabel metal2 s 50498 -960 50610 480 8 wbs_dat_o[10]
port 599 nsew default tristate
rlabel metal2 s 53994 -960 54106 480 8 wbs_dat_o[11]
port 600 nsew default tristate
rlabel metal2 s 57582 -960 57694 480 8 wbs_dat_o[12]
port 601 nsew default tristate
rlabel metal2 s 61170 -960 61282 480 8 wbs_dat_o[13]
port 602 nsew default tristate
rlabel metal2 s 64758 -960 64870 480 8 wbs_dat_o[14]
port 603 nsew default tristate
rlabel metal2 s 68254 -960 68366 480 8 wbs_dat_o[15]
port 604 nsew default tristate
rlabel metal2 s 71842 -960 71954 480 8 wbs_dat_o[16]
port 605 nsew default tristate
rlabel metal2 s 75430 -960 75542 480 8 wbs_dat_o[17]
port 606 nsew default tristate
rlabel metal2 s 79018 -960 79130 480 8 wbs_dat_o[18]
port 607 nsew default tristate
rlabel metal2 s 82606 -960 82718 480 8 wbs_dat_o[19]
port 608 nsew default tristate
rlabel metal2 s 14802 -960 14914 480 8 wbs_dat_o[1]
port 609 nsew default tristate
rlabel metal2 s 86102 -960 86214 480 8 wbs_dat_o[20]
port 610 nsew default tristate
rlabel metal2 s 89690 -960 89802 480 8 wbs_dat_o[21]
port 611 nsew default tristate
rlabel metal2 s 93278 -960 93390 480 8 wbs_dat_o[22]
port 612 nsew default tristate
rlabel metal2 s 96866 -960 96978 480 8 wbs_dat_o[23]
port 613 nsew default tristate
rlabel metal2 s 100454 -960 100566 480 8 wbs_dat_o[24]
port 614 nsew default tristate
rlabel metal2 s 103950 -960 104062 480 8 wbs_dat_o[25]
port 615 nsew default tristate
rlabel metal2 s 107538 -960 107650 480 8 wbs_dat_o[26]
port 616 nsew default tristate
rlabel metal2 s 111126 -960 111238 480 8 wbs_dat_o[27]
port 617 nsew default tristate
rlabel metal2 s 114714 -960 114826 480 8 wbs_dat_o[28]
port 618 nsew default tristate
rlabel metal2 s 118210 -960 118322 480 8 wbs_dat_o[29]
port 619 nsew default tristate
rlabel metal2 s 19494 -960 19606 480 8 wbs_dat_o[2]
port 620 nsew default tristate
rlabel metal2 s 121798 -960 121910 480 8 wbs_dat_o[30]
port 621 nsew default tristate
rlabel metal2 s 125386 -960 125498 480 8 wbs_dat_o[31]
port 622 nsew default tristate
rlabel metal2 s 24278 -960 24390 480 8 wbs_dat_o[3]
port 623 nsew default tristate
rlabel metal2 s 29062 -960 29174 480 8 wbs_dat_o[4]
port 624 nsew default tristate
rlabel metal2 s 32650 -960 32762 480 8 wbs_dat_o[5]
port 625 nsew default tristate
rlabel metal2 s 36146 -960 36258 480 8 wbs_dat_o[6]
port 626 nsew default tristate
rlabel metal2 s 39734 -960 39846 480 8 wbs_dat_o[7]
port 627 nsew default tristate
rlabel metal2 s 43322 -960 43434 480 8 wbs_dat_o[8]
port 628 nsew default tristate
rlabel metal2 s 46910 -960 47022 480 8 wbs_dat_o[9]
port 629 nsew default tristate
rlabel metal2 s 11214 -960 11326 480 8 wbs_sel_i[0]
port 630 nsew default input
rlabel metal2 s 15998 -960 16110 480 8 wbs_sel_i[1]
port 631 nsew default input
rlabel metal2 s 20690 -960 20802 480 8 wbs_sel_i[2]
port 632 nsew default input
rlabel metal2 s 25474 -960 25586 480 8 wbs_sel_i[3]
port 633 nsew default input
rlabel metal2 s 5234 -960 5346 480 8 wbs_stb_i
port 634 nsew default input
rlabel metal2 s 6430 -960 6542 480 8 wbs_we_i
port 635 nsew default input
rlabel metal5 s -1996 -924 585920 -324 8 vccd1
port 636 nsew default input
rlabel metal5 s -2936 -1864 586860 -1264 8 vssd1
port 637 nsew default input
rlabel metal5 s -3876 -2804 587800 -2204 8 vccd2
port 638 nsew default input
rlabel metal5 s -4816 -3744 588740 -3144 8 vssd2
port 639 nsew default input
rlabel metal5 s -5756 -4684 589680 -4084 8 vdda1
port 640 nsew default input
rlabel metal5 s -6696 -5624 590620 -5024 8 vssa1
port 641 nsew default input
rlabel metal5 s -7636 -6564 591560 -5964 8 vdda2
port 642 nsew default input
rlabel metal5 s -8576 -7504 592500 -6904 8 vssa2
port 643 nsew default input
<< properties >>
string FIXED_BBOX 0 0 584000 704000
<< end >>
