VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO spinet5
  CLASS BLOCK ;
  FOREIGN spinet5 ;
  ORIGIN 0.000 0.000 ;
  SIZE 333.390 BY 344.110 ;
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 187.770 340.110 188.050 344.110 ;
    END
  END clk
  PIN io_in[0]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 315.650 340.110 315.930 344.110 ;
    END
  END io_in[0]
  PIN io_in[10]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 87.080 4.000 87.680 ;
    END
  END io_in[10]
  PIN io_in[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 340.110 45.450 344.110 ;
    END
  END io_in[11]
  PIN io_in[12]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 329.390 233.960 333.390 234.560 ;
    END
  END io_in[12]
  PIN io_in[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 130.730 0.000 131.010 4.000 ;
    END
  END io_in[13]
  PIN io_in[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 159.250 0.000 159.530 4.000 ;
    END
  END io_in[14]
  PIN io_in[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 329.390 276.120 333.390 276.720 ;
    END
  END io_in[15]
  PIN io_in[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 201.570 340.110 201.850 344.110 ;
    END
  END io_in[16]
  PIN io_in[17]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 44.920 4.000 45.520 ;
    END
  END io_in[17]
  PIN io_in[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END io_in[18]
  PIN io_in[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 273.330 340.110 273.610 344.110 ;
    END
  END io_in[19]
  PIN io_in[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 173.050 0.000 173.330 4.000 ;
    END
  END io_in[1]
  PIN io_in[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 116.930 340.110 117.210 344.110 ;
    END
  END io_in[20]
  PIN io_in[21]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 329.390 213.560 333.390 214.160 ;
    END
  END io_in[21]
  PIN io_in[22]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 30.450 0.000 30.730 4.000 ;
    END
  END io_in[22]
  PIN io_in[23]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 108.840 4.000 109.440 ;
    END
  END io_in[23]
  PIN io_in[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 216.290 340.110 216.570 344.110 ;
    END
  END io_in[24]
  PIN io_in[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 272.410 0.000 272.690 4.000 ;
    END
  END io_in[25]
  PIN io_in[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 329.390 44.920 333.390 45.520 ;
    END
  END io_in[26]
  PIN io_in[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.160 4.000 193.760 ;
    END
  END io_in[27]
  PIN io_in[28]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 329.450 340.110 329.730 344.110 ;
    END
  END io_in[28]
  PIN io_in[29]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 130.730 340.110 131.010 344.110 ;
    END
  END io_in[29]
  PIN io_in[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END io_in[2]
  PIN io_in[30]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END io_in[30]
  PIN io_in[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 73.690 0.000 73.970 4.000 ;
    END
  END io_in[31]
  PIN io_in[32]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 329.390 297.880 333.390 298.480 ;
    END
  END io_in[32]
  PIN io_in[33]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 16.650 340.110 16.930 344.110 ;
    END
  END io_in[33]
  PIN io_in[34]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 31.370 340.110 31.650 344.110 ;
    END
  END io_in[34]
  PIN io_in[35]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 258.610 340.110 258.890 344.110 ;
    END
  END io_in[35]
  PIN io_in[36]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 59.890 340.110 60.170 344.110 ;
    END
  END io_in[36]
  PIN io_in[37]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 329.450 0.000 329.730 4.000 ;
    END
  END io_in[37]
  PIN io_in[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.720 4.000 256.320 ;
    END
  END io_in[3]
  PIN io_in[4]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 329.390 66.680 333.390 67.280 ;
    END
  END io_in[4]
  PIN io_in[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 340.110 3.130 344.110 ;
    END
  END io_in[5]
  PIN io_in[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 58.970 0.000 59.250 4.000 ;
    END
  END io_in[6]
  PIN io_in[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END io_in[7]
  PIN io_in[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 187.770 0.000 188.050 4.000 ;
    END
  END io_in[8]
  PIN io_in[9]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 24.520 4.000 25.120 ;
    END
  END io_in[9]
  PIN io_out[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END io_out[0]
  PIN io_out[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END io_out[10]
  PIN io_out[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 230.090 340.110 230.370 344.110 ;
    END
  END io_out[11]
  PIN io_out[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 16.650 0.000 16.930 4.000 ;
    END
  END io_out[12]
  PIN io_out[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 329.390 191.800 333.390 192.400 ;
    END
  END io_out[13]
  PIN io_out[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 300.930 0.000 301.210 4.000 ;
    END
  END io_out[14]
  PIN io_out[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 173.050 340.110 173.330 344.110 ;
    END
  END io_out[15]
  PIN io_out[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 329.390 318.280 333.390 318.880 ;
    END
  END io_out[16]
  PIN io_out[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 329.390 171.400 333.390 172.000 ;
    END
  END io_out[17]
  PIN io_out[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 329.390 24.520 333.390 25.120 ;
    END
  END io_out[18]
  PIN io_out[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END io_out[19]
  PIN io_out[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 88.410 340.110 88.690 344.110 ;
    END
  END io_out[1]
  PIN io_out[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 329.390 149.640 333.390 150.240 ;
    END
  END io_out[20]
  PIN io_out[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 329.390 129.240 333.390 129.840 ;
    END
  END io_out[21]
  PIN io_out[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 159.250 340.110 159.530 344.110 ;
    END
  END io_out[22]
  PIN io_out[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 301.850 340.110 302.130 344.110 ;
    END
  END io_out[23]
  PIN io_out[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 213.560 4.000 214.160 ;
    END
  END io_out[24]
  PIN io_out[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END io_out[25]
  PIN io_out[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 276.120 4.000 276.720 ;
    END
  END io_out[26]
  PIN io_out[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.210 0.000 102.490 4.000 ;
    END
  END io_out[27]
  PIN io_out[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END io_out[28]
  PIN io_out[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 297.880 4.000 298.480 ;
    END
  END io_out[29]
  PIN io_out[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 201.570 0.000 201.850 4.000 ;
    END
  END io_out[2]
  PIN io_out[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 258.610 0.000 258.890 4.000 ;
    END
  END io_out[30]
  PIN io_out[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 244.810 340.110 245.090 344.110 ;
    END
  END io_out[31]
  PIN io_out[32]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 151.000 4.000 151.600 ;
    END
  END io_out[32]
  PIN io_out[33]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 329.390 87.080 333.390 87.680 ;
    END
  END io_out[33]
  PIN io_out[34]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 235.320 4.000 235.920 ;
    END
  END io_out[34]
  PIN io_out[35]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 144.530 340.110 144.810 344.110 ;
    END
  END io_out[35]
  PIN io_out[36]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 329.390 107.480 333.390 108.080 ;
    END
  END io_out[36]
  PIN io_out[37]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 171.400 4.000 172.000 ;
    END
  END io_out[37]
  PIN io_out[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 230.090 0.000 230.370 4.000 ;
    END
  END io_out[3]
  PIN io_out[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 102.210 340.110 102.490 344.110 ;
    END
  END io_out[4]
  PIN io_out[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 287.130 0.000 287.410 4.000 ;
    END
  END io_out[5]
  PIN io_out[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 243.890 0.000 244.170 4.000 ;
    END
  END io_out[6]
  PIN io_out[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 287.130 340.110 287.410 344.110 ;
    END
  END io_out[7]
  PIN io_out[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 329.390 255.720 333.390 256.320 ;
    END
  END io_out[8]
  PIN io_out[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 73.690 340.110 73.970 344.110 ;
    END
  END io_out[9]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 144.530 0.000 144.810 4.000 ;
    END
  END rst
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 332.080 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 332.080 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 327.520 331.925 ;
      LAYER met1 ;
        RECT 2.830 10.640 329.750 332.080 ;
      LAYER met2 ;
        RECT 3.410 339.830 16.370 340.110 ;
        RECT 17.210 339.830 31.090 340.110 ;
        RECT 31.930 339.830 44.890 340.110 ;
        RECT 45.730 339.830 59.610 340.110 ;
        RECT 60.450 339.830 73.410 340.110 ;
        RECT 74.250 339.830 88.130 340.110 ;
        RECT 88.970 339.830 101.930 340.110 ;
        RECT 102.770 339.830 116.650 340.110 ;
        RECT 117.490 339.830 130.450 340.110 ;
        RECT 131.290 339.830 144.250 340.110 ;
        RECT 145.090 339.830 158.970 340.110 ;
        RECT 159.810 339.830 172.770 340.110 ;
        RECT 173.610 339.830 187.490 340.110 ;
        RECT 188.330 339.830 201.290 340.110 ;
        RECT 202.130 339.830 216.010 340.110 ;
        RECT 216.850 339.830 229.810 340.110 ;
        RECT 230.650 339.830 244.530 340.110 ;
        RECT 245.370 339.830 258.330 340.110 ;
        RECT 259.170 339.830 273.050 340.110 ;
        RECT 273.890 339.830 286.850 340.110 ;
        RECT 287.690 339.830 301.570 340.110 ;
        RECT 302.410 339.830 315.370 340.110 ;
        RECT 316.210 339.830 329.170 340.110 ;
        RECT 2.860 4.280 329.720 339.830 ;
        RECT 3.410 4.000 16.370 4.280 ;
        RECT 17.210 4.000 30.170 4.280 ;
        RECT 31.010 4.000 44.890 4.280 ;
        RECT 45.730 4.000 58.690 4.280 ;
        RECT 59.530 4.000 73.410 4.280 ;
        RECT 74.250 4.000 87.210 4.280 ;
        RECT 88.050 4.000 101.930 4.280 ;
        RECT 102.770 4.000 115.730 4.280 ;
        RECT 116.570 4.000 130.450 4.280 ;
        RECT 131.290 4.000 144.250 4.280 ;
        RECT 145.090 4.000 158.970 4.280 ;
        RECT 159.810 4.000 172.770 4.280 ;
        RECT 173.610 4.000 187.490 4.280 ;
        RECT 188.330 4.000 201.290 4.280 ;
        RECT 202.130 4.000 215.090 4.280 ;
        RECT 215.930 4.000 229.810 4.280 ;
        RECT 230.650 4.000 243.610 4.280 ;
        RECT 244.450 4.000 258.330 4.280 ;
        RECT 259.170 4.000 272.130 4.280 ;
        RECT 272.970 4.000 286.850 4.280 ;
        RECT 287.690 4.000 300.650 4.280 ;
        RECT 301.490 4.000 315.370 4.280 ;
        RECT 316.210 4.000 329.170 4.280 ;
      LAYER met3 ;
        RECT 4.000 319.280 329.390 332.005 ;
        RECT 4.400 317.880 328.990 319.280 ;
        RECT 4.000 298.880 329.390 317.880 ;
        RECT 4.400 297.480 328.990 298.880 ;
        RECT 4.000 277.120 329.390 297.480 ;
        RECT 4.400 275.720 328.990 277.120 ;
        RECT 4.000 256.720 329.390 275.720 ;
        RECT 4.400 255.320 328.990 256.720 ;
        RECT 4.000 236.320 329.390 255.320 ;
        RECT 4.400 234.960 329.390 236.320 ;
        RECT 4.400 234.920 328.990 234.960 ;
        RECT 4.000 233.560 328.990 234.920 ;
        RECT 4.000 214.560 329.390 233.560 ;
        RECT 4.400 213.160 328.990 214.560 ;
        RECT 4.000 194.160 329.390 213.160 ;
        RECT 4.400 192.800 329.390 194.160 ;
        RECT 4.400 192.760 328.990 192.800 ;
        RECT 4.000 191.400 328.990 192.760 ;
        RECT 4.000 172.400 329.390 191.400 ;
        RECT 4.400 171.000 328.990 172.400 ;
        RECT 4.000 152.000 329.390 171.000 ;
        RECT 4.400 150.640 329.390 152.000 ;
        RECT 4.400 150.600 328.990 150.640 ;
        RECT 4.000 149.240 328.990 150.600 ;
        RECT 4.000 130.240 329.390 149.240 ;
        RECT 4.400 128.840 328.990 130.240 ;
        RECT 4.000 109.840 329.390 128.840 ;
        RECT 4.400 108.480 329.390 109.840 ;
        RECT 4.400 108.440 328.990 108.480 ;
        RECT 4.000 107.080 328.990 108.440 ;
        RECT 4.000 88.080 329.390 107.080 ;
        RECT 4.400 86.680 328.990 88.080 ;
        RECT 4.000 67.680 329.390 86.680 ;
        RECT 4.400 66.280 328.990 67.680 ;
        RECT 4.000 45.920 329.390 66.280 ;
        RECT 4.400 44.520 328.990 45.920 ;
        RECT 4.000 25.520 329.390 44.520 ;
        RECT 4.400 24.120 328.990 25.520 ;
        RECT 4.000 10.715 329.390 24.120 ;
      LAYER met4 ;
        RECT 174.640 10.640 253.040 332.080 ;
  END
END spinet5
END LIBRARY

