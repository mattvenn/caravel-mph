VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO asic_freq
  CLASS BLOCK ;
  FOREIGN asic_freq ;
  ORIGIN 0.000 0.000 ;
  SIZE 389.335 BY 400.055 ;
  PIN addr[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 385.335 206.760 389.335 207.360 ;
    END
  END addr[0]
  PIN addr[1]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 318.280 4.000 318.880 ;
    END
  END addr[1]
  PIN addr[2]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 247.570 396.055 247.850 400.055 ;
    END
  END addr[2]
  PIN addr[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 385.335 363.160 389.335 363.760 ;
    END
  END addr[3]
  PIN clk
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 35.050 396.055 35.330 400.055 ;
    END
  END clk
  PIN col_drvs[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 191.800 4.000 192.400 ;
    END
  END col_drvs[0]
  PIN col_drvs[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 119.690 0.000 119.970 4.000 ;
    END
  END col_drvs[1]
  PIN col_drvs[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 385.570 0.000 385.850 4.000 ;
    END
  END col_drvs[2]
  PIN col_drvs[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 385.335 190.440 389.335 191.040 ;
    END
  END col_drvs[3]
  PIN col_drvs[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 50.360 4.000 50.960 ;
    END
  END col_drvs[4]
  PIN col_drvs[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END col_drvs[5]
  PIN col_drvs[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 385.335 111.560 389.335 112.160 ;
    END
  END col_drvs[6]
  PIN col_drvs[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 129.810 0.000 130.090 4.000 ;
    END
  END col_drvs[7]
  PIN col_drvs[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 385.335 285.640 389.335 286.240 ;
    END
  END col_drvs[8]
  PIN o[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 353.370 0.000 353.650 4.000 ;
    END
  END o[0]
  PIN o[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 141.770 396.055 142.050 400.055 ;
    END
  END o[10]
  PIN o[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 258.610 396.055 258.890 400.055 ;
    END
  END o[11]
  PIN o[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 385.335 175.480 389.335 176.080 ;
    END
  END o[12]
  PIN o[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 204.330 0.000 204.610 4.000 ;
    END
  END o[13]
  PIN o[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 267.810 0.000 268.090 4.000 ;
    END
  END o[14]
  PIN o[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 300.930 396.055 301.210 400.055 ;
    END
  END o[15]
  PIN o[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 385.335 49.000 389.335 49.600 ;
    END
  END o[16]
  PIN o[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 385.335 269.320 389.335 269.920 ;
    END
  END o[17]
  PIN o[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 162.010 0.000 162.290 4.000 ;
    END
  END o[18]
  PIN o[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 270.680 4.000 271.280 ;
    END
  END o[19]
  PIN o[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 55.290 0.000 55.570 4.000 ;
    END
  END o[1]
  PIN o[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 385.335 17.720 389.335 18.320 ;
    END
  END o[20]
  PIN o[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 385.570 396.055 385.850 400.055 ;
    END
  END o[21]
  PIN o[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 162.930 396.055 163.210 400.055 ;
    END
  END o[22]
  PIN o[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 205.250 396.055 205.530 400.055 ;
    END
  END o[23]
  PIN o[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 385.335 348.200 389.335 348.800 ;
    END
  END o[24]
  PIN o[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 246.650 0.000 246.930 4.000 ;
    END
  END o[25]
  PIN o[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 333.130 396.055 333.410 400.055 ;
    END
  END o[26]
  PIN o[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 278.850 0.000 279.130 4.000 ;
    END
  END o[27]
  PIN o[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 375.450 396.055 375.730 400.055 ;
    END
  END o[28]
  PIN o[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END o[29]
  PIN o[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 34.130 0.000 34.410 4.000 ;
    END
  END o[2]
  PIN o[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 140.850 0.000 141.130 4.000 ;
    END
  END o[30]
  PIN o[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 301.960 4.000 302.560 ;
    END
  END o[31]
  PIN o[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 87.490 0.000 87.770 4.000 ;
    END
  END o[3]
  PIN o[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 97.960 4.000 98.560 ;
    END
  END o[4]
  PIN o[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 385.335 159.160 389.335 159.760 ;
    END
  END o[5]
  PIN o[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END o[6]
  PIN o[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 342.330 0.000 342.610 4.000 ;
    END
  END o[7]
  PIN o[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END o[8]
  PIN o[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 385.335 221.720 389.335 222.320 ;
    END
  END o[9]
  PIN oc[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 287.000 4.000 287.600 ;
    END
  END oc[0]
  PIN oc[10]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 332.210 0.000 332.490 4.000 ;
    END
  END oc[10]
  PIN oc[11]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END oc[11]
  PIN oc[12]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 194.210 396.055 194.490 400.055 ;
    END
  END oc[12]
  PIN oc[13]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 385.335 316.920 389.335 317.520 ;
    END
  END oc[13]
  PIN oc[14]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 160.520 4.000 161.120 ;
    END
  END oc[14]
  PIN oc[15]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 311.050 0.000 311.330 4.000 ;
    END
  END oc[15]
  PIN oc[16]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 385.335 238.040 389.335 238.640 ;
    END
  END oc[16]
  PIN oc[17]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 385.335 80.280 389.335 80.880 ;
    END
  END oc[17]
  PIN oc[18]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END oc[18]
  PIN oc[19]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 239.400 4.000 240.000 ;
    END
  END oc[19]
  PIN oc[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 343.250 396.055 343.530 400.055 ;
    END
  END oc[1]
  PIN oc[20]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 76.450 0.000 76.730 4.000 ;
    END
  END oc[20]
  PIN oc[21]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 364.410 396.055 364.690 400.055 ;
    END
  END oc[21]
  PIN oc[22]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 354.290 396.055 354.570 400.055 ;
    END
  END oc[22]
  PIN oc[23]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 254.360 4.000 254.960 ;
    END
  END oc[23]
  PIN oc[24]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 2.850 396.055 3.130 400.055 ;
    END
  END oc[24]
  PIN oc[25]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END oc[25]
  PIN oc[26]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 279.770 396.055 280.050 400.055 ;
    END
  END oc[26]
  PIN oc[27]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 289.890 0.000 290.170 4.000 ;
    END
  END oc[27]
  PIN oc[28]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.930 396.055 25.210 400.055 ;
    END
  END oc[28]
  PIN oc[29]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 385.335 253.000 389.335 253.600 ;
    END
  END oc[29]
  PIN oc[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 98.530 396.055 98.810 400.055 ;
    END
  END oc[2]
  PIN oc[30]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 289.890 396.055 290.170 400.055 ;
    END
  END oc[30]
  PIN oc[31]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 19.080 4.000 19.680 ;
    END
  END oc[31]
  PIN oc[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 385.335 300.600 389.335 301.200 ;
    END
  END oc[3]
  PIN oc[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.920 4.000 113.520 ;
    END
  END oc[4]
  PIN oc[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 130.730 396.055 131.010 400.055 ;
    END
  END oc[5]
  PIN oc[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 67.250 396.055 67.530 400.055 ;
    END
  END oc[6]
  PIN oc[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 374.530 0.000 374.810 4.000 ;
    END
  END oc[7]
  PIN oc[8]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 385.335 331.880 389.335 332.480 ;
    END
  END oc[8]
  PIN oc[9]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 108.650 0.000 108.930 4.000 ;
    END
  END oc[9]
  PIN rst
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 385.335 127.880 389.335 128.480 ;
    END
  END rst
  PIN samplee
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 268.730 396.055 269.010 400.055 ;
    END
  END samplee
  PIN seg_drvs[0]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 46.090 396.055 46.370 400.055 ;
    END
  END seg_drvs[0]
  PIN seg_drvs[1]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 66.680 4.000 67.280 ;
    END
  END seg_drvs[1]
  PIN seg_drvs[2]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 0.000 223.080 4.000 223.680 ;
    END
  END seg_drvs[2]
  PIN seg_drvs[3]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 109.570 396.055 109.850 400.055 ;
    END
  END seg_drvs[3]
  PIN seg_drvs[4]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 24.010 0.000 24.290 4.000 ;
    END
  END seg_drvs[4]
  PIN seg_drvs[5]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 183.170 0.000 183.450 4.000 ;
    END
  END seg_drvs[5]
  PIN seg_drvs[6]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 311.970 396.055 312.250 400.055 ;
    END
  END seg_drvs[6]
  PIN seg_drvs[7]
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met3 ;
        RECT 385.335 65.320 389.335 65.920 ;
    END
  END seg_drvs[7]
  PIN strobe
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 349.560 4.000 350.160 ;
    END
  END strobe
  PIN tx
    DIRECTION OUTPUT TRISTATE ;
    PORT
      LAYER met2 ;
        RECT 215.370 0.000 215.650 4.000 ;
    END
  END tx
  PIN value[0]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 385.335 96.600 389.335 97.200 ;
    END
  END value[0]
  PIN value[10]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 56.210 396.055 56.490 400.055 ;
    END
  END value[10]
  PIN value[11]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 77.370 396.055 77.650 400.055 ;
    END
  END value[11]
  PIN value[12]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 236.530 0.000 236.810 4.000 ;
    END
  END value[12]
  PIN value[13]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 363.490 0.000 363.770 4.000 ;
    END
  END value[13]
  PIN value[14]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 322.090 396.055 322.370 400.055 ;
    END
  END value[14]
  PIN value[15]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 385.335 34.040 389.335 34.640 ;
    END
  END value[15]
  PIN value[16]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 194.210 0.000 194.490 4.000 ;
    END
  END value[16]
  PIN value[17]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 88.410 396.055 88.690 400.055 ;
    END
  END value[17]
  PIN value[18]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 321.170 0.000 321.450 4.000 ;
    END
  END value[18]
  PIN value[19]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 300.010 0.000 300.290 4.000 ;
    END
  END value[19]
  PIN value[1]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 184.090 396.055 184.370 400.055 ;
    END
  END value[1]
  PIN value[20]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 151.890 396.055 152.170 400.055 ;
    END
  END value[20]
  PIN value[21]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 173.050 396.055 173.330 400.055 ;
    END
  END value[21]
  PIN value[22]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 145.560 4.000 146.160 ;
    END
  END value[22]
  PIN value[23]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 237.450 396.055 237.730 400.055 ;
    END
  END value[23]
  PIN value[24]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 150.970 0.000 151.250 4.000 ;
    END
  END value[24]
  PIN value[25]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 2.850 0.000 3.130 4.000 ;
    END
  END value[25]
  PIN value[26]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 385.335 379.480 389.335 380.080 ;
    END
  END value[26]
  PIN value[27]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 208.120 4.000 208.720 ;
    END
  END value[27]
  PIN value[28]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 35.400 4.000 36.000 ;
    END
  END value[28]
  PIN value[29]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 385.335 144.200 389.335 144.800 ;
    END
  END value[29]
  PIN value[2]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 364.520 4.000 365.120 ;
    END
  END value[2]
  PIN value[30]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 13.890 396.055 14.170 400.055 ;
    END
  END value[30]
  PIN value[31]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 120.610 396.055 120.890 400.055 ;
    END
  END value[31]
  PIN value[3]
    DIRECTION INPUT ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END value[3]
  PIN value[4]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 66.330 0.000 66.610 4.000 ;
    END
  END value[4]
  PIN value[5]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 12.970 0.000 13.250 4.000 ;
    END
  END value[5]
  PIN value[6]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 216.290 396.055 216.570 400.055 ;
    END
  END value[6]
  PIN value[7]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 226.410 396.055 226.690 400.055 ;
    END
  END value[7]
  PIN value[8]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 98.530 0.000 98.810 4.000 ;
    END
  END value[8]
  PIN value[9]
    DIRECTION INPUT ;
    PORT
      LAYER met2 ;
        RECT 172.130 0.000 172.410 4.000 ;
    END
  END value[9]
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 389.200 ;
    END
  END VPWR
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 389.200 ;
    END
  END VGND
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 384.415 389.045 ;
      LAYER met1 ;
        RECT 2.830 4.460 385.870 389.200 ;
      LAYER met2 ;
        RECT 3.410 395.775 13.610 396.055 ;
        RECT 14.450 395.775 24.650 396.055 ;
        RECT 25.490 395.775 34.770 396.055 ;
        RECT 35.610 395.775 45.810 396.055 ;
        RECT 46.650 395.775 55.930 396.055 ;
        RECT 56.770 395.775 66.970 396.055 ;
        RECT 67.810 395.775 77.090 396.055 ;
        RECT 77.930 395.775 88.130 396.055 ;
        RECT 88.970 395.775 98.250 396.055 ;
        RECT 99.090 395.775 109.290 396.055 ;
        RECT 110.130 395.775 120.330 396.055 ;
        RECT 121.170 395.775 130.450 396.055 ;
        RECT 131.290 395.775 141.490 396.055 ;
        RECT 142.330 395.775 151.610 396.055 ;
        RECT 152.450 395.775 162.650 396.055 ;
        RECT 163.490 395.775 172.770 396.055 ;
        RECT 173.610 395.775 183.810 396.055 ;
        RECT 184.650 395.775 193.930 396.055 ;
        RECT 194.770 395.775 204.970 396.055 ;
        RECT 205.810 395.775 216.010 396.055 ;
        RECT 216.850 395.775 226.130 396.055 ;
        RECT 226.970 395.775 237.170 396.055 ;
        RECT 238.010 395.775 247.290 396.055 ;
        RECT 248.130 395.775 258.330 396.055 ;
        RECT 259.170 395.775 268.450 396.055 ;
        RECT 269.290 395.775 279.490 396.055 ;
        RECT 280.330 395.775 289.610 396.055 ;
        RECT 290.450 395.775 300.650 396.055 ;
        RECT 301.490 395.775 311.690 396.055 ;
        RECT 312.530 395.775 321.810 396.055 ;
        RECT 322.650 395.775 332.850 396.055 ;
        RECT 333.690 395.775 342.970 396.055 ;
        RECT 343.810 395.775 354.010 396.055 ;
        RECT 354.850 395.775 364.130 396.055 ;
        RECT 364.970 395.775 375.170 396.055 ;
        RECT 376.010 395.775 385.290 396.055 ;
        RECT 2.860 4.280 385.840 395.775 ;
        RECT 3.410 4.000 12.690 4.280 ;
        RECT 13.530 4.000 23.730 4.280 ;
        RECT 24.570 4.000 33.850 4.280 ;
        RECT 34.690 4.000 44.890 4.280 ;
        RECT 45.730 4.000 55.010 4.280 ;
        RECT 55.850 4.000 66.050 4.280 ;
        RECT 66.890 4.000 76.170 4.280 ;
        RECT 77.010 4.000 87.210 4.280 ;
        RECT 88.050 4.000 98.250 4.280 ;
        RECT 99.090 4.000 108.370 4.280 ;
        RECT 109.210 4.000 119.410 4.280 ;
        RECT 120.250 4.000 129.530 4.280 ;
        RECT 130.370 4.000 140.570 4.280 ;
        RECT 141.410 4.000 150.690 4.280 ;
        RECT 151.530 4.000 161.730 4.280 ;
        RECT 162.570 4.000 171.850 4.280 ;
        RECT 172.690 4.000 182.890 4.280 ;
        RECT 183.730 4.000 193.930 4.280 ;
        RECT 194.770 4.000 204.050 4.280 ;
        RECT 204.890 4.000 215.090 4.280 ;
        RECT 215.930 4.000 225.210 4.280 ;
        RECT 226.050 4.000 236.250 4.280 ;
        RECT 237.090 4.000 246.370 4.280 ;
        RECT 247.210 4.000 257.410 4.280 ;
        RECT 258.250 4.000 267.530 4.280 ;
        RECT 268.370 4.000 278.570 4.280 ;
        RECT 279.410 4.000 289.610 4.280 ;
        RECT 290.450 4.000 299.730 4.280 ;
        RECT 300.570 4.000 310.770 4.280 ;
        RECT 311.610 4.000 320.890 4.280 ;
        RECT 321.730 4.000 331.930 4.280 ;
        RECT 332.770 4.000 342.050 4.280 ;
        RECT 342.890 4.000 353.090 4.280 ;
        RECT 353.930 4.000 363.210 4.280 ;
        RECT 364.050 4.000 374.250 4.280 ;
        RECT 375.090 4.000 385.290 4.280 ;
      LAYER met3 ;
        RECT 4.000 381.840 385.335 389.125 ;
        RECT 4.400 380.480 385.335 381.840 ;
        RECT 4.400 380.440 384.935 380.480 ;
        RECT 4.000 379.080 384.935 380.440 ;
        RECT 4.000 365.520 385.335 379.080 ;
        RECT 4.400 364.160 385.335 365.520 ;
        RECT 4.400 364.120 384.935 364.160 ;
        RECT 4.000 362.760 384.935 364.120 ;
        RECT 4.000 350.560 385.335 362.760 ;
        RECT 4.400 349.200 385.335 350.560 ;
        RECT 4.400 349.160 384.935 349.200 ;
        RECT 4.000 347.800 384.935 349.160 ;
        RECT 4.000 334.240 385.335 347.800 ;
        RECT 4.400 332.880 385.335 334.240 ;
        RECT 4.400 332.840 384.935 332.880 ;
        RECT 4.000 331.480 384.935 332.840 ;
        RECT 4.000 319.280 385.335 331.480 ;
        RECT 4.400 317.920 385.335 319.280 ;
        RECT 4.400 317.880 384.935 317.920 ;
        RECT 4.000 316.520 384.935 317.880 ;
        RECT 4.000 302.960 385.335 316.520 ;
        RECT 4.400 301.600 385.335 302.960 ;
        RECT 4.400 301.560 384.935 301.600 ;
        RECT 4.000 300.200 384.935 301.560 ;
        RECT 4.000 288.000 385.335 300.200 ;
        RECT 4.400 286.640 385.335 288.000 ;
        RECT 4.400 286.600 384.935 286.640 ;
        RECT 4.000 285.240 384.935 286.600 ;
        RECT 4.000 271.680 385.335 285.240 ;
        RECT 4.400 270.320 385.335 271.680 ;
        RECT 4.400 270.280 384.935 270.320 ;
        RECT 4.000 268.920 384.935 270.280 ;
        RECT 4.000 255.360 385.335 268.920 ;
        RECT 4.400 254.000 385.335 255.360 ;
        RECT 4.400 253.960 384.935 254.000 ;
        RECT 4.000 252.600 384.935 253.960 ;
        RECT 4.000 240.400 385.335 252.600 ;
        RECT 4.400 239.040 385.335 240.400 ;
        RECT 4.400 239.000 384.935 239.040 ;
        RECT 4.000 237.640 384.935 239.000 ;
        RECT 4.000 224.080 385.335 237.640 ;
        RECT 4.400 222.720 385.335 224.080 ;
        RECT 4.400 222.680 384.935 222.720 ;
        RECT 4.000 221.320 384.935 222.680 ;
        RECT 4.000 209.120 385.335 221.320 ;
        RECT 4.400 207.760 385.335 209.120 ;
        RECT 4.400 207.720 384.935 207.760 ;
        RECT 4.000 206.360 384.935 207.720 ;
        RECT 4.000 192.800 385.335 206.360 ;
        RECT 4.400 191.440 385.335 192.800 ;
        RECT 4.400 191.400 384.935 191.440 ;
        RECT 4.000 190.040 384.935 191.400 ;
        RECT 4.000 177.840 385.335 190.040 ;
        RECT 4.400 176.480 385.335 177.840 ;
        RECT 4.400 176.440 384.935 176.480 ;
        RECT 4.000 175.080 384.935 176.440 ;
        RECT 4.000 161.520 385.335 175.080 ;
        RECT 4.400 160.160 385.335 161.520 ;
        RECT 4.400 160.120 384.935 160.160 ;
        RECT 4.000 158.760 384.935 160.120 ;
        RECT 4.000 146.560 385.335 158.760 ;
        RECT 4.400 145.200 385.335 146.560 ;
        RECT 4.400 145.160 384.935 145.200 ;
        RECT 4.000 143.800 384.935 145.160 ;
        RECT 4.000 130.240 385.335 143.800 ;
        RECT 4.400 128.880 385.335 130.240 ;
        RECT 4.400 128.840 384.935 128.880 ;
        RECT 4.000 127.480 384.935 128.840 ;
        RECT 4.000 113.920 385.335 127.480 ;
        RECT 4.400 112.560 385.335 113.920 ;
        RECT 4.400 112.520 384.935 112.560 ;
        RECT 4.000 111.160 384.935 112.520 ;
        RECT 4.000 98.960 385.335 111.160 ;
        RECT 4.400 97.600 385.335 98.960 ;
        RECT 4.400 97.560 384.935 97.600 ;
        RECT 4.000 96.200 384.935 97.560 ;
        RECT 4.000 82.640 385.335 96.200 ;
        RECT 4.400 81.280 385.335 82.640 ;
        RECT 4.400 81.240 384.935 81.280 ;
        RECT 4.000 79.880 384.935 81.240 ;
        RECT 4.000 67.680 385.335 79.880 ;
        RECT 4.400 66.320 385.335 67.680 ;
        RECT 4.400 66.280 384.935 66.320 ;
        RECT 4.000 64.920 384.935 66.280 ;
        RECT 4.000 51.360 385.335 64.920 ;
        RECT 4.400 50.000 385.335 51.360 ;
        RECT 4.400 49.960 384.935 50.000 ;
        RECT 4.000 48.600 384.935 49.960 ;
        RECT 4.000 36.400 385.335 48.600 ;
        RECT 4.400 35.040 385.335 36.400 ;
        RECT 4.400 35.000 384.935 35.040 ;
        RECT 4.000 33.640 384.935 35.000 ;
        RECT 4.000 20.080 385.335 33.640 ;
        RECT 4.400 18.720 385.335 20.080 ;
        RECT 4.400 18.680 384.935 18.720 ;
        RECT 4.000 17.320 384.935 18.680 ;
        RECT 4.000 10.715 385.335 17.320 ;
      LAYER met4 ;
        RECT 100.575 10.640 329.840 389.200 ;
  END
END asic_freq
END LIBRARY

